//685x685 
// Code your testbench here 
// or browse Examples 
// Verilog test bench for HHT with buffer 
`timescale 1ns/1ps 
module testbench; 
  parameter V_SIZE = 9; 
  parameter COL_SIZE = 1967 ; 
reg Clk,Rst,WR,mem_init; 
reg [31:0] dataIn1,dataIn2,csize; 
reg [31:0]v_values_base; 
wire [31:0]addr1,addr2; 
wire [4:0] regaddr1,regaddr2; 
reg[31:0] cpu_addr;
wire hht;
wire [31:0]val[0:8]; 
reg [31:0]wdata_col_base; 
wire [31:0] dataOut; 
reg fe_init; 
reg wn,rn,RD; 
wire [4:0]adata; 
wire [31:0] rdata; 
 // Instantiate memory module 
//  memmodel m1 (addr,dataIn,dataOut,WR,Clk,Rst); 
//  mem_buffer m1 (dataOut, full, empty, Clk, Rst, wn, rn, dataIn); 
control t1 (Clk,wdata_col_base,v_values_base,addr1,addr2,dataIn1,dataIn2,Rst,RD,csize,cpu_addr,hht,regaddr1,regaddr2,rdata,adata); ;  
//frontend t1 (Clk,Rst,fe_init,wdata_col_base,data_req,dataIn,init, 
//{m_cols[0],m_cols[1],m_cols[2],m_cols[3],m_cols[4]}, 
//done,wn); 
initial begin 
Clk = 1'b0; 
  RD = 1'b1; 
 #15; 
Rst = 1'b0; 
cpu_addr = 32'd126;
  v_values_base = 32'd2; 
  wdata_col_base = 32'd6870 ; 
  csize = COL_SIZE; 
 fe_init = 1'b1; 
#15 Rst = 1'b1; 
// RD = 1'b0; 
// RD = 1'b1; 
 #518000; 
$finish; 
end 
always @(*) begin 
//$display("%b,%b",t1.fe1.count,t1.fe1.vdata_req); 
case(addr1)  
32'd6870: dataIn1 = 32'd1
; 
32'd6871: dataIn1 = 32'd4
; 
32'd6872: dataIn1 = 32'd5
; 
32'd6873: dataIn1 = 32'd10
; 
32'd6874: dataIn1 = 32'd2
; 
32'd6875: dataIn1 = 32'd3
; 
32'd6876: dataIn1 = 32'd7
; 
32'd6877: dataIn1 = 32'd161
; 
32'd6878: dataIn1 = 32'd3
; 
32'd6879: dataIn1 = 32'd6
; 
32'd6880: dataIn1 = 32'd9
; 
32'd6881: dataIn1 = 32'd4
; 
32'd6882: dataIn1 = 32'd12
; 
32'd6883: dataIn1 = 32'd185
; 
32'd6884: dataIn1 = 32'd5
; 
32'd6885: dataIn1 = 32'd6
; 
32'd6886: dataIn1 = 32'd7
; 
32'd6887: dataIn1 = 32'd10
; 
32'd6888: dataIn1 = 32'd217
; 
32'd6889: dataIn1 = 32'd8
; 
32'd6890: dataIn1 = 32'd9
; 
32'd6891: dataIn1 = 32'd217
; 
32'd6892: dataIn1 = 32'd229
; 
32'd6893: dataIn1 = 32'd9
; 
32'd6894: dataIn1 = 32'd10
; 
32'd6895: dataIn1 = 32'd11
; 
32'd6896: dataIn1 = 32'd11
; 
32'd6897: dataIn1 = 32'd186
; 
32'd6898: dataIn1 = 32'd12
; 
32'd6899: dataIn1 = 32'd13
; 
32'd6900: dataIn1 = 32'd17
; 
32'd6901: dataIn1 = 32'd53
; 
32'd6902: dataIn1 = 32'd176
; 
32'd6903: dataIn1 = 32'd13
; 
32'd6904: dataIn1 = 32'd15
; 
32'd6905: dataIn1 = 32'd176
; 
32'd6906: dataIn1 = 32'd14
; 
32'd6907: dataIn1 = 32'd17
; 
32'd6908: dataIn1 = 32'd19
; 
32'd6909: dataIn1 = 32'd160
; 
32'd6910: dataIn1 = 32'd15
; 
32'd6911: dataIn1 = 32'd22
; 
32'd6912: dataIn1 = 32'd16
; 
32'd6913: dataIn1 = 32'd162
; 
32'd6914: dataIn1 = 32'd178
; 
32'd6915: dataIn1 = 32'd17
; 
32'd6916: dataIn1 = 32'd18
; 
32'd6917: dataIn1 = 32'd19
; 
32'd6918: dataIn1 = 32'd18
; 
32'd6919: dataIn1 = 32'd19
; 
32'd6920: dataIn1 = 32'd19
; 
32'd6921: dataIn1 = 32'd53
; 
32'd6922: dataIn1 = 32'd55
; 
32'd6923: dataIn1 = 32'd20
; 
32'd6924: dataIn1 = 32'd22
; 
32'd6925: dataIn1 = 32'd124
; 
32'd6926: dataIn1 = 32'd178
; 
32'd6927: dataIn1 = 32'd21
; 
32'd6928: dataIn1 = 32'd22
; 
32'd6929: dataIn1 = 32'd23
; 
32'd6930: dataIn1 = 32'd137
; 
32'd6931: dataIn1 = 32'd178
; 
32'd6932: dataIn1 = 32'd22
; 
32'd6933: dataIn1 = 32'd23
; 
32'd6934: dataIn1 = 32'd125
; 
32'd6935: dataIn1 = 32'd24
; 
32'd6936: dataIn1 = 32'd48
; 
32'd6937: dataIn1 = 32'd50
; 
32'd6938: dataIn1 = 32'd51
; 
32'd6939: dataIn1 = 32'd25
; 
32'd6940: dataIn1 = 32'd27
; 
32'd6941: dataIn1 = 32'd28
; 
32'd6942: dataIn1 = 32'd163
; 
32'd6943: dataIn1 = 32'd26
; 
32'd6944: dataIn1 = 32'd43
; 
32'd6945: dataIn1 = 32'd189
; 
32'd6946: dataIn1 = 32'd208
; 
32'd6947: dataIn1 = 32'd27
; 
32'd6948: dataIn1 = 32'd43
; 
32'd6949: dataIn1 = 32'd182
; 
32'd6950: dataIn1 = 32'd28
; 
32'd6951: dataIn1 = 32'd43
; 
32'd6952: dataIn1 = 32'd182
; 
32'd6953: dataIn1 = 32'd189
; 
32'd6954: dataIn1 = 32'd29
; 
32'd6955: dataIn1 = 32'd30
; 
32'd6956: dataIn1 = 32'd46
; 
32'd6957: dataIn1 = 32'd30
; 
32'd6958: dataIn1 = 32'd31
; 
32'd6959: dataIn1 = 32'd32
; 
32'd6960: dataIn1 = 32'd189
; 
32'd6961: dataIn1 = 32'd31
; 
32'd6962: dataIn1 = 32'd35
; 
32'd6963: dataIn1 = 32'd32
; 
32'd6964: dataIn1 = 32'd52
; 
32'd6965: dataIn1 = 32'd33
; 
32'd6966: dataIn1 = 32'd35
; 
32'd6967: dataIn1 = 32'd47
; 
32'd6968: dataIn1 = 32'd183
; 
32'd6969: dataIn1 = 32'd34
; 
32'd6970: dataIn1 = 32'd46
; 
32'd6971: dataIn1 = 32'd47
; 
32'd6972: dataIn1 = 32'd35
; 
32'd6973: dataIn1 = 32'd36
; 
32'd6974: dataIn1 = 32'd38
; 
32'd6975: dataIn1 = 32'd175
; 
32'd6976: dataIn1 = 32'd37
; 
32'd6977: dataIn1 = 32'd38
; 
32'd6978: dataIn1 = 32'd211
; 
32'd6979: dataIn1 = 32'd38
; 
32'd6980: dataIn1 = 32'd40
; 
32'd6981: dataIn1 = 32'd58
; 
32'd6982: dataIn1 = 32'd39
; 
32'd6983: dataIn1 = 32'd40
; 
32'd6984: dataIn1 = 32'd40
; 
32'd6985: dataIn1 = 32'd41
; 
32'd6986: dataIn1 = 32'd541
; 
32'd6987: dataIn1 = 32'd41
; 
32'd6988: dataIn1 = 32'd42
; 
32'd6989: dataIn1 = 32'd173
; 
32'd6990: dataIn1 = 32'd43
; 
32'd6991: dataIn1 = 32'd46
; 
32'd6992: dataIn1 = 32'd189
; 
32'd6993: dataIn1 = 32'd44
; 
32'd6994: dataIn1 = 32'd45
; 
32'd6995: dataIn1 = 32'd47
; 
32'd6996: dataIn1 = 32'd49
; 
32'd6997: dataIn1 = 32'd51
; 
32'd6998: dataIn1 = 32'd45
; 
32'd6999: dataIn1 = 32'd46
; 
32'd7000: dataIn1 = 32'd47
; 
32'd7001: dataIn1 = 32'd52
; 
32'd7002: dataIn1 = 32'd182
; 
32'd7003: dataIn1 = 32'd46
; 
32'd7004: dataIn1 = 32'd157
; 
32'd7005: dataIn1 = 32'd47
; 
32'd7006: dataIn1 = 32'd48
; 
32'd7007: dataIn1 = 32'd49
; 
32'd7008: dataIn1 = 32'd50
; 
32'd7009: dataIn1 = 32'd49
; 
32'd7010: dataIn1 = 32'd50
; 
32'd7011: dataIn1 = 32'd182
; 
32'd7012: dataIn1 = 32'd50
; 
32'd7013: dataIn1 = 32'd51
; 
32'd7014: dataIn1 = 32'd52
; 
32'd7015: dataIn1 = 32'd53
; 
32'd7016: dataIn1 = 32'd54
; 
32'd7017: dataIn1 = 32'd54
; 
32'd7018: dataIn1 = 32'd55
; 
32'd7019: dataIn1 = 32'd185
; 
32'd7020: dataIn1 = 32'd55
; 
32'd7021: dataIn1 = 32'd56
; 
32'd7022: dataIn1 = 32'd60
; 
32'd7023: dataIn1 = 32'd61
; 
32'd7024: dataIn1 = 32'd189
; 
32'd7025: dataIn1 = 32'd57
; 
32'd7026: dataIn1 = 32'd61
; 
32'd7027: dataIn1 = 32'd190
; 
32'd7028: dataIn1 = 32'd58
; 
32'd7029: dataIn1 = 32'd59
; 
32'd7030: dataIn1 = 32'd59
; 
32'd7031: dataIn1 = 32'd61
; 
32'd7032: dataIn1 = 32'd60
; 
32'd7033: dataIn1 = 32'd211
; 
32'd7034: dataIn1 = 32'd61
; 
32'd7035: dataIn1 = 32'd62
; 
32'd7036: dataIn1 = 32'd64
; 
32'd7037: dataIn1 = 32'd67
; 
32'd7038: dataIn1 = 32'd63
; 
32'd7039: dataIn1 = 32'd64
; 
32'd7040: dataIn1 = 32'd65
; 
32'd7041: dataIn1 = 32'd66
; 
32'd7042: dataIn1 = 32'd64
; 
32'd7043: dataIn1 = 32'd65
; 
32'd7044: dataIn1 = 32'd67
; 
32'd7045: dataIn1 = 32'd184
; 
32'd7046: dataIn1 = 32'd65
; 
32'd7047: dataIn1 = 32'd66
; 
32'd7048: dataIn1 = 32'd616
; 
32'd7049: dataIn1 = 32'd67
; 
32'd7050: dataIn1 = 32'd68
; 
32'd7051: dataIn1 = 32'd88
; 
32'd7052: dataIn1 = 32'd90
; 
32'd7053: dataIn1 = 32'd94
; 
32'd7054: dataIn1 = 32'd69
; 
32'd7055: dataIn1 = 32'd70
; 
32'd7056: dataIn1 = 32'd71
; 
32'd7057: dataIn1 = 32'd74
; 
32'd7058: dataIn1 = 32'd91
; 
32'd7059: dataIn1 = 32'd103
; 
32'd7060: dataIn1 = 32'd70
; 
32'd7061: dataIn1 = 32'd93
; 
32'd7062: dataIn1 = 32'd98
; 
32'd7063: dataIn1 = 32'd126
; 
32'd7064: dataIn1 = 32'd129
; 
32'd7065: dataIn1 = 32'd143
; 
32'd7066: dataIn1 = 32'd171
; 
32'd7067: dataIn1 = 32'd207
; 
32'd7068: dataIn1 = 32'd71
; 
32'd7069: dataIn1 = 32'd91
; 
32'd7070: dataIn1 = 32'd96
; 
32'd7071: dataIn1 = 32'd97
; 
32'd7072: dataIn1 = 32'd106
; 
32'd7073: dataIn1 = 32'd72
; 
32'd7074: dataIn1 = 32'd75
; 
32'd7075: dataIn1 = 32'd107
; 
32'd7076: dataIn1 = 32'd152
; 
32'd7077: dataIn1 = 32'd73
; 
32'd7078: dataIn1 = 32'd81
; 
32'd7079: dataIn1 = 32'd83
; 
32'd7080: dataIn1 = 32'd89
; 
32'd7081: dataIn1 = 32'd74
; 
32'd7082: dataIn1 = 32'd78
; 
32'd7083: dataIn1 = 32'd80
; 
32'd7084: dataIn1 = 32'd75
; 
32'd7085: dataIn1 = 32'd103
; 
32'd7086: dataIn1 = 32'd107
; 
32'd7087: dataIn1 = 32'd123
; 
32'd7088: dataIn1 = 32'd127
; 
32'd7089: dataIn1 = 32'd76
; 
32'd7090: dataIn1 = 32'd101
; 
32'd7091: dataIn1 = 32'd131
; 
32'd7092: dataIn1 = 32'd153
; 
32'd7093: dataIn1 = 32'd77
; 
32'd7094: dataIn1 = 32'd95
; 
32'd7095: dataIn1 = 32'd117
; 
32'd7096: dataIn1 = 32'd132
; 
32'd7097: dataIn1 = 32'd158
; 
32'd7098: dataIn1 = 32'd78
; 
32'd7099: dataIn1 = 32'd85
; 
32'd7100: dataIn1 = 32'd96
; 
32'd7101: dataIn1 = 32'd97
; 
32'd7102: dataIn1 = 32'd106
; 
32'd7103: dataIn1 = 32'd79
; 
32'd7104: dataIn1 = 32'd81
; 
32'd7105: dataIn1 = 32'd84
; 
32'd7106: dataIn1 = 32'd88
; 
32'd7107: dataIn1 = 32'd117
; 
32'd7108: dataIn1 = 32'd151
; 
32'd7109: dataIn1 = 32'd80
; 
32'd7110: dataIn1 = 32'd82
; 
32'd7111: dataIn1 = 32'd85
; 
32'd7112: dataIn1 = 32'd97
; 
32'd7113: dataIn1 = 32'd101
; 
32'd7114: dataIn1 = 32'd81
; 
32'd7115: dataIn1 = 32'd83
; 
32'd7116: dataIn1 = 32'd148
; 
32'd7117: dataIn1 = 32'd151
; 
32'd7118: dataIn1 = 32'd82
; 
32'd7119: dataIn1 = 32'd96
; 
32'd7120: dataIn1 = 32'd101
; 
32'd7121: dataIn1 = 32'd83
; 
32'd7122: dataIn1 = 32'd103
; 
32'd7123: dataIn1 = 32'd127
; 
32'd7124: dataIn1 = 32'd149
; 
32'd7125: dataIn1 = 32'd84
; 
32'd7126: dataIn1 = 32'd86
; 
32'd7127: dataIn1 = 32'd99
; 
32'd7128: dataIn1 = 32'd104
; 
32'd7129: dataIn1 = 32'd148
; 
32'd7130: dataIn1 = 32'd85
; 
32'd7131: dataIn1 = 32'd97
; 
32'd7132: dataIn1 = 32'd106
; 
32'd7133: dataIn1 = 32'd146
; 
32'd7134: dataIn1 = 32'd86
; 
32'd7135: dataIn1 = 32'd87
; 
32'd7136: dataIn1 = 32'd88
; 
32'd7137: dataIn1 = 32'd87
; 
32'd7138: dataIn1 = 32'd99
; 
32'd7139: dataIn1 = 32'd102
; 
32'd7140: dataIn1 = 32'd105
; 
32'd7141: dataIn1 = 32'd110
; 
32'd7142: dataIn1 = 32'd111
; 
32'd7143: dataIn1 = 32'd148
; 
32'd7144: dataIn1 = 32'd149
; 
32'd7145: dataIn1 = 32'd88
; 
32'd7146: dataIn1 = 32'd95
; 
32'd7147: dataIn1 = 32'd102
; 
32'd7148: dataIn1 = 32'd89
; 
32'd7149: dataIn1 = 32'd92
; 
32'd7150: dataIn1 = 32'd96
; 
32'd7151: dataIn1 = 32'd90
; 
32'd7152: dataIn1 = 32'd131
; 
32'd7153: dataIn1 = 32'd158
; 
32'd7154: dataIn1 = 32'd159
; 
32'd7155: dataIn1 = 32'd91
; 
32'd7156: dataIn1 = 32'd144
; 
32'd7157: dataIn1 = 32'd92
; 
32'd7158: dataIn1 = 32'd117
; 
32'd7159: dataIn1 = 32'd146
; 
32'd7160: dataIn1 = 32'd93
; 
32'd7161: dataIn1 = 32'd98
; 
32'd7162: dataIn1 = 32'd177
; 
32'd7163: dataIn1 = 32'd193
; 
32'd7164: dataIn1 = 32'd94
; 
32'd7165: dataIn1 = 32'd131
; 
32'd7166: dataIn1 = 32'd154
; 
32'd7167: dataIn1 = 32'd95
; 
32'd7168: dataIn1 = 32'd104
; 
32'd7169: dataIn1 = 32'd105
; 
32'd7170: dataIn1 = 32'd117
; 
32'd7171: dataIn1 = 32'd151
; 
32'd7172: dataIn1 = 32'd159
; 
32'd7173: dataIn1 = 32'd96
; 
32'd7174: dataIn1 = 32'd146
; 
32'd7175: dataIn1 = 32'd97
; 
32'd7176: dataIn1 = 32'd98
; 
32'd7177: dataIn1 = 32'd106
; 
32'd7178: dataIn1 = 32'd98
; 
32'd7179: dataIn1 = 32'd128
; 
32'd7180: dataIn1 = 32'd129
; 
32'd7181: dataIn1 = 32'd99
; 
32'd7182: dataIn1 = 32'd100
; 
32'd7183: dataIn1 = 32'd102
; 
32'd7184: dataIn1 = 32'd105
; 
32'd7185: dataIn1 = 32'd100
; 
32'd7186: dataIn1 = 32'd118
; 
32'd7187: dataIn1 = 32'd134
; 
32'd7188: dataIn1 = 32'd142
; 
32'd7189: dataIn1 = 32'd147
; 
32'd7190: dataIn1 = 32'd101
; 
32'd7191: dataIn1 = 32'd102
; 
32'd7192: dataIn1 = 32'd110
; 
32'd7193: dataIn1 = 32'd111
; 
32'd7194: dataIn1 = 32'd136
; 
32'd7195: dataIn1 = 32'd103
; 
32'd7196: dataIn1 = 32'd144
; 
32'd7197: dataIn1 = 32'd152
; 
32'd7198: dataIn1 = 32'd104
; 
32'd7199: dataIn1 = 32'd151
; 
32'd7200: dataIn1 = 32'd105
; 
32'd7201: dataIn1 = 32'd132
; 
32'd7202: dataIn1 = 32'd106
; 
32'd7203: dataIn1 = 32'd107
; 
32'd7204: dataIn1 = 32'd108
; 
32'd7205: dataIn1 = 32'd115
; 
32'd7206: dataIn1 = 32'd123
; 
32'd7207: dataIn1 = 32'd108
; 
32'd7208: dataIn1 = 32'd114
; 
32'd7209: dataIn1 = 32'd115
; 
32'd7210: dataIn1 = 32'd121
; 
32'd7211: dataIn1 = 32'd123
; 
32'd7212: dataIn1 = 32'd124
; 
32'd7213: dataIn1 = 32'd109
; 
32'd7214: dataIn1 = 32'd111
; 
32'd7215: dataIn1 = 32'd115
; 
32'd7216: dataIn1 = 32'd116
; 
32'd7217: dataIn1 = 32'd123
; 
32'd7218: dataIn1 = 32'd110
; 
32'd7219: dataIn1 = 32'd111
; 
32'd7220: dataIn1 = 32'd113
; 
32'd7221: dataIn1 = 32'd136
; 
32'd7222: dataIn1 = 32'd140
; 
32'd7223: dataIn1 = 32'd111
; 
32'd7224: dataIn1 = 32'd112
; 
32'd7225: dataIn1 = 32'd113
; 
32'd7226: dataIn1 = 32'd116
; 
32'd7227: dataIn1 = 32'd120
; 
32'd7228: dataIn1 = 32'd138
; 
32'd7229: dataIn1 = 32'd140
; 
32'd7230: dataIn1 = 32'd141
; 
32'd7231: dataIn1 = 32'd112
; 
32'd7232: dataIn1 = 32'd113
; 
32'd7233: dataIn1 = 32'd134
; 
32'd7234: dataIn1 = 32'd136
; 
32'd7235: dataIn1 = 32'd113
; 
32'd7236: dataIn1 = 32'd116
; 
32'd7237: dataIn1 = 32'd122
; 
32'd7238: dataIn1 = 32'd133
; 
32'd7239: dataIn1 = 32'd134
; 
32'd7240: dataIn1 = 32'd135
; 
32'd7241: dataIn1 = 32'd138
; 
32'd7242: dataIn1 = 32'd140
; 
32'd7243: dataIn1 = 32'd114
; 
32'd7244: dataIn1 = 32'd115
; 
32'd7245: dataIn1 = 32'd122
; 
32'd7246: dataIn1 = 32'd135
; 
32'd7247: dataIn1 = 32'd139
; 
32'd7248: dataIn1 = 32'd115
; 
32'd7249: dataIn1 = 32'd116
; 
32'd7250: dataIn1 = 32'd119
; 
32'd7251: dataIn1 = 32'd121
; 
32'd7252: dataIn1 = 32'd123
; 
32'd7253: dataIn1 = 32'd124
; 
32'd7254: dataIn1 = 32'd116
; 
32'd7255: dataIn1 = 32'd123
; 
32'd7256: dataIn1 = 32'd138
; 
32'd7257: dataIn1 = 32'd140
; 
32'd7258: dataIn1 = 32'd117
; 
32'd7259: dataIn1 = 32'd118
; 
32'd7260: dataIn1 = 32'd132
; 
32'd7261: dataIn1 = 32'd118
; 
32'd7262: dataIn1 = 32'd145
; 
32'd7263: dataIn1 = 32'd150
; 
32'd7264: dataIn1 = 32'd155
; 
32'd7265: dataIn1 = 32'd119
; 
32'd7266: dataIn1 = 32'd120
; 
32'd7267: dataIn1 = 32'd123
; 
32'd7268: dataIn1 = 32'd125
; 
32'd7269: dataIn1 = 32'd126
; 
32'd7270: dataIn1 = 32'd137
; 
32'd7271: dataIn1 = 32'd141
; 
32'd7272: dataIn1 = 32'd143
; 
32'd7273: dataIn1 = 32'd120
; 
32'd7274: dataIn1 = 32'd150
; 
32'd7275: dataIn1 = 32'd121
; 
32'd7276: dataIn1 = 32'd125
; 
32'd7277: dataIn1 = 32'd122
; 
32'd7278: dataIn1 = 32'd135
; 
32'd7279: dataIn1 = 32'd139
; 
32'd7280: dataIn1 = 32'd140
; 
32'd7281: dataIn1 = 32'd123
; 
32'd7282: dataIn1 = 32'd124
; 
32'd7283: dataIn1 = 32'd125
; 
32'd7284: dataIn1 = 32'd126
; 
32'd7285: dataIn1 = 32'd127
; 
32'd7286: dataIn1 = 32'd127
; 
32'd7287: dataIn1 = 32'd152
; 
32'd7288: dataIn1 = 32'd128
; 
32'd7289: dataIn1 = 32'd129
; 
32'd7290: dataIn1 = 32'd153
; 
32'd7291: dataIn1 = 32'd129
; 
32'd7292: dataIn1 = 32'd145
; 
32'd7293: dataIn1 = 32'd147
; 
32'd7294: dataIn1 = 32'd130
; 
32'd7295: dataIn1 = 32'd131
; 
32'd7296: dataIn1 = 32'd153
; 
32'd7297: dataIn1 = 32'd155
; 
32'd7298: dataIn1 = 32'd131
; 
32'd7299: dataIn1 = 32'd154
; 
32'd7300: dataIn1 = 32'd132
; 
32'd7301: dataIn1 = 32'd133
; 
32'd7302: dataIn1 = 32'd134
; 
32'd7303: dataIn1 = 32'd138
; 
32'd7304: dataIn1 = 32'd134
; 
32'd7305: dataIn1 = 32'd140
; 
32'd7306: dataIn1 = 32'd135
; 
32'd7307: dataIn1 = 32'd138
; 
32'd7308: dataIn1 = 32'd139
; 
32'd7309: dataIn1 = 32'd136
; 
32'd7310: dataIn1 = 32'd137
; 
32'd7311: dataIn1 = 32'd138
; 
32'd7312: dataIn1 = 32'd140
; 
32'd7313: dataIn1 = 32'd139
; 
32'd7314: dataIn1 = 32'd140
; 
32'd7315: dataIn1 = 32'd140
; 
32'd7316: dataIn1 = 32'd141
; 
32'd7317: dataIn1 = 32'd142
; 
32'd7318: dataIn1 = 32'd150
; 
32'd7319: dataIn1 = 32'd143
; 
32'd7320: dataIn1 = 32'd144
; 
32'd7321: dataIn1 = 32'd144
; 
32'd7322: dataIn1 = 32'd145
; 
32'd7323: dataIn1 = 32'd146
; 
32'd7324: dataIn1 = 32'd146
; 
32'd7325: dataIn1 = 32'd147
; 
32'd7326: dataIn1 = 32'd148
; 
32'd7327: dataIn1 = 32'd148
; 
32'd7328: dataIn1 = 32'd149
; 
32'd7329: dataIn1 = 32'd149
; 
32'd7330: dataIn1 = 32'd150
; 
32'd7331: dataIn1 = 32'd151
; 
32'd7332: dataIn1 = 32'd151
; 
32'd7333: dataIn1 = 32'd152
; 
32'd7334: dataIn1 = 32'd153
; 
32'd7335: dataIn1 = 32'd154
; 
32'd7336: dataIn1 = 32'd155
; 
32'd7337: dataIn1 = 32'd156
; 
32'd7338: dataIn1 = 32'd156
; 
32'd7339: dataIn1 = 32'd158
; 
32'd7340: dataIn1 = 32'd159
; 
32'd7341: dataIn1 = 32'd157
; 
32'd7342: dataIn1 = 32'd158
; 
32'd7343: dataIn1 = 32'd159
; 
32'd7344: dataIn1 = 32'd160
; 
32'd7345: dataIn1 = 32'd185
; 
32'd7346: dataIn1 = 32'd161
; 
32'd7347: dataIn1 = 32'd205
; 
32'd7348: dataIn1 = 32'd162
; 
32'd7349: dataIn1 = 32'd188
; 
32'd7350: dataIn1 = 32'd163
; 
32'd7351: dataIn1 = 32'd164
; 
32'd7352: dataIn1 = 32'd165
; 
32'd7353: dataIn1 = 32'd188
; 
32'd7354: dataIn1 = 32'd203
; 
32'd7355: dataIn1 = 32'd164
; 
32'd7356: dataIn1 = 32'd165
; 
32'd7357: dataIn1 = 32'd201
; 
32'd7358: dataIn1 = 32'd166
; 
32'd7359: dataIn1 = 32'd167
; 
32'd7360: dataIn1 = 32'd219
; 
32'd7361: dataIn1 = 32'd167
; 
32'd7362: dataIn1 = 32'd194
; 
32'd7363: dataIn1 = 32'd195
; 
32'd7364: dataIn1 = 32'd168
; 
32'd7365: dataIn1 = 32'd178
; 
32'd7366: dataIn1 = 32'd183
; 
32'd7367: dataIn1 = 32'd169
; 
32'd7368: dataIn1 = 32'd170
; 
32'd7369: dataIn1 = 32'd171
; 
32'd7370: dataIn1 = 32'd172
; 
32'd7371: dataIn1 = 32'd216
; 
32'd7372: dataIn1 = 32'd170
; 
32'd7373: dataIn1 = 32'd189
; 
32'd7374: dataIn1 = 32'd211
; 
32'd7375: dataIn1 = 32'd171
; 
32'd7376: dataIn1 = 32'd184
; 
32'd7377: dataIn1 = 32'd193
; 
32'd7378: dataIn1 = 32'd210
; 
32'd7379: dataIn1 = 32'd172
; 
32'd7380: dataIn1 = 32'd173
; 
32'd7381: dataIn1 = 32'd174
; 
32'd7382: dataIn1 = 32'd184
; 
32'd7383: dataIn1 = 32'd193
; 
32'd7384: dataIn1 = 32'd628
; 
32'd7385: dataIn1 = 32'd631
; 
32'd7386: dataIn1 = 32'd173
; 
32'd7387: dataIn1 = 32'd174
; 
32'd7388: dataIn1 = 32'd175
; 
32'd7389: dataIn1 = 32'd190
; 
32'd7390: dataIn1 = 32'd174
; 
32'd7391: dataIn1 = 32'd175
; 
32'd7392: dataIn1 = 32'd190
; 
32'd7393: dataIn1 = 32'd667
; 
32'd7394: dataIn1 = 32'd176
; 
32'd7395: dataIn1 = 32'd177
; 
32'd7396: dataIn1 = 32'd193
; 
32'd7397: dataIn1 = 32'd178
; 
32'd7398: dataIn1 = 32'd179
; 
32'd7399: dataIn1 = 32'd180
; 
32'd7400: dataIn1 = 32'd208
; 
32'd7401: dataIn1 = 32'd180
; 
32'd7402: dataIn1 = 32'd184
; 
32'd7403: dataIn1 = 32'd192
; 
32'd7404: dataIn1 = 32'd212
; 
32'd7405: dataIn1 = 32'd626
; 
32'd7406: dataIn1 = 32'd181
; 
32'd7407: dataIn1 = 32'd188
; 
32'd7408: dataIn1 = 32'd215
; 
32'd7409: dataIn1 = 32'd182
; 
32'd7410: dataIn1 = 32'd204
; 
32'd7411: dataIn1 = 32'd183
; 
32'd7412: dataIn1 = 32'd215
; 
32'd7413: dataIn1 = 32'd184
; 
32'd7414: dataIn1 = 32'd185
; 
32'd7415: dataIn1 = 32'd188
; 
32'd7416: dataIn1 = 32'd206
; 
32'd7417: dataIn1 = 32'd186
; 
32'd7418: dataIn1 = 32'd205
; 
32'd7419: dataIn1 = 32'd213
; 
32'd7420: dataIn1 = 32'd187
; 
32'd7421: dataIn1 = 32'd194
; 
32'd7422: dataIn1 = 32'd188
; 
32'd7423: dataIn1 = 32'd191
; 
32'd7424: dataIn1 = 32'd189
; 
32'd7425: dataIn1 = 32'd190
; 
32'd7426: dataIn1 = 32'd518
; 
32'd7427: dataIn1 = 32'd191
; 
32'd7428: dataIn1 = 32'd205
; 
32'd7429: dataIn1 = 32'd206
; 
32'd7430: dataIn1 = 32'd192
; 
32'd7431: dataIn1 = 32'd193
; 
32'd7432: dataIn1 = 32'd193
; 
32'd7433: dataIn1 = 32'd210
; 
32'd7434: dataIn1 = 32'd214
; 
32'd7435: dataIn1 = 32'd194
; 
32'd7436: dataIn1 = 32'd196
; 
32'd7437: dataIn1 = 32'd195
; 
32'd7438: dataIn1 = 32'd203
; 
32'd7439: dataIn1 = 32'd196
; 
32'd7440: dataIn1 = 32'd197
; 
32'd7441: dataIn1 = 32'd198
; 
32'd7442: dataIn1 = 32'd685
; 
32'd7443: dataIn1 = 32'd197
; 
32'd7444: dataIn1 = 32'd290
; 
32'd7445: dataIn1 = 32'd198
; 
32'd7446: dataIn1 = 32'd199
; 
32'd7447: dataIn1 = 32'd200
; 
32'd7448: dataIn1 = 32'd199
; 
32'd7449: dataIn1 = 32'd421
; 
32'd7450: dataIn1 = 32'd200
; 
32'd7451: dataIn1 = 32'd201
; 
32'd7452: dataIn1 = 32'd204
; 
32'd7453: dataIn1 = 32'd201
; 
32'd7454: dataIn1 = 32'd202
; 
32'd7455: dataIn1 = 32'd203
; 
32'd7456: dataIn1 = 32'd209
; 
32'd7457: dataIn1 = 32'd213
; 
32'd7458: dataIn1 = 32'd203
; 
32'd7459: dataIn1 = 32'd204
; 
32'd7460: dataIn1 = 32'd205
; 
32'd7461: dataIn1 = 32'd212
; 
32'd7462: dataIn1 = 32'd206
; 
32'd7463: dataIn1 = 32'd207
; 
32'd7464: dataIn1 = 32'd214
; 
32'd7465: dataIn1 = 32'd215
; 
32'd7466: dataIn1 = 32'd216
; 
32'd7467: dataIn1 = 32'd208
; 
32'd7468: dataIn1 = 32'd209
; 
32'd7469: dataIn1 = 32'd210
; 
32'd7470: dataIn1 = 32'd211
; 
32'd7471: dataIn1 = 32'd212
; 
32'd7472: dataIn1 = 32'd213
; 
32'd7473: dataIn1 = 32'd215
; 
32'd7474: dataIn1 = 32'd213
; 
32'd7475: dataIn1 = 32'd214
; 
32'd7476: dataIn1 = 32'd215
; 
32'd7477: dataIn1 = 32'd216
; 
32'd7478: dataIn1 = 32'd217
; 
32'd7479: dataIn1 = 32'd218
; 
32'd7480: dataIn1 = 32'd268
; 
32'd7481: dataIn1 = 32'd218
; 
32'd7482: dataIn1 = 32'd219
; 
32'd7483: dataIn1 = 32'd220
; 
32'd7484: dataIn1 = 32'd237
; 
32'd7485: dataIn1 = 32'd671
; 
32'd7486: dataIn1 = 32'd672
; 
32'd7487: dataIn1 = 32'd219
; 
32'd7488: dataIn1 = 32'd672
; 
32'd7489: dataIn1 = 32'd220
; 
32'd7490: dataIn1 = 32'd267
; 
32'd7491: dataIn1 = 32'd670
; 
32'd7492: dataIn1 = 32'd671
; 
32'd7493: dataIn1 = 32'd221
; 
32'd7494: dataIn1 = 32'd233
; 
32'd7495: dataIn1 = 32'd235
; 
32'd7496: dataIn1 = 32'd236
; 
32'd7497: dataIn1 = 32'd222
; 
32'd7498: dataIn1 = 32'd256
; 
32'd7499: dataIn1 = 32'd223
; 
32'd7500: dataIn1 = 32'd224
; 
32'd7501: dataIn1 = 32'd226
; 
32'd7502: dataIn1 = 32'd265
; 
32'd7503: dataIn1 = 32'd673
; 
32'd7504: dataIn1 = 32'd224
; 
32'd7505: dataIn1 = 32'd225
; 
32'd7506: dataIn1 = 32'd225
; 
32'd7507: dataIn1 = 32'd229
; 
32'd7508: dataIn1 = 32'd265
; 
32'd7509: dataIn1 = 32'd266
; 
32'd7510: dataIn1 = 32'd673
; 
32'd7511: dataIn1 = 32'd226
; 
32'd7512: dataIn1 = 32'd227
; 
32'd7513: dataIn1 = 32'd228
; 
32'd7514: dataIn1 = 32'd230
; 
32'd7515: dataIn1 = 32'd673
; 
32'd7516: dataIn1 = 32'd227
; 
32'd7517: dataIn1 = 32'd231
; 
32'd7518: dataIn1 = 32'd232
; 
32'd7519: dataIn1 = 32'd233
; 
32'd7520: dataIn1 = 32'd228
; 
32'd7521: dataIn1 = 32'd236
; 
32'd7522: dataIn1 = 32'd266
; 
32'd7523: dataIn1 = 32'd229
; 
32'd7524: dataIn1 = 32'd256
; 
32'd7525: dataIn1 = 32'd265
; 
32'd7526: dataIn1 = 32'd266
; 
32'd7527: dataIn1 = 32'd268
; 
32'd7528: dataIn1 = 32'd230
; 
32'd7529: dataIn1 = 32'd231
; 
32'd7530: dataIn1 = 32'd232
; 
32'd7531: dataIn1 = 32'd234
; 
32'd7532: dataIn1 = 32'd235
; 
32'd7533: dataIn1 = 32'd236
; 
32'd7534: dataIn1 = 32'd256
; 
32'd7535: dataIn1 = 32'd265
; 
32'd7536: dataIn1 = 32'd231
; 
32'd7537: dataIn1 = 32'd232
; 
32'd7538: dataIn1 = 32'd233
; 
32'd7539: dataIn1 = 32'd234
; 
32'd7540: dataIn1 = 32'd234
; 
32'd7541: dataIn1 = 32'd235
; 
32'd7542: dataIn1 = 32'd236
; 
32'd7543: dataIn1 = 32'd253
; 
32'd7544: dataIn1 = 32'd237
; 
32'd7545: dataIn1 = 32'd238
; 
32'd7546: dataIn1 = 32'd252
; 
32'd7547: dataIn1 = 32'd269
; 
32'd7548: dataIn1 = 32'd238
; 
32'd7549: dataIn1 = 32'd239
; 
32'd7550: dataIn1 = 32'd240
; 
32'd7551: dataIn1 = 32'd253
; 
32'd7552: dataIn1 = 32'd261
; 
32'd7553: dataIn1 = 32'd239
; 
32'd7554: dataIn1 = 32'd240
; 
32'd7555: dataIn1 = 32'd241
; 
32'd7556: dataIn1 = 32'd242
; 
32'd7557: dataIn1 = 32'd253
; 
32'd7558: dataIn1 = 32'd261
; 
32'd7559: dataIn1 = 32'd675
; 
32'd7560: dataIn1 = 32'd240
; 
32'd7561: dataIn1 = 32'd241
; 
32'd7562: dataIn1 = 32'd261
; 
32'd7563: dataIn1 = 32'd262
; 
32'd7564: dataIn1 = 32'd675
; 
32'd7565: dataIn1 = 32'd241
; 
32'd7566: dataIn1 = 32'd243
; 
32'd7567: dataIn1 = 32'd253
; 
32'd7568: dataIn1 = 32'd259
; 
32'd7569: dataIn1 = 32'd262
; 
32'd7570: dataIn1 = 32'd675
; 
32'd7571: dataIn1 = 32'd677
; 
32'd7572: dataIn1 = 32'd242
; 
32'd7573: dataIn1 = 32'd264
; 
32'd7574: dataIn1 = 32'd674
; 
32'd7575: dataIn1 = 32'd243
; 
32'd7576: dataIn1 = 32'd246
; 
32'd7577: dataIn1 = 32'd255
; 
32'd7578: dataIn1 = 32'd679
; 
32'd7579: dataIn1 = 32'd680
; 
32'd7580: dataIn1 = 32'd244
; 
32'd7581: dataIn1 = 32'd245
; 
32'd7582: dataIn1 = 32'd676
; 
32'd7583: dataIn1 = 32'd678
; 
32'd7584: dataIn1 = 32'd245
; 
32'd7585: dataIn1 = 32'd261
; 
32'd7586: dataIn1 = 32'd676
; 
32'd7587: dataIn1 = 32'd677
; 
32'd7588: dataIn1 = 32'd678
; 
32'd7589: dataIn1 = 32'd246
; 
32'd7590: dataIn1 = 32'd247
; 
32'd7591: dataIn1 = 32'd254
; 
32'd7592: dataIn1 = 32'd255
; 
32'd7593: dataIn1 = 32'd676
; 
32'd7594: dataIn1 = 32'd679
; 
32'd7595: dataIn1 = 32'd680
; 
32'd7596: dataIn1 = 32'd247
; 
32'd7597: dataIn1 = 32'd248
; 
32'd7598: dataIn1 = 32'd255
; 
32'd7599: dataIn1 = 32'd259
; 
32'd7600: dataIn1 = 32'd680
; 
32'd7601: dataIn1 = 32'd681
; 
32'd7602: dataIn1 = 32'd248
; 
32'd7603: dataIn1 = 32'd254
; 
32'd7604: dataIn1 = 32'd249
; 
32'd7605: dataIn1 = 32'd259
; 
32'd7606: dataIn1 = 32'd684
; 
32'd7607: dataIn1 = 32'd250
; 
32'd7608: dataIn1 = 32'd251
; 
32'd7609: dataIn1 = 32'd255
; 
32'd7610: dataIn1 = 32'd251
; 
32'd7611: dataIn1 = 32'd255
; 
32'd7612: dataIn1 = 32'd252
; 
32'd7613: dataIn1 = 32'd256
; 
32'd7614: dataIn1 = 32'd260
; 
32'd7615: dataIn1 = 32'd253
; 
32'd7616: dataIn1 = 32'd268
; 
32'd7617: dataIn1 = 32'd677
; 
32'd7618: dataIn1 = 32'd254
; 
32'd7619: dataIn1 = 32'd258
; 
32'd7620: dataIn1 = 32'd269
; 
32'd7621: dataIn1 = 32'd255
; 
32'd7622: dataIn1 = 32'd679
; 
32'd7623: dataIn1 = 32'd680
; 
32'd7624: dataIn1 = 32'd683
; 
32'd7625: dataIn1 = 32'd256
; 
32'd7626: dataIn1 = 32'd257
; 
32'd7627: dataIn1 = 32'd258
; 
32'd7628: dataIn1 = 32'd258
; 
32'd7629: dataIn1 = 32'd259
; 
32'd7630: dataIn1 = 32'd259
; 
32'd7631: dataIn1 = 32'd684
; 
32'd7632: dataIn1 = 32'd260
; 
32'd7633: dataIn1 = 32'd263
; 
32'd7634: dataIn1 = 32'd268
; 
32'd7635: dataIn1 = 32'd669
; 
32'd7636: dataIn1 = 32'd261
; 
32'd7637: dataIn1 = 32'd262
; 
32'd7638: dataIn1 = 32'd262
; 
32'd7639: dataIn1 = 32'd264
; 
32'd7640: dataIn1 = 32'd675
; 
32'd7641: dataIn1 = 32'd677
; 
32'd7642: dataIn1 = 32'd263
; 
32'd7643: dataIn1 = 32'd264
; 
32'd7644: dataIn1 = 32'd264
; 
32'd7645: dataIn1 = 32'd265
; 
32'd7646: dataIn1 = 32'd266
; 
32'd7647: dataIn1 = 32'd266
; 
32'd7648: dataIn1 = 32'd267
; 
32'd7649: dataIn1 = 32'd268
; 
32'd7650: dataIn1 = 32'd269
; 
32'd7651: dataIn1 = 32'd270
; 
32'd7652: dataIn1 = 32'd271
; 
32'd7653: dataIn1 = 32'd273
; 
32'd7654: dataIn1 = 32'd276
; 
32'd7655: dataIn1 = 32'd277
; 
32'd7656: dataIn1 = 32'd278
; 
32'd7657: dataIn1 = 32'd280
; 
32'd7658: dataIn1 = 32'd283
; 
32'd7659: dataIn1 = 32'd287
; 
32'd7660: dataIn1 = 32'd297
; 
32'd7661: dataIn1 = 32'd271
; 
32'd7662: dataIn1 = 32'd275
; 
32'd7663: dataIn1 = 32'd277
; 
32'd7664: dataIn1 = 32'd280
; 
32'd7665: dataIn1 = 32'd272
; 
32'd7666: dataIn1 = 32'd274
; 
32'd7667: dataIn1 = 32'd273
; 
32'd7668: dataIn1 = 32'd274
; 
32'd7669: dataIn1 = 32'd277
; 
32'd7670: dataIn1 = 32'd278
; 
32'd7671: dataIn1 = 32'd280
; 
32'd7672: dataIn1 = 32'd274
; 
32'd7673: dataIn1 = 32'd277
; 
32'd7674: dataIn1 = 32'd278
; 
32'd7675: dataIn1 = 32'd275
; 
32'd7676: dataIn1 = 32'd277
; 
32'd7677: dataIn1 = 32'd278
; 
32'd7678: dataIn1 = 32'd276
; 
32'd7679: dataIn1 = 32'd280
; 
32'd7680: dataIn1 = 32'd281
; 
32'd7681: dataIn1 = 32'd283
; 
32'd7682: dataIn1 = 32'd284
; 
32'd7683: dataIn1 = 32'd277
; 
32'd7684: dataIn1 = 32'd278
; 
32'd7685: dataIn1 = 32'd280
; 
32'd7686: dataIn1 = 32'd278
; 
32'd7687: dataIn1 = 32'd279
; 
32'd7688: dataIn1 = 32'd287
; 
32'd7689: dataIn1 = 32'd297
; 
32'd7690: dataIn1 = 32'd279
; 
32'd7691: dataIn1 = 32'd290
; 
32'd7692: dataIn1 = 32'd280
; 
32'd7693: dataIn1 = 32'd281
; 
32'd7694: dataIn1 = 32'd282
; 
32'd7695: dataIn1 = 32'd283
; 
32'd7696: dataIn1 = 32'd284
; 
32'd7697: dataIn1 = 32'd289
; 
32'd7698: dataIn1 = 32'd290
; 
32'd7699: dataIn1 = 32'd295
; 
32'd7700: dataIn1 = 32'd282
; 
32'd7701: dataIn1 = 32'd296
; 
32'd7702: dataIn1 = 32'd301
; 
32'd7703: dataIn1 = 32'd310
; 
32'd7704: dataIn1 = 32'd311
; 
32'd7705: dataIn1 = 32'd312
; 
32'd7706: dataIn1 = 32'd283
; 
32'd7707: dataIn1 = 32'd289
; 
32'd7708: dataIn1 = 32'd290
; 
32'd7709: dataIn1 = 32'd295
; 
32'd7710: dataIn1 = 32'd297
; 
32'd7711: dataIn1 = 32'd284
; 
32'd7712: dataIn1 = 32'd285
; 
32'd7713: dataIn1 = 32'd286
; 
32'd7714: dataIn1 = 32'd288
; 
32'd7715: dataIn1 = 32'd289
; 
32'd7716: dataIn1 = 32'd291
; 
32'd7717: dataIn1 = 32'd293
; 
32'd7718: dataIn1 = 32'd295
; 
32'd7719: dataIn1 = 32'd296
; 
32'd7720: dataIn1 = 32'd297
; 
32'd7721: dataIn1 = 32'd298
; 
32'd7722: dataIn1 = 32'd286
; 
32'd7723: dataIn1 = 32'd295
; 
32'd7724: dataIn1 = 32'd297
; 
32'd7725: dataIn1 = 32'd298
; 
32'd7726: dataIn1 = 32'd315
; 
32'd7727: dataIn1 = 32'd287
; 
32'd7728: dataIn1 = 32'd293
; 
32'd7729: dataIn1 = 32'd295
; 
32'd7730: dataIn1 = 32'd297
; 
32'd7731: dataIn1 = 32'd288
; 
32'd7732: dataIn1 = 32'd291
; 
32'd7733: dataIn1 = 32'd293
; 
32'd7734: dataIn1 = 32'd298
; 
32'd7735: dataIn1 = 32'd307
; 
32'd7736: dataIn1 = 32'd289
; 
32'd7737: dataIn1 = 32'd290
; 
32'd7738: dataIn1 = 32'd293
; 
32'd7739: dataIn1 = 32'd295
; 
32'd7740: dataIn1 = 32'd297
; 
32'd7741: dataIn1 = 32'd298
; 
32'd7742: dataIn1 = 32'd290
; 
32'd7743: dataIn1 = 32'd292
; 
32'd7744: dataIn1 = 32'd295
; 
32'd7745: dataIn1 = 32'd309
; 
32'd7746: dataIn1 = 32'd291
; 
32'd7747: dataIn1 = 32'd292
; 
32'd7748: dataIn1 = 32'd294
; 
32'd7749: dataIn1 = 32'd298
; 
32'd7750: dataIn1 = 32'd315
; 
32'd7751: dataIn1 = 32'd292
; 
32'd7752: dataIn1 = 32'd309
; 
32'd7753: dataIn1 = 32'd293
; 
32'd7754: dataIn1 = 32'd294
; 
32'd7755: dataIn1 = 32'd294
; 
32'd7756: dataIn1 = 32'd295
; 
32'd7757: dataIn1 = 32'd296
; 
32'd7758: dataIn1 = 32'd297
; 
32'd7759: dataIn1 = 32'd298
; 
32'd7760: dataIn1 = 32'd311
; 
32'd7761: dataIn1 = 32'd296
; 
32'd7762: dataIn1 = 32'd301
; 
32'd7763: dataIn1 = 32'd310
; 
32'd7764: dataIn1 = 32'd311
; 
32'd7765: dataIn1 = 32'd312
; 
32'd7766: dataIn1 = 32'd297
; 
32'd7767: dataIn1 = 32'd298
; 
32'd7768: dataIn1 = 32'd298
; 
32'd7769: dataIn1 = 32'd299
; 
32'd7770: dataIn1 = 32'd300
; 
32'd7771: dataIn1 = 32'd303
; 
32'd7772: dataIn1 = 32'd305
; 
32'd7773: dataIn1 = 32'd314
; 
32'd7774: dataIn1 = 32'd300
; 
32'd7775: dataIn1 = 32'd305
; 
32'd7776: dataIn1 = 32'd306
; 
32'd7777: dataIn1 = 32'd308
; 
32'd7778: dataIn1 = 32'd301
; 
32'd7779: dataIn1 = 32'd310
; 
32'd7780: dataIn1 = 32'd311
; 
32'd7781: dataIn1 = 32'd312
; 
32'd7782: dataIn1 = 32'd302
; 
32'd7783: dataIn1 = 32'd313
; 
32'd7784: dataIn1 = 32'd303
; 
32'd7785: dataIn1 = 32'd305
; 
32'd7786: dataIn1 = 32'd304
; 
32'd7787: dataIn1 = 32'd308
; 
32'd7788: dataIn1 = 32'd313
; 
32'd7789: dataIn1 = 32'd305
; 
32'd7790: dataIn1 = 32'd306
; 
32'd7791: dataIn1 = 32'd312
; 
32'd7792: dataIn1 = 32'd306
; 
32'd7793: dataIn1 = 32'd308
; 
32'd7794: dataIn1 = 32'd312
; 
32'd7795: dataIn1 = 32'd313
; 
32'd7796: dataIn1 = 32'd307
; 
32'd7797: dataIn1 = 32'd310
; 
32'd7798: dataIn1 = 32'd308
; 
32'd7799: dataIn1 = 32'd309
; 
32'd7800: dataIn1 = 32'd309
; 
32'd7801: dataIn1 = 32'd310
; 
32'd7802: dataIn1 = 32'd311
; 
32'd7803: dataIn1 = 32'd312
; 
32'd7804: dataIn1 = 32'd315
; 
32'd7805: dataIn1 = 32'd311
; 
32'd7806: dataIn1 = 32'd312
; 
32'd7807: dataIn1 = 32'd312
; 
32'd7808: dataIn1 = 32'd313
; 
32'd7809: dataIn1 = 32'd313
; 
32'd7810: dataIn1 = 32'd314
; 
32'd7811: dataIn1 = 32'd315
; 
32'd7812: dataIn1 = 32'd316
; 
32'd7813: dataIn1 = 32'd408
; 
32'd7814: dataIn1 = 32'd317
; 
32'd7815: dataIn1 = 32'd318
; 
32'd7816: dataIn1 = 32'd324
; 
32'd7817: dataIn1 = 32'd339
; 
32'd7818: dataIn1 = 32'd343
; 
32'd7819: dataIn1 = 32'd344
; 
32'd7820: dataIn1 = 32'd357
; 
32'd7821: dataIn1 = 32'd363
; 
32'd7822: dataIn1 = 32'd373
; 
32'd7823: dataIn1 = 32'd431
; 
32'd7824: dataIn1 = 32'd435
; 
32'd7825: dataIn1 = 32'd441
; 
32'd7826: dataIn1 = 32'd446
; 
32'd7827: dataIn1 = 32'd318
; 
32'd7828: dataIn1 = 32'd435
; 
32'd7829: dataIn1 = 32'd446
; 
32'd7830: dataIn1 = 32'd319
; 
32'd7831: dataIn1 = 32'd320
; 
32'd7832: dataIn1 = 32'd360
; 
32'd7833: dataIn1 = 32'd363
; 
32'd7834: dataIn1 = 32'd364
; 
32'd7835: dataIn1 = 32'd320
; 
32'd7836: dataIn1 = 32'd321
; 
32'd7837: dataIn1 = 32'd322
; 
32'd7838: dataIn1 = 32'd321
; 
32'd7839: dataIn1 = 32'd322
; 
32'd7840: dataIn1 = 32'd323
; 
32'd7841: dataIn1 = 32'd324
; 
32'd7842: dataIn1 = 32'd427
; 
32'd7843: dataIn1 = 32'd438
; 
32'd7844: dataIn1 = 32'd442
; 
32'd7845: dataIn1 = 32'd322
; 
32'd7846: dataIn1 = 32'd323
; 
32'd7847: dataIn1 = 32'd437
; 
32'd7848: dataIn1 = 32'd438
; 
32'd7849: dataIn1 = 32'd440
; 
32'd7850: dataIn1 = 32'd442
; 
32'd7851: dataIn1 = 32'd446
; 
32'd7852: dataIn1 = 32'd324
; 
32'd7853: dataIn1 = 32'd427
; 
32'd7854: dataIn1 = 32'd442
; 
32'd7855: dataIn1 = 32'd446
; 
32'd7856: dataIn1 = 32'd325
; 
32'd7857: dataIn1 = 32'd339
; 
32'd7858: dataIn1 = 32'd427
; 
32'd7859: dataIn1 = 32'd445
; 
32'd7860: dataIn1 = 32'd446
; 
32'd7861: dataIn1 = 32'd326
; 
32'd7862: dataIn1 = 32'd328
; 
32'd7863: dataIn1 = 32'd339
; 
32'd7864: dataIn1 = 32'd445
; 
32'd7865: dataIn1 = 32'd327
; 
32'd7866: dataIn1 = 32'd328
; 
32'd7867: dataIn1 = 32'd409
; 
32'd7868: dataIn1 = 32'd328
; 
32'd7869: dataIn1 = 32'd330
; 
32'd7870: dataIn1 = 32'd409
; 
32'd7871: dataIn1 = 32'd430
; 
32'd7872: dataIn1 = 32'd436
; 
32'd7873: dataIn1 = 32'd329
; 
32'd7874: dataIn1 = 32'd336
; 
32'd7875: dataIn1 = 32'd424
; 
32'd7876: dataIn1 = 32'd430
; 
32'd7877: dataIn1 = 32'd330
; 
32'd7878: dataIn1 = 32'd331
; 
32'd7879: dataIn1 = 32'd336
; 
32'd7880: dataIn1 = 32'd331
; 
32'd7881: dataIn1 = 32'd336
; 
32'd7882: dataIn1 = 32'd424
; 
32'd7883: dataIn1 = 32'd436
; 
32'd7884: dataIn1 = 32'd332
; 
32'd7885: dataIn1 = 32'd333
; 
32'd7886: dataIn1 = 32'd347
; 
32'd7887: dataIn1 = 32'd333
; 
32'd7888: dataIn1 = 32'd334
; 
32'd7889: dataIn1 = 32'd335
; 
32'd7890: dataIn1 = 32'd336
; 
32'd7891: dataIn1 = 32'd424
; 
32'd7892: dataIn1 = 32'd334
; 
32'd7893: dataIn1 = 32'd336
; 
32'd7894: dataIn1 = 32'd335
; 
32'd7895: dataIn1 = 32'd336
; 
32'd7896: dataIn1 = 32'd424
; 
32'd7897: dataIn1 = 32'd336
; 
32'd7898: dataIn1 = 32'd337
; 
32'd7899: dataIn1 = 32'd338
; 
32'd7900: dataIn1 = 32'd344
; 
32'd7901: dataIn1 = 32'd337
; 
32'd7902: dataIn1 = 32'd338
; 
32'd7903: dataIn1 = 32'd345
; 
32'd7904: dataIn1 = 32'd349
; 
32'd7905: dataIn1 = 32'd338
; 
32'd7906: dataIn1 = 32'd345
; 
32'd7907: dataIn1 = 32'd339
; 
32'd7908: dataIn1 = 32'd340
; 
32'd7909: dataIn1 = 32'd341
; 
32'd7910: dataIn1 = 32'd340
; 
32'd7911: dataIn1 = 32'd341
; 
32'd7912: dataIn1 = 32'd427
; 
32'd7913: dataIn1 = 32'd341
; 
32'd7914: dataIn1 = 32'd342
; 
32'd7915: dataIn1 = 32'd357
; 
32'd7916: dataIn1 = 32'd360
; 
32'd7917: dataIn1 = 32'd362
; 
32'd7918: dataIn1 = 32'd428
; 
32'd7919: dataIn1 = 32'd441
; 
32'd7920: dataIn1 = 32'd342
; 
32'd7921: dataIn1 = 32'd347
; 
32'd7922: dataIn1 = 32'd343
; 
32'd7923: dataIn1 = 32'd344
; 
32'd7924: dataIn1 = 32'd345
; 
32'd7925: dataIn1 = 32'd357
; 
32'd7926: dataIn1 = 32'd431
; 
32'd7927: dataIn1 = 32'd441
; 
32'd7928: dataIn1 = 32'd344
; 
32'd7929: dataIn1 = 32'd345
; 
32'd7930: dataIn1 = 32'd373
; 
32'd7931: dataIn1 = 32'd345
; 
32'd7932: dataIn1 = 32'd346
; 
32'd7933: dataIn1 = 32'd354
; 
32'd7934: dataIn1 = 32'd375
; 
32'd7935: dataIn1 = 32'd346
; 
32'd7936: dataIn1 = 32'd348
; 
32'd7937: dataIn1 = 32'd347
; 
32'd7938: dataIn1 = 32'd352
; 
32'd7939: dataIn1 = 32'd443
; 
32'd7940: dataIn1 = 32'd348
; 
32'd7941: dataIn1 = 32'd349
; 
32'd7942: dataIn1 = 32'd349
; 
32'd7943: dataIn1 = 32'd353
; 
32'd7944: dataIn1 = 32'd354
; 
32'd7945: dataIn1 = 32'd433
; 
32'd7946: dataIn1 = 32'd434
; 
32'd7947: dataIn1 = 32'd443
; 
32'd7948: dataIn1 = 32'd350
; 
32'd7949: dataIn1 = 32'd351
; 
32'd7950: dataIn1 = 32'd368
; 
32'd7951: dataIn1 = 32'd381
; 
32'd7952: dataIn1 = 32'd382
; 
32'd7953: dataIn1 = 32'd433
; 
32'd7954: dataIn1 = 32'd434
; 
32'd7955: dataIn1 = 32'd351
; 
32'd7956: dataIn1 = 32'd353
; 
32'd7957: dataIn1 = 32'd352
; 
32'd7958: dataIn1 = 32'd353
; 
32'd7959: dataIn1 = 32'd376
; 
32'd7960: dataIn1 = 32'd353
; 
32'd7961: dataIn1 = 32'd381
; 
32'd7962: dataIn1 = 32'd354
; 
32'd7963: dataIn1 = 32'd375
; 
32'd7964: dataIn1 = 32'd355
; 
32'd7965: dataIn1 = 32'd356
; 
32'd7966: dataIn1 = 32'd366
; 
32'd7967: dataIn1 = 32'd367
; 
32'd7968: dataIn1 = 32'd370
; 
32'd7969: dataIn1 = 32'd373
; 
32'd7970: dataIn1 = 32'd429
; 
32'd7971: dataIn1 = 32'd431
; 
32'd7972: dataIn1 = 32'd356
; 
32'd7973: dataIn1 = 32'd358
; 
32'd7974: dataIn1 = 32'd357
; 
32'd7975: dataIn1 = 32'd358
; 
32'd7976: dataIn1 = 32'd360
; 
32'd7977: dataIn1 = 32'd429
; 
32'd7978: dataIn1 = 32'd441
; 
32'd7979: dataIn1 = 32'd358
; 
32'd7980: dataIn1 = 32'd360
; 
32'd7981: dataIn1 = 32'd429
; 
32'd7982: dataIn1 = 32'd359
; 
32'd7983: dataIn1 = 32'd360
; 
32'd7984: dataIn1 = 32'd361
; 
32'd7985: dataIn1 = 32'd363
; 
32'd7986: dataIn1 = 32'd366
; 
32'd7987: dataIn1 = 32'd429
; 
32'd7988: dataIn1 = 32'd360
; 
32'd7989: dataIn1 = 32'd441
; 
32'd7990: dataIn1 = 32'd361
; 
32'd7991: dataIn1 = 32'd363
; 
32'd7992: dataIn1 = 32'd362
; 
32'd7993: dataIn1 = 32'd363
; 
32'd7994: dataIn1 = 32'd364
; 
32'd7995: dataIn1 = 32'd364
; 
32'd7996: dataIn1 = 32'd365
; 
32'd7997: dataIn1 = 32'd365
; 
32'd7998: dataIn1 = 32'd399
; 
32'd7999: dataIn1 = 32'd366
; 
32'd8000: dataIn1 = 32'd367
; 
32'd8001: dataIn1 = 32'd402
; 
32'd8002: dataIn1 = 32'd429
; 
32'd8003: dataIn1 = 32'd367
; 
32'd8004: dataIn1 = 32'd369
; 
32'd8005: dataIn1 = 32'd402
; 
32'd8006: dataIn1 = 32'd404
; 
32'd8007: dataIn1 = 32'd429
; 
32'd8008: dataIn1 = 32'd368
; 
32'd8009: dataIn1 = 32'd369
; 
32'd8010: dataIn1 = 32'd372
; 
32'd8011: dataIn1 = 32'd370
; 
32'd8012: dataIn1 = 32'd372
; 
32'd8013: dataIn1 = 32'd371
; 
32'd8014: dataIn1 = 32'd372
; 
32'd8015: dataIn1 = 32'd431
; 
32'd8016: dataIn1 = 32'd372
; 
32'd8017: dataIn1 = 32'd398
; 
32'd8018: dataIn1 = 32'd404
; 
32'd8019: dataIn1 = 32'd373
; 
32'd8020: dataIn1 = 32'd375
; 
32'd8021: dataIn1 = 32'd431
; 
32'd8022: dataIn1 = 32'd374
; 
32'd8023: dataIn1 = 32'd378
; 
32'd8024: dataIn1 = 32'd375
; 
32'd8025: dataIn1 = 32'd377
; 
32'd8026: dataIn1 = 32'd398
; 
32'd8027: dataIn1 = 32'd411
; 
32'd8028: dataIn1 = 32'd376
; 
32'd8029: dataIn1 = 32'd378
; 
32'd8030: dataIn1 = 32'd392
; 
32'd8031: dataIn1 = 32'd448
; 
32'd8032: dataIn1 = 32'd377
; 
32'd8033: dataIn1 = 32'd380
; 
32'd8034: dataIn1 = 32'd381
; 
32'd8035: dataIn1 = 32'd384
; 
32'd8036: dataIn1 = 32'd385
; 
32'd8037: dataIn1 = 32'd390
; 
32'd8038: dataIn1 = 32'd447
; 
32'd8039: dataIn1 = 32'd378
; 
32'd8040: dataIn1 = 32'd379
; 
32'd8041: dataIn1 = 32'd388
; 
32'd8042: dataIn1 = 32'd390
; 
32'd8043: dataIn1 = 32'd447
; 
32'd8044: dataIn1 = 32'd379
; 
32'd8045: dataIn1 = 32'd387
; 
32'd8046: dataIn1 = 32'd380
; 
32'd8047: dataIn1 = 32'd381
; 
32'd8048: dataIn1 = 32'd381
; 
32'd8049: dataIn1 = 32'd383
; 
32'd8050: dataIn1 = 32'd382
; 
32'd8051: dataIn1 = 32'd383
; 
32'd8052: dataIn1 = 32'd383
; 
32'd8053: dataIn1 = 32'd384
; 
32'd8054: dataIn1 = 32'd384
; 
32'd8055: dataIn1 = 32'd385
; 
32'd8056: dataIn1 = 32'd390
; 
32'd8057: dataIn1 = 32'd447
; 
32'd8058: dataIn1 = 32'd386
; 
32'd8059: dataIn1 = 32'd388
; 
32'd8060: dataIn1 = 32'd387
; 
32'd8061: dataIn1 = 32'd388
; 
32'd8062: dataIn1 = 32'd393
; 
32'd8063: dataIn1 = 32'd447
; 
32'd8064: dataIn1 = 32'd388
; 
32'd8065: dataIn1 = 32'd389
; 
32'd8066: dataIn1 = 32'd393
; 
32'd8067: dataIn1 = 32'd389
; 
32'd8068: dataIn1 = 32'd390
; 
32'd8069: dataIn1 = 32'd393
; 
32'd8070: dataIn1 = 32'd390
; 
32'd8071: dataIn1 = 32'd391
; 
32'd8072: dataIn1 = 32'd391
; 
32'd8073: dataIn1 = 32'd394
; 
32'd8074: dataIn1 = 32'd392
; 
32'd8075: dataIn1 = 32'd393
; 
32'd8076: dataIn1 = 32'd406
; 
32'd8077: dataIn1 = 32'd393
; 
32'd8078: dataIn1 = 32'd394
; 
32'd8079: dataIn1 = 32'd395
; 
32'd8080: dataIn1 = 32'd398
; 
32'd8081: dataIn1 = 32'd403
; 
32'd8082: dataIn1 = 32'd404
; 
32'd8083: dataIn1 = 32'd411
; 
32'd8084: dataIn1 = 32'd431
; 
32'd8085: dataIn1 = 32'd394
; 
32'd8086: dataIn1 = 32'd395
; 
32'd8087: dataIn1 = 32'd396
; 
32'd8088: dataIn1 = 32'd395
; 
32'd8089: dataIn1 = 32'd398
; 
32'd8090: dataIn1 = 32'd404
; 
32'd8091: dataIn1 = 32'd411
; 
32'd8092: dataIn1 = 32'd396
; 
32'd8093: dataIn1 = 32'd397
; 
32'd8094: dataIn1 = 32'd397
; 
32'd8095: dataIn1 = 32'd410
; 
32'd8096: dataIn1 = 32'd398
; 
32'd8097: dataIn1 = 32'd403
; 
32'd8098: dataIn1 = 32'd404
; 
32'd8099: dataIn1 = 32'd411
; 
32'd8100: dataIn1 = 32'd399
; 
32'd8101: dataIn1 = 32'd401
; 
32'd8102: dataIn1 = 32'd402
; 
32'd8103: dataIn1 = 32'd400
; 
32'd8104: dataIn1 = 32'd401
; 
32'd8105: dataIn1 = 32'd403
; 
32'd8106: dataIn1 = 32'd401
; 
32'd8107: dataIn1 = 32'd408
; 
32'd8108: dataIn1 = 32'd402
; 
32'd8109: dataIn1 = 32'd429
; 
32'd8110: dataIn1 = 32'd403
; 
32'd8111: dataIn1 = 32'd404
; 
32'd8112: dataIn1 = 32'd407
; 
32'd8113: dataIn1 = 32'd411
; 
32'd8114: dataIn1 = 32'd404
; 
32'd8115: dataIn1 = 32'd411
; 
32'd8116: dataIn1 = 32'd429
; 
32'd8117: dataIn1 = 32'd405
; 
32'd8118: dataIn1 = 32'd407
; 
32'd8119: dataIn1 = 32'd408
; 
32'd8120: dataIn1 = 32'd406
; 
32'd8121: dataIn1 = 32'd407
; 
32'd8122: dataIn1 = 32'd421
; 
32'd8123: dataIn1 = 32'd428
; 
32'd8124: dataIn1 = 32'd407
; 
32'd8125: dataIn1 = 32'd410
; 
32'd8126: dataIn1 = 32'd412
; 
32'd8127: dataIn1 = 32'd413
; 
32'd8128: dataIn1 = 32'd408
; 
32'd8129: dataIn1 = 32'd416
; 
32'd8130: dataIn1 = 32'd409
; 
32'd8131: dataIn1 = 32'd410
; 
32'd8132: dataIn1 = 32'd411
; 
32'd8133: dataIn1 = 32'd414
; 
32'd8134: dataIn1 = 32'd417
; 
32'd8135: dataIn1 = 32'd411
; 
32'd8136: dataIn1 = 32'd412
; 
32'd8137: dataIn1 = 32'd413
; 
32'd8138: dataIn1 = 32'd413
; 
32'd8139: dataIn1 = 32'd414
; 
32'd8140: dataIn1 = 32'd417
; 
32'd8141: dataIn1 = 32'd414
; 
32'd8142: dataIn1 = 32'd415
; 
32'd8143: dataIn1 = 32'd417
; 
32'd8144: dataIn1 = 32'd415
; 
32'd8145: dataIn1 = 32'd416
; 
32'd8146: dataIn1 = 32'd417
; 
32'd8147: dataIn1 = 32'd425
; 
32'd8148: dataIn1 = 32'd416
; 
32'd8149: dataIn1 = 32'd417
; 
32'd8150: dataIn1 = 32'd417
; 
32'd8151: dataIn1 = 32'd418
; 
32'd8152: dataIn1 = 32'd419
; 
32'd8153: dataIn1 = 32'd418
; 
32'd8154: dataIn1 = 32'd422
; 
32'd8155: dataIn1 = 32'd419
; 
32'd8156: dataIn1 = 32'd420
; 
32'd8157: dataIn1 = 32'd422
; 
32'd8158: dataIn1 = 32'd420
; 
32'd8159: dataIn1 = 32'd423
; 
32'd8160: dataIn1 = 32'd421
; 
32'd8161: dataIn1 = 32'd422
; 
32'd8162: dataIn1 = 32'd422
; 
32'd8163: dataIn1 = 32'd423
; 
32'd8164: dataIn1 = 32'd424
; 
32'd8165: dataIn1 = 32'd430
; 
32'd8166: dataIn1 = 32'd425
; 
32'd8167: dataIn1 = 32'd426
; 
32'd8168: dataIn1 = 32'd427
; 
32'd8169: dataIn1 = 32'd524
; 
32'd8170: dataIn1 = 32'd427
; 
32'd8171: dataIn1 = 32'd442
; 
32'd8172: dataIn1 = 32'd428
; 
32'd8173: dataIn1 = 32'd429
; 
32'd8174: dataIn1 = 32'd429
; 
32'd8175: dataIn1 = 32'd430
; 
32'd8176: dataIn1 = 32'd431
; 
32'd8177: dataIn1 = 32'd432
; 
32'd8178: dataIn1 = 32'd444
; 
32'd8179: dataIn1 = 32'd446
; 
32'd8180: dataIn1 = 32'd433
; 
32'd8181: dataIn1 = 32'd434
; 
32'd8182: dataIn1 = 32'd435
; 
32'd8183: dataIn1 = 32'd444
; 
32'd8184: dataIn1 = 32'd446
; 
32'd8185: dataIn1 = 32'd436
; 
32'd8186: dataIn1 = 32'd437
; 
32'd8187: dataIn1 = 32'd438
; 
32'd8188: dataIn1 = 32'd438
; 
32'd8189: dataIn1 = 32'd504
; 
32'd8190: dataIn1 = 32'd439
; 
32'd8191: dataIn1 = 32'd440
; 
32'd8192: dataIn1 = 32'd456
; 
32'd8193: dataIn1 = 32'd440
; 
32'd8194: dataIn1 = 32'd456
; 
32'd8195: dataIn1 = 32'd441
; 
32'd8196: dataIn1 = 32'd442
; 
32'd8197: dataIn1 = 32'd443
; 
32'd8198: dataIn1 = 32'd444
; 
32'd8199: dataIn1 = 32'd445
; 
32'd8200: dataIn1 = 32'd446
; 
32'd8201: dataIn1 = 32'd445
; 
32'd8202: dataIn1 = 32'd446
; 
32'd8203: dataIn1 = 32'd447
; 
32'd8204: dataIn1 = 32'd448
; 
32'd8205: dataIn1 = 32'd448
; 
32'd8206: dataIn1 = 32'd449
; 
32'd8207: dataIn1 = 32'd463
; 
32'd8208: dataIn1 = 32'd465
; 
32'd8209: dataIn1 = 32'd502
; 
32'd8210: dataIn1 = 32'd450
; 
32'd8211: dataIn1 = 32'd466
; 
32'd8212: dataIn1 = 32'd467
; 
32'd8213: dataIn1 = 32'd482
; 
32'd8214: dataIn1 = 32'd451
; 
32'd8215: dataIn1 = 32'd457
; 
32'd8216: dataIn1 = 32'd460
; 
32'd8217: dataIn1 = 32'd668
; 
32'd8218: dataIn1 = 32'd452
; 
32'd8219: dataIn1 = 32'd453
; 
32'd8220: dataIn1 = 32'd454
; 
32'd8221: dataIn1 = 32'd455
; 
32'd8222: dataIn1 = 32'd534
; 
32'd8223: dataIn1 = 32'd453
; 
32'd8224: dataIn1 = 32'd454
; 
32'd8225: dataIn1 = 32'd486
; 
32'd8226: dataIn1 = 32'd512
; 
32'd8227: dataIn1 = 32'd533
; 
32'd8228: dataIn1 = 32'd454
; 
32'd8229: dataIn1 = 32'd471
; 
32'd8230: dataIn1 = 32'd475
; 
32'd8231: dataIn1 = 32'd455
; 
32'd8232: dataIn1 = 32'd462
; 
32'd8233: dataIn1 = 32'd535
; 
32'd8234: dataIn1 = 32'd456
; 
32'd8235: dataIn1 = 32'd466
; 
32'd8236: dataIn1 = 32'd484
; 
32'd8237: dataIn1 = 32'd504
; 
32'd8238: dataIn1 = 32'd457
; 
32'd8239: dataIn1 = 32'd461
; 
32'd8240: dataIn1 = 32'd458
; 
32'd8241: dataIn1 = 32'd466
; 
32'd8242: dataIn1 = 32'd467
; 
32'd8243: dataIn1 = 32'd542
; 
32'd8244: dataIn1 = 32'd459
; 
32'd8245: dataIn1 = 32'd460
; 
32'd8246: dataIn1 = 32'd479
; 
32'd8247: dataIn1 = 32'd668
; 
32'd8248: dataIn1 = 32'd460
; 
32'd8249: dataIn1 = 32'd461
; 
32'd8250: dataIn1 = 32'd462
; 
32'd8251: dataIn1 = 32'd518
; 
32'd8252: dataIn1 = 32'd461
; 
32'd8253: dataIn1 = 32'd465
; 
32'd8254: dataIn1 = 32'd477
; 
32'd8255: dataIn1 = 32'd542
; 
32'd8256: dataIn1 = 32'd462
; 
32'd8257: dataIn1 = 32'd463
; 
32'd8258: dataIn1 = 32'd465
; 
32'd8259: dataIn1 = 32'd463
; 
32'd8260: dataIn1 = 32'd557
; 
32'd8261: dataIn1 = 32'd464
; 
32'd8262: dataIn1 = 32'd473
; 
32'd8263: dataIn1 = 32'd479
; 
32'd8264: dataIn1 = 32'd665
; 
32'd8265: dataIn1 = 32'd465
; 
32'd8266: dataIn1 = 32'd477
; 
32'd8267: dataIn1 = 32'd518
; 
32'd8268: dataIn1 = 32'd466
; 
32'd8269: dataIn1 = 32'd467
; 
32'd8270: dataIn1 = 32'd472
; 
32'd8271: dataIn1 = 32'd477
; 
32'd8272: dataIn1 = 32'd484
; 
32'd8273: dataIn1 = 32'd543
; 
32'd8274: dataIn1 = 32'd468
; 
32'd8275: dataIn1 = 32'd476
; 
32'd8276: dataIn1 = 32'd481
; 
32'd8277: dataIn1 = 32'd501
; 
32'd8278: dataIn1 = 32'd469
; 
32'd8279: dataIn1 = 32'd474
; 
32'd8280: dataIn1 = 32'd665
; 
32'd8281: dataIn1 = 32'd667
; 
32'd8282: dataIn1 = 32'd470
; 
32'd8283: dataIn1 = 32'd478
; 
32'd8284: dataIn1 = 32'd485
; 
32'd8285: dataIn1 = 32'd546
; 
32'd8286: dataIn1 = 32'd597
; 
32'd8287: dataIn1 = 32'd598
; 
32'd8288: dataIn1 = 32'd471
; 
32'd8289: dataIn1 = 32'd475
; 
32'd8290: dataIn1 = 32'd547
; 
32'd8291: dataIn1 = 32'd472
; 
32'd8292: dataIn1 = 32'd477
; 
32'd8293: dataIn1 = 32'd482
; 
32'd8294: dataIn1 = 32'd489
; 
32'd8295: dataIn1 = 32'd523
; 
32'd8296: dataIn1 = 32'd473
; 
32'd8297: dataIn1 = 32'd478
; 
32'd8298: dataIn1 = 32'd483
; 
32'd8299: dataIn1 = 32'd666
; 
32'd8300: dataIn1 = 32'd474
; 
32'd8301: dataIn1 = 32'd479
; 
32'd8302: dataIn1 = 32'd525
; 
32'd8303: dataIn1 = 32'd666
; 
32'd8304: dataIn1 = 32'd475
; 
32'd8305: dataIn1 = 32'd597
; 
32'd8306: dataIn1 = 32'd476
; 
32'd8307: dataIn1 = 32'd481
; 
32'd8308: dataIn1 = 32'd488
; 
32'd8309: dataIn1 = 32'd477
; 
32'd8310: dataIn1 = 32'd531
; 
32'd8311: dataIn1 = 32'd478
; 
32'd8312: dataIn1 = 32'd577
; 
32'd8313: dataIn1 = 32'd597
; 
32'd8314: dataIn1 = 32'd479
; 
32'd8315: dataIn1 = 32'd480
; 
32'd8316: dataIn1 = 32'd480
; 
32'd8317: dataIn1 = 32'd525
; 
32'd8318: dataIn1 = 32'd667
; 
32'd8319: dataIn1 = 32'd481
; 
32'd8320: dataIn1 = 32'd489
; 
32'd8321: dataIn1 = 32'd523
; 
32'd8322: dataIn1 = 32'd526
; 
32'd8323: dataIn1 = 32'd482
; 
32'd8324: dataIn1 = 32'd489
; 
32'd8325: dataIn1 = 32'd519
; 
32'd8326: dataIn1 = 32'd523
; 
32'd8327: dataIn1 = 32'd483
; 
32'd8328: dataIn1 = 32'd485
; 
32'd8329: dataIn1 = 32'd484
; 
32'd8330: dataIn1 = 32'd519
; 
32'd8331: dataIn1 = 32'd485
; 
32'd8332: dataIn1 = 32'd545
; 
32'd8333: dataIn1 = 32'd546
; 
32'd8334: dataIn1 = 32'd486
; 
32'd8335: dataIn1 = 32'd487
; 
32'd8336: dataIn1 = 32'd495
; 
32'd8337: dataIn1 = 32'd497
; 
32'd8338: dataIn1 = 32'd499
; 
32'd8339: dataIn1 = 32'd500
; 
32'd8340: dataIn1 = 32'd501
; 
32'd8341: dataIn1 = 32'd512
; 
32'd8342: dataIn1 = 32'd487
; 
32'd8343: dataIn1 = 32'd502
; 
32'd8344: dataIn1 = 32'd521
; 
32'd8345: dataIn1 = 32'd538
; 
32'd8346: dataIn1 = 32'd488
; 
32'd8347: dataIn1 = 32'd489
; 
32'd8348: dataIn1 = 32'd499
; 
32'd8349: dataIn1 = 32'd489
; 
32'd8350: dataIn1 = 32'd491
; 
32'd8351: dataIn1 = 32'd492
; 
32'd8352: dataIn1 = 32'd503
; 
32'd8353: dataIn1 = 32'd508
; 
32'd8354: dataIn1 = 32'd519
; 
32'd8355: dataIn1 = 32'd523
; 
32'd8356: dataIn1 = 32'd536
; 
32'd8357: dataIn1 = 32'd490
; 
32'd8358: dataIn1 = 32'd514
; 
32'd8359: dataIn1 = 32'd521
; 
32'd8360: dataIn1 = 32'd527
; 
32'd8361: dataIn1 = 32'd529
; 
32'd8362: dataIn1 = 32'd491
; 
32'd8363: dataIn1 = 32'd502
; 
32'd8364: dataIn1 = 32'd522
; 
32'd8365: dataIn1 = 32'd492
; 
32'd8366: dataIn1 = 32'd498
; 
32'd8367: dataIn1 = 32'd503
; 
32'd8368: dataIn1 = 32'd508
; 
32'd8369: dataIn1 = 32'd520
; 
32'd8370: dataIn1 = 32'd536
; 
32'd8371: dataIn1 = 32'd540
; 
32'd8372: dataIn1 = 32'd493
; 
32'd8373: dataIn1 = 32'd506
; 
32'd8374: dataIn1 = 32'd509
; 
32'd8375: dataIn1 = 32'd515
; 
32'd8376: dataIn1 = 32'd494
; 
32'd8377: dataIn1 = 32'd511
; 
32'd8378: dataIn1 = 32'd495
; 
32'd8379: dataIn1 = 32'd517
; 
32'd8380: dataIn1 = 32'd544
; 
32'd8381: dataIn1 = 32'd496
; 
32'd8382: dataIn1 = 32'd497
; 
32'd8383: dataIn1 = 32'd509
; 
32'd8384: dataIn1 = 32'd520
; 
32'd8385: dataIn1 = 32'd497
; 
32'd8386: dataIn1 = 32'd498
; 
32'd8387: dataIn1 = 32'd500
; 
32'd8388: dataIn1 = 32'd521
; 
32'd8389: dataIn1 = 32'd498
; 
32'd8390: dataIn1 = 32'd520
; 
32'd8391: dataIn1 = 32'd540
; 
32'd8392: dataIn1 = 32'd499
; 
32'd8393: dataIn1 = 32'd500
; 
32'd8394: dataIn1 = 32'd500
; 
32'd8395: dataIn1 = 32'd501
; 
32'd8396: dataIn1 = 32'd502
; 
32'd8397: dataIn1 = 32'd502
; 
32'd8398: dataIn1 = 32'd526
; 
32'd8399: dataIn1 = 32'd503
; 
32'd8400: dataIn1 = 32'd540
; 
32'd8401: dataIn1 = 32'd504
; 
32'd8402: dataIn1 = 32'd505
; 
32'd8403: dataIn1 = 32'd505
; 
32'd8404: dataIn1 = 32'd508
; 
32'd8405: dataIn1 = 32'd506
; 
32'd8406: dataIn1 = 32'd508
; 
32'd8407: dataIn1 = 32'd507
; 
32'd8408: dataIn1 = 32'd508
; 
32'd8409: dataIn1 = 32'd508
; 
32'd8410: dataIn1 = 32'd536
; 
32'd8411: dataIn1 = 32'd509
; 
32'd8412: dataIn1 = 32'd529
; 
32'd8413: dataIn1 = 32'd510
; 
32'd8414: dataIn1 = 32'd515
; 
32'd8415: dataIn1 = 32'd517
; 
32'd8416: dataIn1 = 32'd511
; 
32'd8417: dataIn1 = 32'd512
; 
32'd8418: dataIn1 = 32'd517
; 
32'd8419: dataIn1 = 32'd528
; 
32'd8420: dataIn1 = 32'd512
; 
32'd8421: dataIn1 = 32'd513
; 
32'd8422: dataIn1 = 32'd515
; 
32'd8423: dataIn1 = 32'd544
; 
32'd8424: dataIn1 = 32'd514
; 
32'd8425: dataIn1 = 32'd516
; 
32'd8426: dataIn1 = 32'd532
; 
32'd8427: dataIn1 = 32'd538
; 
32'd8428: dataIn1 = 32'd515
; 
32'd8429: dataIn1 = 32'd516
; 
32'd8430: dataIn1 = 32'd516
; 
32'd8431: dataIn1 = 32'd517
; 
32'd8432: dataIn1 = 32'd544
; 
32'd8433: dataIn1 = 32'd518
; 
32'd8434: dataIn1 = 32'd531
; 
32'd8435: dataIn1 = 32'd519
; 
32'd8436: dataIn1 = 32'd520
; 
32'd8437: dataIn1 = 32'd527
; 
32'd8438: dataIn1 = 32'd521
; 
32'd8439: dataIn1 = 32'd522
; 
32'd8440: dataIn1 = 32'd523
; 
32'd8441: dataIn1 = 32'd526
; 
32'd8442: dataIn1 = 32'd531
; 
32'd8443: dataIn1 = 32'd523
; 
32'd8444: dataIn1 = 32'd524
; 
32'd8445: dataIn1 = 32'd537
; 
32'd8446: dataIn1 = 32'd543
; 
32'd8447: dataIn1 = 32'd525
; 
32'd8448: dataIn1 = 32'd558
; 
32'd8449: dataIn1 = 32'd526
; 
32'd8450: dataIn1 = 32'd527
; 
32'd8451: dataIn1 = 32'd529
; 
32'd8452: dataIn1 = 32'd530
; 
32'd8453: dataIn1 = 32'd528
; 
32'd8454: dataIn1 = 32'd529
; 
32'd8455: dataIn1 = 32'd530
; 
32'd8456: dataIn1 = 32'd536
; 
32'd8457: dataIn1 = 32'd531
; 
32'd8458: dataIn1 = 32'd543
; 
32'd8459: dataIn1 = 32'd532
; 
32'd8460: dataIn1 = 32'd533
; 
32'd8461: dataIn1 = 32'd533
; 
32'd8462: dataIn1 = 32'd534
; 
32'd8463: dataIn1 = 32'd534
; 
32'd8464: dataIn1 = 32'd535
; 
32'd8465: dataIn1 = 32'd535
; 
32'd8466: dataIn1 = 32'd557
; 
32'd8467: dataIn1 = 32'd536
; 
32'd8468: dataIn1 = 32'd537
; 
32'd8469: dataIn1 = 32'd537
; 
32'd8470: dataIn1 = 32'd538
; 
32'd8471: dataIn1 = 32'd544
; 
32'd8472: dataIn1 = 32'd539
; 
32'd8473: dataIn1 = 32'd577
; 
32'd8474: dataIn1 = 32'd598
; 
32'd8475: dataIn1 = 32'd540
; 
32'd8476: dataIn1 = 32'd541
; 
32'd8477: dataIn1 = 32'd542
; 
32'd8478: dataIn1 = 32'd542
; 
32'd8479: dataIn1 = 32'd543
; 
32'd8480: dataIn1 = 32'd544
; 
32'd8481: dataIn1 = 32'd545
; 
32'd8482: dataIn1 = 32'd546
; 
32'd8483: dataIn1 = 32'd547
; 
32'd8484: dataIn1 = 32'd548
; 
32'd8485: dataIn1 = 32'd549
; 
32'd8486: dataIn1 = 32'd546
; 
32'd8487: dataIn1 = 32'd547
; 
32'd8488: dataIn1 = 32'd548
; 
32'd8489: dataIn1 = 32'd597
; 
32'd8490: dataIn1 = 32'd549
; 
32'd8491: dataIn1 = 32'd597
; 
32'd8492: dataIn1 = 32'd550
; 
32'd8493: dataIn1 = 32'd551
; 
32'd8494: dataIn1 = 32'd555
; 
32'd8495: dataIn1 = 32'd563
; 
32'd8496: dataIn1 = 32'd612
; 
32'd8497: dataIn1 = 32'd636
; 
32'd8498: dataIn1 = 32'd643
; 
32'd8499: dataIn1 = 32'd654
; 
32'd8500: dataIn1 = 32'd551
; 
32'd8501: dataIn1 = 32'd653
; 
32'd8502: dataIn1 = 32'd552
; 
32'd8503: dataIn1 = 32'd553
; 
32'd8504: dataIn1 = 32'd554
; 
32'd8505: dataIn1 = 32'd579
; 
32'd8506: dataIn1 = 32'd630
; 
32'd8507: dataIn1 = 32'd641
; 
32'd8508: dataIn1 = 32'd553
; 
32'd8509: dataIn1 = 32'd583
; 
32'd8510: dataIn1 = 32'd584
; 
32'd8511: dataIn1 = 32'd591
; 
32'd8512: dataIn1 = 32'd605
; 
32'd8513: dataIn1 = 32'd649
; 
32'd8514: dataIn1 = 32'd650
; 
32'd8515: dataIn1 = 32'd554
; 
32'd8516: dataIn1 = 32'd578
; 
32'd8517: dataIn1 = 32'd591
; 
32'd8518: dataIn1 = 32'd607
; 
32'd8519: dataIn1 = 32'd612
; 
32'd8520: dataIn1 = 32'd617
; 
32'd8521: dataIn1 = 32'd623
; 
32'd8522: dataIn1 = 32'd634
; 
32'd8523: dataIn1 = 32'd658
; 
32'd8524: dataIn1 = 32'd555
; 
32'd8525: dataIn1 = 32'd614
; 
32'd8526: dataIn1 = 32'd627
; 
32'd8527: dataIn1 = 32'd556
; 
32'd8528: dataIn1 = 32'd558
; 
32'd8529: dataIn1 = 32'd612
; 
32'd8530: dataIn1 = 32'd627
; 
32'd8531: dataIn1 = 32'd632
; 
32'd8532: dataIn1 = 32'd635
; 
32'd8533: dataIn1 = 32'd557
; 
32'd8534: dataIn1 = 32'd558
; 
32'd8535: dataIn1 = 32'd639
; 
32'd8536: dataIn1 = 32'd558
; 
32'd8537: dataIn1 = 32'd559
; 
32'd8538: dataIn1 = 32'd561
; 
32'd8539: dataIn1 = 32'd577
; 
32'd8540: dataIn1 = 32'd601
; 
32'd8541: dataIn1 = 32'd617
; 
32'd8542: dataIn1 = 32'd560
; 
32'd8543: dataIn1 = 32'd562
; 
32'd8544: dataIn1 = 32'd577
; 
32'd8545: dataIn1 = 32'd578
; 
32'd8546: dataIn1 = 32'd600
; 
32'd8547: dataIn1 = 32'd561
; 
32'd8548: dataIn1 = 32'd566
; 
32'd8549: dataIn1 = 32'd567
; 
32'd8550: dataIn1 = 32'd579
; 
32'd8551: dataIn1 = 32'd562
; 
32'd8552: dataIn1 = 32'd563
; 
32'd8553: dataIn1 = 32'd565
; 
32'd8554: dataIn1 = 32'd577
; 
32'd8555: dataIn1 = 32'd603
; 
32'd8556: dataIn1 = 32'd563
; 
32'd8557: dataIn1 = 32'd564
; 
32'd8558: dataIn1 = 32'd648
; 
32'd8559: dataIn1 = 32'd564
; 
32'd8560: dataIn1 = 32'd565
; 
32'd8561: dataIn1 = 32'd570
; 
32'd8562: dataIn1 = 32'd613
; 
32'd8563: dataIn1 = 32'd614
; 
32'd8564: dataIn1 = 32'd565
; 
32'd8565: dataIn1 = 32'd570
; 
32'd8566: dataIn1 = 32'd624
; 
32'd8567: dataIn1 = 32'd643
; 
32'd8568: dataIn1 = 32'd566
; 
32'd8569: dataIn1 = 32'd568
; 
32'd8570: dataIn1 = 32'd569
; 
32'd8571: dataIn1 = 32'd625
; 
32'd8572: dataIn1 = 32'd642
; 
32'd8573: dataIn1 = 32'd567
; 
32'd8574: dataIn1 = 32'd569
; 
32'd8575: dataIn1 = 32'd576
; 
32'd8576: dataIn1 = 32'd645
; 
32'd8577: dataIn1 = 32'd568
; 
32'd8578: dataIn1 = 32'd570
; 
32'd8579: dataIn1 = 32'd569
; 
32'd8580: dataIn1 = 32'd570
; 
32'd8581: dataIn1 = 32'd613
; 
32'd8582: dataIn1 = 32'd614
; 
32'd8583: dataIn1 = 32'd570
; 
32'd8584: dataIn1 = 32'd571
; 
32'd8585: dataIn1 = 32'd640
; 
32'd8586: dataIn1 = 32'd663
; 
32'd8587: dataIn1 = 32'd571
; 
32'd8588: dataIn1 = 32'd593
; 
32'd8589: dataIn1 = 32'd652
; 
32'd8590: dataIn1 = 32'd572
; 
32'd8591: dataIn1 = 32'd573
; 
32'd8592: dataIn1 = 32'd593
; 
32'd8593: dataIn1 = 32'd660
; 
32'd8594: dataIn1 = 32'd573
; 
32'd8595: dataIn1 = 32'd616
; 
32'd8596: dataIn1 = 32'd647
; 
32'd8597: dataIn1 = 32'd648
; 
32'd8598: dataIn1 = 32'd574
; 
32'd8599: dataIn1 = 32'd601
; 
32'd8600: dataIn1 = 32'd618
; 
32'd8601: dataIn1 = 32'd637
; 
32'd8602: dataIn1 = 32'd575
; 
32'd8603: dataIn1 = 32'd577
; 
32'd8604: dataIn1 = 32'd600
; 
32'd8605: dataIn1 = 32'd601
; 
32'd8606: dataIn1 = 32'd576
; 
32'd8607: dataIn1 = 32'd618
; 
32'd8608: dataIn1 = 32'd659
; 
32'd8609: dataIn1 = 32'd577
; 
32'd8610: dataIn1 = 32'd578
; 
32'd8611: dataIn1 = 32'd590
; 
32'd8612: dataIn1 = 32'd595
; 
32'd8613: dataIn1 = 32'd579
; 
32'd8614: dataIn1 = 32'd605
; 
32'd8615: dataIn1 = 32'd625
; 
32'd8616: dataIn1 = 32'd580
; 
32'd8617: dataIn1 = 32'd581
; 
32'd8618: dataIn1 = 32'd583
; 
32'd8619: dataIn1 = 32'd581
; 
32'd8620: dataIn1 = 32'd582
; 
32'd8621: dataIn1 = 32'd586
; 
32'd8622: dataIn1 = 32'd611
; 
32'd8623: dataIn1 = 32'd619
; 
32'd8624: dataIn1 = 32'd582
; 
32'd8625: dataIn1 = 32'd583
; 
32'd8626: dataIn1 = 32'd649
; 
32'd8627: dataIn1 = 32'd583
; 
32'd8628: dataIn1 = 32'd603
; 
32'd8629: dataIn1 = 32'd606
; 
32'd8630: dataIn1 = 32'd584
; 
32'd8631: dataIn1 = 32'd606
; 
32'd8632: dataIn1 = 32'd622
; 
32'd8633: dataIn1 = 32'd585
; 
32'd8634: dataIn1 = 32'd619
; 
32'd8635: dataIn1 = 32'd622
; 
32'd8636: dataIn1 = 32'd646
; 
32'd8637: dataIn1 = 32'd586
; 
32'd8638: dataIn1 = 32'd587
; 
32'd8639: dataIn1 = 32'd661
; 
32'd8640: dataIn1 = 32'd587
; 
32'd8641: dataIn1 = 32'd589
; 
32'd8642: dataIn1 = 32'd606
; 
32'd8643: dataIn1 = 32'd588
; 
32'd8644: dataIn1 = 32'd589
; 
32'd8645: dataIn1 = 32'd644
; 
32'd8646: dataIn1 = 32'd646
; 
32'd8647: dataIn1 = 32'd589
; 
32'd8648: dataIn1 = 32'd590
; 
32'd8649: dataIn1 = 32'd592
; 
32'd8650: dataIn1 = 32'd609
; 
32'd8651: dataIn1 = 32'd590
; 
32'd8652: dataIn1 = 32'd617
; 
32'd8653: dataIn1 = 32'd623
; 
32'd8654: dataIn1 = 32'd658
; 
32'd8655: dataIn1 = 32'd591
; 
32'd8656: dataIn1 = 32'd603
; 
32'd8657: dataIn1 = 32'd629
; 
32'd8658: dataIn1 = 32'd653
; 
32'd8659: dataIn1 = 32'd592
; 
32'd8660: dataIn1 = 32'd594
; 
32'd8661: dataIn1 = 32'd595
; 
32'd8662: dataIn1 = 32'd608
; 
32'd8663: dataIn1 = 32'd593
; 
32'd8664: dataIn1 = 32'd652
; 
32'd8665: dataIn1 = 32'd594
; 
32'd8666: dataIn1 = 32'd595
; 
32'd8667: dataIn1 = 32'd596
; 
32'd8668: dataIn1 = 32'd602
; 
32'd8669: dataIn1 = 32'd595
; 
32'd8670: dataIn1 = 32'd596
; 
32'd8671: dataIn1 = 32'd597
; 
32'd8672: dataIn1 = 32'd602
; 
32'd8673: dataIn1 = 32'd607
; 
32'd8674: dataIn1 = 32'd597
; 
32'd8675: dataIn1 = 32'd602
; 
32'd8676: dataIn1 = 32'd598
; 
32'd8677: dataIn1 = 32'd599
; 
32'd8678: dataIn1 = 32'd604
; 
32'd8679: dataIn1 = 32'd611
; 
32'd8680: dataIn1 = 32'd619
; 
32'd8681: dataIn1 = 32'd646
; 
32'd8682: dataIn1 = 32'd651
; 
32'd8683: dataIn1 = 32'd600
; 
32'd8684: dataIn1 = 32'd647
; 
32'd8685: dataIn1 = 32'd601
; 
32'd8686: dataIn1 = 32'd602
; 
32'd8687: dataIn1 = 32'd603
; 
32'd8688: dataIn1 = 32'd624
; 
32'd8689: dataIn1 = 32'd604
; 
32'd8690: dataIn1 = 32'd605
; 
32'd8691: dataIn1 = 32'd650
; 
32'd8692: dataIn1 = 32'd605
; 
32'd8693: dataIn1 = 32'd644
; 
32'd8694: dataIn1 = 32'd651
; 
32'd8695: dataIn1 = 32'd606
; 
32'd8696: dataIn1 = 32'd607
; 
32'd8697: dataIn1 = 32'd608
; 
32'd8698: dataIn1 = 32'd621
; 
32'd8699: dataIn1 = 32'd655
; 
32'd8700: dataIn1 = 32'd608
; 
32'd8701: dataIn1 = 32'd609
; 
32'd8702: dataIn1 = 32'd609
; 
32'd8703: dataIn1 = 32'd610
; 
32'd8704: dataIn1 = 32'd623
; 
32'd8705: dataIn1 = 32'd658
; 
32'd8706: dataIn1 = 32'd610
; 
32'd8707: dataIn1 = 32'd622
; 
32'd8708: dataIn1 = 32'd662
; 
32'd8709: dataIn1 = 32'd611
; 
32'd8710: dataIn1 = 32'd649
; 
32'd8711: dataIn1 = 32'd661
; 
32'd8712: dataIn1 = 32'd612
; 
32'd8713: dataIn1 = 32'd645
; 
32'd8714: dataIn1 = 32'd664
; 
32'd8715: dataIn1 = 32'd613
; 
32'd8716: dataIn1 = 32'd614
; 
32'd8717: dataIn1 = 32'd645
; 
32'd8718: dataIn1 = 32'd614
; 
32'd8719: dataIn1 = 32'd615
; 
32'd8720: dataIn1 = 32'd616
; 
32'd8721: dataIn1 = 32'd636
; 
32'd8722: dataIn1 = 32'd648
; 
32'd8723: dataIn1 = 32'd616
; 
32'd8724: dataIn1 = 32'd618
; 
32'd8725: dataIn1 = 32'd620
; 
32'd8726: dataIn1 = 32'd637
; 
32'd8727: dataIn1 = 32'd659
; 
32'd8728: dataIn1 = 32'd617
; 
32'd8729: dataIn1 = 32'd618
; 
32'd8730: dataIn1 = 32'd652
; 
32'd8731: dataIn1 = 32'd619
; 
32'd8732: dataIn1 = 32'd650
; 
32'd8733: dataIn1 = 32'd620
; 
32'd8734: dataIn1 = 32'd652
; 
32'd8735: dataIn1 = 32'd621
; 
32'd8736: dataIn1 = 32'd655
; 
32'd8737: dataIn1 = 32'd622
; 
32'd8738: dataIn1 = 32'd661
; 
32'd8739: dataIn1 = 32'd623
; 
32'd8740: dataIn1 = 32'd624
; 
32'd8741: dataIn1 = 32'd625
; 
32'd8742: dataIn1 = 32'd629
; 
32'd8743: dataIn1 = 32'd625
; 
32'd8744: dataIn1 = 32'd630
; 
32'd8745: dataIn1 = 32'd626
; 
32'd8746: dataIn1 = 32'd627
; 
32'd8747: dataIn1 = 32'd633
; 
32'd8748: dataIn1 = 32'd627
; 
32'd8749: dataIn1 = 32'd636
; 
32'd8750: dataIn1 = 32'd628
; 
32'd8751: dataIn1 = 32'd637
; 
32'd8752: dataIn1 = 32'd654
; 
32'd8753: dataIn1 = 32'd629
; 
32'd8754: dataIn1 = 32'd630
; 
32'd8755: dataIn1 = 32'd630
; 
32'd8756: dataIn1 = 32'd631
; 
32'd8757: dataIn1 = 32'd645
; 
32'd8758: dataIn1 = 32'd632
; 
32'd8759: dataIn1 = 32'd638
; 
32'd8760: dataIn1 = 32'd639
; 
32'd8761: dataIn1 = 32'd666
; 
32'd8762: dataIn1 = 32'd633
; 
32'd8763: dataIn1 = 32'd634
; 
32'd8764: dataIn1 = 32'd656
; 
32'd8765: dataIn1 = 32'd634
; 
32'd8766: dataIn1 = 32'd635
; 
32'd8767: dataIn1 = 32'd636
; 
32'd8768: dataIn1 = 32'd637
; 
32'd8769: dataIn1 = 32'd647
; 
32'd8770: dataIn1 = 32'd638
; 
32'd8771: dataIn1 = 32'd657
; 
32'd8772: dataIn1 = 32'd664
; 
32'd8773: dataIn1 = 32'd639
; 
32'd8774: dataIn1 = 32'd640
; 
32'd8775: dataIn1 = 32'd645
; 
32'd8776: dataIn1 = 32'd641
; 
32'd8777: dataIn1 = 32'd642
; 
32'd8778: dataIn1 = 32'd645
; 
32'd8779: dataIn1 = 32'd642
; 
32'd8780: dataIn1 = 32'd643
; 
32'd8781: dataIn1 = 32'd644
; 
32'd8782: dataIn1 = 32'd662
; 
32'd8783: dataIn1 = 32'd645
; 
32'd8784: dataIn1 = 32'd659
; 
32'd8785: dataIn1 = 32'd664
; 
32'd8786: dataIn1 = 32'd646
; 
32'd8787: dataIn1 = 32'd647
; 
32'd8788: dataIn1 = 32'd648
; 
32'd8789: dataIn1 = 32'd649
; 
32'd8790: dataIn1 = 32'd650
; 
32'd8791: dataIn1 = 32'd651
; 
32'd8792: dataIn1 = 32'd652
; 
32'd8793: dataIn1 = 32'd653
; 
32'd8794: dataIn1 = 32'd663
; 
32'd8795: dataIn1 = 32'd664
; 
32'd8796: dataIn1 = 32'd654
; 
32'd8797: dataIn1 = 32'd655
; 
32'd8798: dataIn1 = 32'd656
; 
32'd8799: dataIn1 = 32'd657
; 
32'd8800: dataIn1 = 32'd657
; 
32'd8801: dataIn1 = 32'd658
; 
32'd8802: dataIn1 = 32'd659
; 
32'd8803: dataIn1 = 32'd660
; 
32'd8804: dataIn1 = 32'd661
; 
32'd8805: dataIn1 = 32'd662
; 
32'd8806: dataIn1 = 32'd663
; 
32'd8807: dataIn1 = 32'd664
; 
32'd8808: dataIn1 = 32'd665
; 
32'd8809: dataIn1 = 32'd666
; 
32'd8810: dataIn1 = 32'd667
; 
32'd8811: dataIn1 = 32'd668
; 
32'd8812: dataIn1 = 32'd669
; 
32'd8813: dataIn1 = 32'd670
; 
32'd8814: dataIn1 = 32'd670
; 
32'd8815: dataIn1 = 32'd671
; 
32'd8816: dataIn1 = 32'd672
; 
32'd8817: dataIn1 = 32'd672
; 
32'd8818: dataIn1 = 32'd673
; 
32'd8819: dataIn1 = 32'd674
; 
32'd8820: dataIn1 = 32'd675
; 
32'd8821: dataIn1 = 32'd675
; 
32'd8822: dataIn1 = 32'd676
; 
32'd8823: dataIn1 = 32'd678
; 
32'd8824: dataIn1 = 32'd677
; 
32'd8825: dataIn1 = 32'd678
; 
32'd8826: dataIn1 = 32'd679
; 
32'd8827: dataIn1 = 32'd679
; 
32'd8828: dataIn1 = 32'd680
; 
32'd8829: dataIn1 = 32'd680
; 
32'd8830: dataIn1 = 32'd681
; 
32'd8831: dataIn1 = 32'd682
; 
32'd8832: dataIn1 = 32'd682
; 
32'd8833: dataIn1 = 32'd683
; 
32'd8834: dataIn1 = 32'd683
; 
32'd8835: dataIn1 = 32'd684
; 
32'd8836: dataIn1 = 32'd685
; 
default:  
	dataIn1 = 32'd99999; 
endcase 
case(addr2) 
32'd2: dataIn2 = 32'd0; 
32'd3: dataIn2 = 32'd1; 
32'd4: dataIn2 = 32'd1; 
32'd5: dataIn2 = 32'd0; 
32'd6: dataIn2 = 32'd1; 
32'd7: dataIn2 = 32'd0; 
32'd8: dataIn2 = 32'd1; 
32'd9: dataIn2 = 32'd1; 
32'd10: dataIn2 = 32'd1; 
32'd11: dataIn2 = 32'd0; 
32'd12: dataIn2 = 32'd0; 
32'd13: dataIn2 = 32'd1; 
32'd14: dataIn2 = 32'd0; 
32'd15: dataIn2 = 32'd0; 
32'd16: dataIn2 = 32'd1; 
32'd17: dataIn2 = 32'd0; 
32'd18: dataIn2 = 32'd0; 
32'd19: dataIn2 = 32'd1; 
32'd20: dataIn2 = 32'd0; 
32'd21: dataIn2 = 32'd1; 
32'd22: dataIn2 = 32'd0; 
32'd23: dataIn2 = 32'd0; 
32'd24: dataIn2 = 32'd0; 
32'd25: dataIn2 = 32'd0; 
32'd26: dataIn2 = 32'd1; 
32'd27: dataIn2 = 32'd1; 
32'd28: dataIn2 = 32'd0; 
32'd29: dataIn2 = 32'd0; 
32'd30: dataIn2 = 32'd0; 
32'd31: dataIn2 = 32'd1; 
32'd32: dataIn2 = 32'd1; 
32'd33: dataIn2 = 32'd1; 
32'd34: dataIn2 = 32'd0; 
32'd35: dataIn2 = 32'd0; 
32'd36: dataIn2 = 32'd1; 
32'd37: dataIn2 = 32'd1; 
32'd38: dataIn2 = 32'd0; 
32'd39: dataIn2 = 32'd0; 
32'd40: dataIn2 = 32'd1; 
32'd41: dataIn2 = 32'd0; 
32'd42: dataIn2 = 32'd1; 
32'd43: dataIn2 = 32'd0; 
32'd44: dataIn2 = 32'd1; 
32'd45: dataIn2 = 32'd0; 
32'd46: dataIn2 = 32'd0; 
32'd47: dataIn2 = 32'd1; 
32'd48: dataIn2 = 32'd0; 
32'd49: dataIn2 = 32'd0; 
32'd50: dataIn2 = 32'd1; 
32'd51: dataIn2 = 32'd1; 
32'd52: dataIn2 = 32'd0; 
32'd53: dataIn2 = 32'd0; 
32'd54: dataIn2 = 32'd0; 
32'd55: dataIn2 = 32'd0; 
32'd56: dataIn2 = 32'd0; 
32'd57: dataIn2 = 32'd1; 
32'd58: dataIn2 = 32'd0; 
32'd59: dataIn2 = 32'd1; 
32'd60: dataIn2 = 32'd1; 
32'd61: dataIn2 = 32'd0; 
32'd62: dataIn2 = 32'd0; 
32'd63: dataIn2 = 32'd0; 
32'd64: dataIn2 = 32'd1; 
32'd65: dataIn2 = 32'd0; 
32'd66: dataIn2 = 32'd1; 
32'd67: dataIn2 = 32'd1; 
32'd68: dataIn2 = 32'd0; 
32'd69: dataIn2 = 32'd1; 
32'd70: dataIn2 = 32'd0; 
32'd71: dataIn2 = 32'd1; 
32'd72: dataIn2 = 32'd1; 
32'd73: dataIn2 = 32'd0; 
32'd74: dataIn2 = 32'd1; 
32'd75: dataIn2 = 32'd0; 
32'd76: dataIn2 = 32'd1; 
32'd77: dataIn2 = 32'd0; 
32'd78: dataIn2 = 32'd0; 
32'd79: dataIn2 = 32'd0; 
32'd80: dataIn2 = 32'd1; 
32'd81: dataIn2 = 32'd0; 
32'd82: dataIn2 = 32'd0; 
32'd83: dataIn2 = 32'd1; 
32'd84: dataIn2 = 32'd1; 
32'd85: dataIn2 = 32'd1; 
32'd86: dataIn2 = 32'd0; 
32'd87: dataIn2 = 32'd1; 
32'd88: dataIn2 = 32'd0; 
32'd89: dataIn2 = 32'd0; 
32'd90: dataIn2 = 32'd0; 
32'd91: dataIn2 = 32'd1; 
32'd92: dataIn2 = 32'd1; 
32'd93: dataIn2 = 32'd1; 
32'd94: dataIn2 = 32'd0; 
32'd95: dataIn2 = 32'd1; 
32'd96: dataIn2 = 32'd1; 
32'd97: dataIn2 = 32'd1; 
32'd98: dataIn2 = 32'd1; 
32'd99: dataIn2 = 32'd0; 
32'd100: dataIn2 = 32'd1; 
32'd101: dataIn2 = 32'd1; 
32'd102: dataIn2 = 32'd0; 
32'd103: dataIn2 = 32'd0; 
32'd104: dataIn2 = 32'd1; 
32'd105: dataIn2 = 32'd1; 
32'd106: dataIn2 = 32'd1; 
32'd107: dataIn2 = 32'd0; 
32'd108: dataIn2 = 32'd0; 
32'd109: dataIn2 = 32'd1; 
32'd110: dataIn2 = 32'd1; 
32'd111: dataIn2 = 32'd1; 
32'd112: dataIn2 = 32'd1; 
32'd113: dataIn2 = 32'd1; 
32'd114: dataIn2 = 32'd0; 
32'd115: dataIn2 = 32'd0; 
32'd116: dataIn2 = 32'd0; 
32'd117: dataIn2 = 32'd0; 
32'd118: dataIn2 = 32'd1; 
32'd119: dataIn2 = 32'd1; 
32'd120: dataIn2 = 32'd1; 
32'd121: dataIn2 = 32'd0; 
32'd122: dataIn2 = 32'd0; 
32'd123: dataIn2 = 32'd0; 
32'd124: dataIn2 = 32'd1; 
32'd125: dataIn2 = 32'd0; 
32'd126: dataIn2 = 32'd0; 
32'd127: dataIn2 = 32'd1; 
32'd128: dataIn2 = 32'd0; 
32'd129: dataIn2 = 32'd0; 
32'd130: dataIn2 = 32'd0; 
32'd131: dataIn2 = 32'd0; 
32'd132: dataIn2 = 32'd1; 
32'd133: dataIn2 = 32'd0; 
32'd134: dataIn2 = 32'd0; 
32'd135: dataIn2 = 32'd1; 
32'd136: dataIn2 = 32'd1; 
32'd137: dataIn2 = 32'd1; 
32'd138: dataIn2 = 32'd1; 
32'd139: dataIn2 = 32'd1; 
32'd140: dataIn2 = 32'd0; 
32'd141: dataIn2 = 32'd0; 
32'd142: dataIn2 = 32'd0; 
32'd143: dataIn2 = 32'd1; 
32'd144: dataIn2 = 32'd0; 
32'd145: dataIn2 = 32'd1; 
32'd146: dataIn2 = 32'd1; 
32'd147: dataIn2 = 32'd0; 
32'd148: dataIn2 = 32'd1; 
32'd149: dataIn2 = 32'd0; 
32'd150: dataIn2 = 32'd1; 
32'd151: dataIn2 = 32'd0; 
32'd152: dataIn2 = 32'd1; 
32'd153: dataIn2 = 32'd1; 
32'd154: dataIn2 = 32'd1; 
32'd155: dataIn2 = 32'd1; 
32'd156: dataIn2 = 32'd1; 
32'd157: dataIn2 = 32'd1; 
32'd158: dataIn2 = 32'd1; 
32'd159: dataIn2 = 32'd1; 
32'd160: dataIn2 = 32'd0; 
32'd161: dataIn2 = 32'd0; 
32'd162: dataIn2 = 32'd0; 
32'd163: dataIn2 = 32'd0; 
32'd164: dataIn2 = 32'd0; 
32'd165: dataIn2 = 32'd0; 
32'd166: dataIn2 = 32'd0; 
32'd167: dataIn2 = 32'd0; 
32'd168: dataIn2 = 32'd0; 
32'd169: dataIn2 = 32'd1; 
32'd170: dataIn2 = 32'd0; 
32'd171: dataIn2 = 32'd1; 
32'd172: dataIn2 = 32'd1; 
32'd173: dataIn2 = 32'd1; 
32'd174: dataIn2 = 32'd1; 
32'd175: dataIn2 = 32'd1; 
32'd176: dataIn2 = 32'd0; 
32'd177: dataIn2 = 32'd0; 
32'd178: dataIn2 = 32'd1; 
32'd179: dataIn2 = 32'd1; 
32'd180: dataIn2 = 32'd0; 
32'd181: dataIn2 = 32'd1; 
32'd182: dataIn2 = 32'd0; 
32'd183: dataIn2 = 32'd0; 
32'd184: dataIn2 = 32'd0; 
32'd185: dataIn2 = 32'd1; 
32'd186: dataIn2 = 32'd0; 
32'd187: dataIn2 = 32'd1; 
32'd188: dataIn2 = 32'd1; 
32'd189: dataIn2 = 32'd0; 
32'd190: dataIn2 = 32'd1; 
32'd191: dataIn2 = 32'd1; 
32'd192: dataIn2 = 32'd1; 
32'd193: dataIn2 = 32'd0; 
32'd194: dataIn2 = 32'd0; 
32'd195: dataIn2 = 32'd1; 
32'd196: dataIn2 = 32'd0; 
32'd197: dataIn2 = 32'd1; 
32'd198: dataIn2 = 32'd0; 
32'd199: dataIn2 = 32'd1; 
32'd200: dataIn2 = 32'd0; 
32'd201: dataIn2 = 32'd0; 
32'd202: dataIn2 = 32'd1; 
32'd203: dataIn2 = 32'd1; 
32'd204: dataIn2 = 32'd1; 
32'd205: dataIn2 = 32'd1; 
32'd206: dataIn2 = 32'd1; 
32'd207: dataIn2 = 32'd1; 
32'd208: dataIn2 = 32'd1; 
32'd209: dataIn2 = 32'd1; 
32'd210: dataIn2 = 32'd1; 
32'd211: dataIn2 = 32'd1; 
32'd212: dataIn2 = 32'd1; 
32'd213: dataIn2 = 32'd1; 
32'd214: dataIn2 = 32'd1; 
32'd215: dataIn2 = 32'd1; 
32'd216: dataIn2 = 32'd1; 
32'd217: dataIn2 = 32'd0; 
32'd218: dataIn2 = 32'd1; 
32'd219: dataIn2 = 32'd0; 
32'd220: dataIn2 = 32'd1; 
32'd221: dataIn2 = 32'd1; 
32'd222: dataIn2 = 32'd0; 
32'd223: dataIn2 = 32'd1; 
32'd224: dataIn2 = 32'd0; 
32'd225: dataIn2 = 32'd1; 
32'd226: dataIn2 = 32'd0; 
32'd227: dataIn2 = 32'd0; 
32'd228: dataIn2 = 32'd0; 
32'd229: dataIn2 = 32'd0; 
32'd230: dataIn2 = 32'd0; 
32'd231: dataIn2 = 32'd1; 
32'd232: dataIn2 = 32'd0; 
32'd233: dataIn2 = 32'd0; 
32'd234: dataIn2 = 32'd0; 
32'd235: dataIn2 = 32'd1; 
32'd236: dataIn2 = 32'd1; 
32'd237: dataIn2 = 32'd1; 
32'd238: dataIn2 = 32'd0; 
32'd239: dataIn2 = 32'd0; 
32'd240: dataIn2 = 32'd0; 
32'd241: dataIn2 = 32'd1; 
32'd242: dataIn2 = 32'd0; 
32'd243: dataIn2 = 32'd0; 
32'd244: dataIn2 = 32'd0; 
32'd245: dataIn2 = 32'd1; 
32'd246: dataIn2 = 32'd1; 
32'd247: dataIn2 = 32'd1; 
32'd248: dataIn2 = 32'd1; 
32'd249: dataIn2 = 32'd0; 
32'd250: dataIn2 = 32'd1; 
32'd251: dataIn2 = 32'd1; 
32'd252: dataIn2 = 32'd0; 
32'd253: dataIn2 = 32'd1; 
32'd254: dataIn2 = 32'd1; 
32'd255: dataIn2 = 32'd1; 
32'd256: dataIn2 = 32'd1; 
32'd257: dataIn2 = 32'd0; 
32'd258: dataIn2 = 32'd0; 
32'd259: dataIn2 = 32'd0; 
32'd260: dataIn2 = 32'd0; 
32'd261: dataIn2 = 32'd0; 
32'd262: dataIn2 = 32'd1; 
32'd263: dataIn2 = 32'd1; 
32'd264: dataIn2 = 32'd1; 
32'd265: dataIn2 = 32'd0; 
32'd266: dataIn2 = 32'd0; 
32'd267: dataIn2 = 32'd0; 
32'd268: dataIn2 = 32'd1; 
32'd269: dataIn2 = 32'd0; 
32'd270: dataIn2 = 32'd1; 
32'd271: dataIn2 = 32'd1; 
32'd272: dataIn2 = 32'd0; 
32'd273: dataIn2 = 32'd0; 
32'd274: dataIn2 = 32'd0; 
32'd275: dataIn2 = 32'd1; 
32'd276: dataIn2 = 32'd0; 
32'd277: dataIn2 = 32'd0; 
32'd278: dataIn2 = 32'd0; 
32'd279: dataIn2 = 32'd0; 
32'd280: dataIn2 = 32'd0; 
32'd281: dataIn2 = 32'd0; 
32'd282: dataIn2 = 32'd0; 
32'd283: dataIn2 = 32'd0; 
32'd284: dataIn2 = 32'd0; 
32'd285: dataIn2 = 32'd1; 
32'd286: dataIn2 = 32'd1; 
32'd287: dataIn2 = 32'd0; 
32'd288: dataIn2 = 32'd0; 
32'd289: dataIn2 = 32'd0; 
32'd290: dataIn2 = 32'd0; 
32'd291: dataIn2 = 32'd0; 
32'd292: dataIn2 = 32'd1; 
32'd293: dataIn2 = 32'd0; 
32'd294: dataIn2 = 32'd0; 
32'd295: dataIn2 = 32'd0; 
32'd296: dataIn2 = 32'd1; 
32'd297: dataIn2 = 32'd0; 
32'd298: dataIn2 = 32'd0; 
32'd299: dataIn2 = 32'd0; 
32'd300: dataIn2 = 32'd0; 
32'd301: dataIn2 = 32'd0; 
32'd302: dataIn2 = 32'd0; 
32'd303: dataIn2 = 32'd1; 
32'd304: dataIn2 = 32'd1; 
32'd305: dataIn2 = 32'd0; 
32'd306: dataIn2 = 32'd1; 
32'd307: dataIn2 = 32'd0; 
32'd308: dataIn2 = 32'd1; 
32'd309: dataIn2 = 32'd1; 
32'd310: dataIn2 = 32'd0; 
32'd311: dataIn2 = 32'd0; 
32'd312: dataIn2 = 32'd0; 
32'd313: dataIn2 = 32'd1; 
32'd314: dataIn2 = 32'd0; 
32'd315: dataIn2 = 32'd1; 
32'd316: dataIn2 = 32'd0; 
32'd317: dataIn2 = 32'd0; 
32'd318: dataIn2 = 32'd0; 
32'd319: dataIn2 = 32'd0; 
32'd320: dataIn2 = 32'd1; 
32'd321: dataIn2 = 32'd1; 
32'd322: dataIn2 = 32'd1; 
32'd323: dataIn2 = 32'd0; 
32'd324: dataIn2 = 32'd1; 
32'd325: dataIn2 = 32'd1; 
32'd326: dataIn2 = 32'd0; 
32'd327: dataIn2 = 32'd1; 
32'd328: dataIn2 = 32'd0; 
32'd329: dataIn2 = 32'd0; 
32'd330: dataIn2 = 32'd0; 
32'd331: dataIn2 = 32'd1; 
32'd332: dataIn2 = 32'd1; 
32'd333: dataIn2 = 32'd1; 
32'd334: dataIn2 = 32'd1; 
32'd335: dataIn2 = 32'd0; 
32'd336: dataIn2 = 32'd1; 
32'd337: dataIn2 = 32'd1; 
32'd338: dataIn2 = 32'd0; 
32'd339: dataIn2 = 32'd1; 
32'd340: dataIn2 = 32'd0; 
32'd341: dataIn2 = 32'd1; 
32'd342: dataIn2 = 32'd1; 
32'd343: dataIn2 = 32'd0; 
32'd344: dataIn2 = 32'd1; 
32'd345: dataIn2 = 32'd0; 
32'd346: dataIn2 = 32'd1; 
32'd347: dataIn2 = 32'd0; 
32'd348: dataIn2 = 32'd0; 
32'd349: dataIn2 = 32'd1; 
32'd350: dataIn2 = 32'd1; 
32'd351: dataIn2 = 32'd1; 
32'd352: dataIn2 = 32'd1; 
32'd353: dataIn2 = 32'd1; 
32'd354: dataIn2 = 32'd1; 
32'd355: dataIn2 = 32'd0; 
32'd356: dataIn2 = 32'd0; 
32'd357: dataIn2 = 32'd1; 
32'd358: dataIn2 = 32'd0; 
32'd359: dataIn2 = 32'd0; 
32'd360: dataIn2 = 32'd0; 
32'd361: dataIn2 = 32'd0; 
32'd362: dataIn2 = 32'd1; 
32'd363: dataIn2 = 32'd0; 
32'd364: dataIn2 = 32'd1; 
32'd365: dataIn2 = 32'd0; 
32'd366: dataIn2 = 32'd0; 
32'd367: dataIn2 = 32'd0; 
32'd368: dataIn2 = 32'd0; 
32'd369: dataIn2 = 32'd1; 
32'd370: dataIn2 = 32'd0; 
32'd371: dataIn2 = 32'd1; 
32'd372: dataIn2 = 32'd1; 
32'd373: dataIn2 = 32'd1; 
32'd374: dataIn2 = 32'd1; 
32'd375: dataIn2 = 32'd0; 
32'd376: dataIn2 = 32'd0; 
32'd377: dataIn2 = 32'd1; 
32'd378: dataIn2 = 32'd0; 
32'd379: dataIn2 = 32'd1; 
32'd380: dataIn2 = 32'd0; 
32'd381: dataIn2 = 32'd1; 
32'd382: dataIn2 = 32'd0; 
32'd383: dataIn2 = 32'd1; 
32'd384: dataIn2 = 32'd0; 
32'd385: dataIn2 = 32'd1; 
32'd386: dataIn2 = 32'd0; 
32'd387: dataIn2 = 32'd1; 
32'd388: dataIn2 = 32'd0; 
32'd389: dataIn2 = 32'd0; 
32'd390: dataIn2 = 32'd0; 
32'd391: dataIn2 = 32'd1; 
32'd392: dataIn2 = 32'd1; 
32'd393: dataIn2 = 32'd0; 
32'd394: dataIn2 = 32'd1; 
32'd395: dataIn2 = 32'd1; 
32'd396: dataIn2 = 32'd0; 
32'd397: dataIn2 = 32'd1; 
32'd398: dataIn2 = 32'd1; 
32'd399: dataIn2 = 32'd0; 
32'd400: dataIn2 = 32'd1; 
32'd401: dataIn2 = 32'd1; 
32'd402: dataIn2 = 32'd0; 
32'd403: dataIn2 = 32'd0; 
32'd404: dataIn2 = 32'd0; 
32'd405: dataIn2 = 32'd0; 
32'd406: dataIn2 = 32'd0; 
32'd407: dataIn2 = 32'd1; 
32'd408: dataIn2 = 32'd1; 
32'd409: dataIn2 = 32'd0; 
32'd410: dataIn2 = 32'd1; 
32'd411: dataIn2 = 32'd0; 
32'd412: dataIn2 = 32'd0; 
32'd413: dataIn2 = 32'd1; 
32'd414: dataIn2 = 32'd1; 
32'd415: dataIn2 = 32'd0; 
32'd416: dataIn2 = 32'd0; 
32'd417: dataIn2 = 32'd1; 
32'd418: dataIn2 = 32'd0; 
32'd419: dataIn2 = 32'd1; 
32'd420: dataIn2 = 32'd0; 
32'd421: dataIn2 = 32'd1; 
32'd422: dataIn2 = 32'd0; 
32'd423: dataIn2 = 32'd0; 
32'd424: dataIn2 = 32'd1; 
32'd425: dataIn2 = 32'd0; 
32'd426: dataIn2 = 32'd0; 
32'd427: dataIn2 = 32'd0; 
32'd428: dataIn2 = 32'd1; 
32'd429: dataIn2 = 32'd1; 
32'd430: dataIn2 = 32'd1; 
32'd431: dataIn2 = 32'd1; 
32'd432: dataIn2 = 32'd0; 
32'd433: dataIn2 = 32'd0; 
32'd434: dataIn2 = 32'd0; 
32'd435: dataIn2 = 32'd1; 
32'd436: dataIn2 = 32'd1; 
32'd437: dataIn2 = 32'd1; 
32'd438: dataIn2 = 32'd0; 
32'd439: dataIn2 = 32'd0; 
32'd440: dataIn2 = 32'd1; 
32'd441: dataIn2 = 32'd0; 
32'd442: dataIn2 = 32'd0; 
32'd443: dataIn2 = 32'd1; 
32'd444: dataIn2 = 32'd0; 
32'd445: dataIn2 = 32'd1; 
32'd446: dataIn2 = 32'd0; 
32'd447: dataIn2 = 32'd1; 
32'd448: dataIn2 = 32'd0; 
32'd449: dataIn2 = 32'd0; 
32'd450: dataIn2 = 32'd1; 
32'd451: dataIn2 = 32'd1; 
32'd452: dataIn2 = 32'd1; 
32'd453: dataIn2 = 32'd1; 
32'd454: dataIn2 = 32'd0; 
32'd455: dataIn2 = 32'd1; 
32'd456: dataIn2 = 32'd0; 
32'd457: dataIn2 = 32'd0; 
32'd458: dataIn2 = 32'd0; 
32'd459: dataIn2 = 32'd0; 
32'd460: dataIn2 = 32'd0; 
32'd461: dataIn2 = 32'd1; 
32'd462: dataIn2 = 32'd1; 
32'd463: dataIn2 = 32'd1; 
32'd464: dataIn2 = 32'd1; 
32'd465: dataIn2 = 32'd0; 
32'd466: dataIn2 = 32'd0; 
32'd467: dataIn2 = 32'd1; 
32'd468: dataIn2 = 32'd1; 
32'd469: dataIn2 = 32'd0; 
32'd470: dataIn2 = 32'd0; 
32'd471: dataIn2 = 32'd0; 
32'd472: dataIn2 = 32'd1; 
32'd473: dataIn2 = 32'd1; 
32'd474: dataIn2 = 32'd1; 
32'd475: dataIn2 = 32'd1; 
32'd476: dataIn2 = 32'd0; 
32'd477: dataIn2 = 32'd1; 
32'd478: dataIn2 = 32'd0; 
32'd479: dataIn2 = 32'd0; 
32'd480: dataIn2 = 32'd1; 
32'd481: dataIn2 = 32'd1; 
32'd482: dataIn2 = 32'd0; 
32'd483: dataIn2 = 32'd1; 
32'd484: dataIn2 = 32'd0; 
32'd485: dataIn2 = 32'd1; 
32'd486: dataIn2 = 32'd1; 
32'd487: dataIn2 = 32'd0; 
32'd488: dataIn2 = 32'd0; 
32'd489: dataIn2 = 32'd1; 
32'd490: dataIn2 = 32'd1; 
32'd491: dataIn2 = 32'd1; 
32'd492: dataIn2 = 32'd0; 
32'd493: dataIn2 = 32'd1; 
32'd494: dataIn2 = 32'd1; 
32'd495: dataIn2 = 32'd0; 
32'd496: dataIn2 = 32'd0; 
32'd497: dataIn2 = 32'd0; 
32'd498: dataIn2 = 32'd0; 
32'd499: dataIn2 = 32'd0; 
32'd500: dataIn2 = 32'd0; 
32'd501: dataIn2 = 32'd0; 
32'd502: dataIn2 = 32'd1; 
32'd503: dataIn2 = 32'd0; 
32'd504: dataIn2 = 32'd0; 
32'd505: dataIn2 = 32'd1; 
32'd506: dataIn2 = 32'd0; 
32'd507: dataIn2 = 32'd1; 
32'd508: dataIn2 = 32'd0; 
32'd509: dataIn2 = 32'd0; 
32'd510: dataIn2 = 32'd0; 
32'd511: dataIn2 = 32'd1; 
32'd512: dataIn2 = 32'd1; 
32'd513: dataIn2 = 32'd1; 
32'd514: dataIn2 = 32'd1; 
32'd515: dataIn2 = 32'd1; 
32'd516: dataIn2 = 32'd0; 
32'd517: dataIn2 = 32'd0; 
32'd518: dataIn2 = 32'd1; 
32'd519: dataIn2 = 32'd1; 
32'd520: dataIn2 = 32'd1; 
32'd521: dataIn2 = 32'd1; 
32'd522: dataIn2 = 32'd0; 
32'd523: dataIn2 = 32'd0; 
32'd524: dataIn2 = 32'd0; 
32'd525: dataIn2 = 32'd1; 
32'd526: dataIn2 = 32'd0; 
32'd527: dataIn2 = 32'd0; 
32'd528: dataIn2 = 32'd0; 
32'd529: dataIn2 = 32'd1; 
32'd530: dataIn2 = 32'd1; 
32'd531: dataIn2 = 32'd1; 
32'd532: dataIn2 = 32'd0; 
32'd533: dataIn2 = 32'd1; 
32'd534: dataIn2 = 32'd1; 
32'd535: dataIn2 = 32'd1; 
32'd536: dataIn2 = 32'd0; 
32'd537: dataIn2 = 32'd1; 
32'd538: dataIn2 = 32'd0; 
32'd539: dataIn2 = 32'd0; 
32'd540: dataIn2 = 32'd0; 
32'd541: dataIn2 = 32'd0; 
32'd542: dataIn2 = 32'd0; 
32'd543: dataIn2 = 32'd0; 
32'd544: dataIn2 = 32'd1; 
32'd545: dataIn2 = 32'd1; 
32'd546: dataIn2 = 32'd1; 
32'd547: dataIn2 = 32'd0; 
32'd548: dataIn2 = 32'd0; 
32'd549: dataIn2 = 32'd1; 
32'd550: dataIn2 = 32'd1; 
32'd551: dataIn2 = 32'd1; 
32'd552: dataIn2 = 32'd1; 
32'd553: dataIn2 = 32'd1; 
32'd554: dataIn2 = 32'd1; 
32'd555: dataIn2 = 32'd0; 
32'd556: dataIn2 = 32'd0; 
32'd557: dataIn2 = 32'd0; 
32'd558: dataIn2 = 32'd0; 
32'd559: dataIn2 = 32'd0; 
32'd560: dataIn2 = 32'd0; 
32'd561: dataIn2 = 32'd1; 
32'd562: dataIn2 = 32'd1; 
32'd563: dataIn2 = 32'd1; 
32'd564: dataIn2 = 32'd0; 
32'd565: dataIn2 = 32'd0; 
32'd566: dataIn2 = 32'd0; 
32'd567: dataIn2 = 32'd0; 
32'd568: dataIn2 = 32'd0; 
32'd569: dataIn2 = 32'd0; 
32'd570: dataIn2 = 32'd0; 
32'd571: dataIn2 = 32'd1; 
32'd572: dataIn2 = 32'd0; 
32'd573: dataIn2 = 32'd1; 
32'd574: dataIn2 = 32'd1; 
32'd575: dataIn2 = 32'd0; 
32'd576: dataIn2 = 32'd0; 
32'd577: dataIn2 = 32'd0; 
32'd578: dataIn2 = 32'd0; 
32'd579: dataIn2 = 32'd1; 
32'd580: dataIn2 = 32'd0; 
32'd581: dataIn2 = 32'd1; 
32'd582: dataIn2 = 32'd0; 
32'd583: dataIn2 = 32'd1; 
32'd584: dataIn2 = 32'd0; 
32'd585: dataIn2 = 32'd1; 
32'd586: dataIn2 = 32'd0; 
32'd587: dataIn2 = 32'd1; 
32'd588: dataIn2 = 32'd0; 
32'd589: dataIn2 = 32'd0; 
32'd590: dataIn2 = 32'd1; 
32'd591: dataIn2 = 32'd0; 
32'd592: dataIn2 = 32'd0; 
32'd593: dataIn2 = 32'd1; 
32'd594: dataIn2 = 32'd0; 
32'd595: dataIn2 = 32'd1; 
32'd596: dataIn2 = 32'd0; 
32'd597: dataIn2 = 32'd0; 
32'd598: dataIn2 = 32'd0; 
32'd599: dataIn2 = 32'd0; 
32'd600: dataIn2 = 32'd0; 
32'd601: dataIn2 = 32'd0; 
32'd602: dataIn2 = 32'd0; 
32'd603: dataIn2 = 32'd0; 
32'd604: dataIn2 = 32'd0; 
32'd605: dataIn2 = 32'd0; 
32'd606: dataIn2 = 32'd1; 
32'd607: dataIn2 = 32'd0; 
32'd608: dataIn2 = 32'd0; 
32'd609: dataIn2 = 32'd0; 
32'd610: dataIn2 = 32'd0; 
32'd611: dataIn2 = 32'd0; 
32'd612: dataIn2 = 32'd1; 
32'd613: dataIn2 = 32'd0; 
32'd614: dataIn2 = 32'd1; 
32'd615: dataIn2 = 32'd1; 
32'd616: dataIn2 = 32'd1; 
32'd617: dataIn2 = 32'd0; 
32'd618: dataIn2 = 32'd1; 
32'd619: dataIn2 = 32'd0; 
32'd620: dataIn2 = 32'd0; 
32'd621: dataIn2 = 32'd1; 
32'd622: dataIn2 = 32'd0; 
32'd623: dataIn2 = 32'd1; 
32'd624: dataIn2 = 32'd1; 
32'd625: dataIn2 = 32'd1; 
32'd626: dataIn2 = 32'd1; 
32'd627: dataIn2 = 32'd0; 
32'd628: dataIn2 = 32'd0; 
32'd629: dataIn2 = 32'd0; 
32'd630: dataIn2 = 32'd0; 
32'd631: dataIn2 = 32'd0; 
32'd632: dataIn2 = 32'd0; 
32'd633: dataIn2 = 32'd1; 
32'd634: dataIn2 = 32'd0; 
32'd635: dataIn2 = 32'd1; 
32'd636: dataIn2 = 32'd0; 
32'd637: dataIn2 = 32'd0; 
32'd638: dataIn2 = 32'd0; 
32'd639: dataIn2 = 32'd1; 
32'd640: dataIn2 = 32'd1; 
32'd641: dataIn2 = 32'd0; 
32'd642: dataIn2 = 32'd0; 
32'd643: dataIn2 = 32'd1; 
32'd644: dataIn2 = 32'd1; 
32'd645: dataIn2 = 32'd0; 
32'd646: dataIn2 = 32'd1; 
32'd647: dataIn2 = 32'd0; 
32'd648: dataIn2 = 32'd1; 
32'd649: dataIn2 = 32'd0; 
32'd650: dataIn2 = 32'd0; 
32'd651: dataIn2 = 32'd0; 
32'd652: dataIn2 = 32'd0; 
32'd653: dataIn2 = 32'd0; 
32'd654: dataIn2 = 32'd1; 
32'd655: dataIn2 = 32'd1; 
32'd656: dataIn2 = 32'd1; 
32'd657: dataIn2 = 32'd0; 
32'd658: dataIn2 = 32'd1; 
32'd659: dataIn2 = 32'd1; 
32'd660: dataIn2 = 32'd1; 
32'd661: dataIn2 = 32'd1; 
32'd662: dataIn2 = 32'd0; 
32'd663: dataIn2 = 32'd0; 
32'd664: dataIn2 = 32'd0; 
32'd665: dataIn2 = 32'd1; 
32'd666: dataIn2 = 32'd1; 
32'd667: dataIn2 = 32'd0; 
32'd668: dataIn2 = 32'd1; 
32'd669: dataIn2 = 32'd0; 
32'd670: dataIn2 = 32'd1; 
32'd671: dataIn2 = 32'd1; 
32'd672: dataIn2 = 32'd0; 
32'd673: dataIn2 = 32'd0; 
32'd674: dataIn2 = 32'd1; 
32'd675: dataIn2 = 32'd1; 
32'd676: dataIn2 = 32'd1; 
32'd677: dataIn2 = 32'd1; 
32'd678: dataIn2 = 32'd0; 
32'd679: dataIn2 = 32'd0; 
32'd680: dataIn2 = 32'd1; 
32'd681: dataIn2 = 32'd1; 
32'd682: dataIn2 = 32'd1; 
32'd683: dataIn2 = 32'd0; 
32'd684: dataIn2 = 32'd1; 
32'd685: dataIn2 = 32'd1; 
32'd686: dataIn2 = 32'd0; 
default: 
	dataIn2 = 32'd99999; 
endcase 
end 
always begin 
#10 Clk = ~Clk; 
end 
//========== VCD ============ 
`ifdef VCD 
initial 
begin 
	$dumpfile("685_bus.vcd");  
	$dumpvars; 
end 
`endif 
//===========RTLVCD ========== 
`ifdef RTLVCD 
initial 
begin 
	$dumpfile("hht_rtl.vcd"); 
	$dumpvars; 
end 
`endif 
endmodule 
