//800x800 
// Code your testbench here 
// or browse Examples 
// Verilog test bench for HHT with buffer 
`timescale 1ns/1ps 
module testbench; 
  parameter V_SIZE = 9; 
  parameter COL_SIZE = 38352 ; 
reg Clk,Rst,WR,mem_init; 
reg [31:0] dataIn1,dataIn2,csize; 
reg [31:0]v_values_base; 
wire [31:0]addr1,addr2; 
wire [4:0] regaddr1,regaddr2; 
reg[31:0] cpu_addr;
wire hht;
wire [31:0]val[0:8]; 
reg [31:0]wdata_col_base; 
wire [31:0] dataOut; 
reg fe_init; 
reg wn,rn,RD; 
wire [4:0]adata; 
wire [31:0] rdata; 
 // Instantiate memory module 
//  memmodel m1 (addr,dataIn,dataOut,WR,Clk,Rst); 
//  mem_buffer m1 (dataOut, full, empty, Clk, Rst, wn, rn, dataIn); 
control t1 (Clk,wdata_col_base,v_values_base,addr1,addr2,dataIn1,dataIn2,Rst,RD,csize,cpu_addr,hht,regaddr1,regaddr2,rdata,adata); ;  
//frontend t1 (Clk,Rst,fe_init,wdata_col_base,data_req,dataIn,init, 
//{m_cols[0],m_cols[1],m_cols[2],m_cols[3],m_cols[4]}, 
//done,wn); 
initial begin 
Clk = 1'b0; 
  RD = 1'b1; 
 #15; 
Rst = 1'b0; 
cpu_addr = 32'd126;
  v_values_base = 32'd2; 
  wdata_col_base = 32'd8020 ; 
  csize = COL_SIZE; 
 fe_init = 1'b1; 
#15 Rst = 1'b1; 
// RD = 1'b0; 
// RD = 1'b1; 
 #7090000; 
$finish; 
end 
always @(*) begin 
//$display("%b,%b",t1.fe1.count,t1.fe1.vdata_req); 
case(addr1)  
32'd8020: dataIn1 = 32'd48
; 
32'd8021: dataIn1 = 32'd53
; 
32'd8022: dataIn1 = 32'd66
; 
32'd8023: dataIn1 = 32'd70
; 
32'd8024: dataIn1 = 32'd154
; 
32'd8025: dataIn1 = 32'd159
; 
32'd8026: dataIn1 = 32'd163
; 
32'd8027: dataIn1 = 32'd170
; 
32'd8028: dataIn1 = 32'd180
; 
32'd8029: dataIn1 = 32'd200
; 
32'd8030: dataIn1 = 32'd206
; 
32'd8031: dataIn1 = 32'd234
; 
32'd8032: dataIn1 = 32'd254
; 
32'd8033: dataIn1 = 32'd289
; 
32'd8034: dataIn1 = 32'd297
; 
32'd8035: dataIn1 = 32'd331
; 
32'd8036: dataIn1 = 32'd345
; 
32'd8037: dataIn1 = 32'd364
; 
32'd8038: dataIn1 = 32'd385
; 
32'd8039: dataIn1 = 32'd394
; 
32'd8040: dataIn1 = 32'd405
; 
32'd8041: dataIn1 = 32'd422
; 
32'd8042: dataIn1 = 32'd430
; 
32'd8043: dataIn1 = 32'd434
; 
32'd8044: dataIn1 = 32'd440
; 
32'd8045: dataIn1 = 32'd471
; 
32'd8046: dataIn1 = 32'd474
; 
32'd8047: dataIn1 = 32'd515
; 
32'd8048: dataIn1 = 32'd557
; 
32'd8049: dataIn1 = 32'd568
; 
32'd8050: dataIn1 = 32'd577
; 
32'd8051: dataIn1 = 32'd622
; 
32'd8052: dataIn1 = 32'd625
; 
32'd8053: dataIn1 = 32'd656
; 
32'd8054: dataIn1 = 32'd658
; 
32'd8055: dataIn1 = 32'd665
; 
32'd8056: dataIn1 = 32'd721
; 
32'd8057: dataIn1 = 32'd751
; 
32'd8058: dataIn1 = 32'd773
; 
32'd8059: dataIn1 = 32'd792
; 
32'd8060: dataIn1 = 32'd7
; 
32'd8061: dataIn1 = 32'd29
; 
32'd8062: dataIn1 = 32'd31
; 
32'd8063: dataIn1 = 32'd33
; 
32'd8064: dataIn1 = 32'd35
; 
32'd8065: dataIn1 = 32'd37
; 
32'd8066: dataIn1 = 32'd46
; 
32'd8067: dataIn1 = 32'd53
; 
32'd8068: dataIn1 = 32'd57
; 
32'd8069: dataIn1 = 32'd60
; 
32'd8070: dataIn1 = 32'd84
; 
32'd8071: dataIn1 = 32'd99
; 
32'd8072: dataIn1 = 32'd151
; 
32'd8073: dataIn1 = 32'd156
; 
32'd8074: dataIn1 = 32'd177
; 
32'd8075: dataIn1 = 32'd204
; 
32'd8076: dataIn1 = 32'd228
; 
32'd8077: dataIn1 = 32'd239
; 
32'd8078: dataIn1 = 32'd248
; 
32'd8079: dataIn1 = 32'd272
; 
32'd8080: dataIn1 = 32'd295
; 
32'd8081: dataIn1 = 32'd305
; 
32'd8082: dataIn1 = 32'd327
; 
32'd8083: dataIn1 = 32'd355
; 
32'd8084: dataIn1 = 32'd360
; 
32'd8085: dataIn1 = 32'd378
; 
32'd8086: dataIn1 = 32'd381
; 
32'd8087: dataIn1 = 32'd394
; 
32'd8088: dataIn1 = 32'd429
; 
32'd8089: dataIn1 = 32'd435
; 
32'd8090: dataIn1 = 32'd440
; 
32'd8091: dataIn1 = 32'd467
; 
32'd8092: dataIn1 = 32'd468
; 
32'd8093: dataIn1 = 32'd502
; 
32'd8094: dataIn1 = 32'd506
; 
32'd8095: dataIn1 = 32'd551
; 
32'd8096: dataIn1 = 32'd558
; 
32'd8097: dataIn1 = 32'd565
; 
32'd8098: dataIn1 = 32'd598
; 
32'd8099: dataIn1 = 32'd614
; 
32'd8100: dataIn1 = 32'd646
; 
32'd8101: dataIn1 = 32'd650
; 
32'd8102: dataIn1 = 32'd658
; 
32'd8103: dataIn1 = 32'd663
; 
32'd8104: dataIn1 = 32'd707
; 
32'd8105: dataIn1 = 32'd727
; 
32'd8106: dataIn1 = 32'd733
; 
32'd8107: dataIn1 = 32'd751
; 
32'd8108: dataIn1 = 32'd777
; 
32'd8109: dataIn1 = 32'd782
; 
32'd8110: dataIn1 = 32'd783
; 
32'd8111: dataIn1 = 32'd23
; 
32'd8112: dataIn1 = 32'd55
; 
32'd8113: dataIn1 = 32'd58
; 
32'd8114: dataIn1 = 32'd61
; 
32'd8115: dataIn1 = 32'd77
; 
32'd8116: dataIn1 = 32'd85
; 
32'd8117: dataIn1 = 32'd94
; 
32'd8118: dataIn1 = 32'd98
; 
32'd8119: dataIn1 = 32'd100
; 
32'd8120: dataIn1 = 32'd109
; 
32'd8121: dataIn1 = 32'd118
; 
32'd8122: dataIn1 = 32'd136
; 
32'd8123: dataIn1 = 32'd139
; 
32'd8124: dataIn1 = 32'd154
; 
32'd8125: dataIn1 = 32'd194
; 
32'd8126: dataIn1 = 32'd202
; 
32'd8127: dataIn1 = 32'd205
; 
32'd8128: dataIn1 = 32'd208
; 
32'd8129: dataIn1 = 32'd215
; 
32'd8130: dataIn1 = 32'd239
; 
32'd8131: dataIn1 = 32'd264
; 
32'd8132: dataIn1 = 32'd282
; 
32'd8133: dataIn1 = 32'd319
; 
32'd8134: dataIn1 = 32'd356
; 
32'd8135: dataIn1 = 32'd374
; 
32'd8136: dataIn1 = 32'd385
; 
32'd8137: dataIn1 = 32'd408
; 
32'd8138: dataIn1 = 32'd417
; 
32'd8139: dataIn1 = 32'd426
; 
32'd8140: dataIn1 = 32'd444
; 
32'd8141: dataIn1 = 32'd459
; 
32'd8142: dataIn1 = 32'd478
; 
32'd8143: dataIn1 = 32'd488
; 
32'd8144: dataIn1 = 32'd503
; 
32'd8145: dataIn1 = 32'd506
; 
32'd8146: dataIn1 = 32'd529
; 
32'd8147: dataIn1 = 32'd532
; 
32'd8148: dataIn1 = 32'd538
; 
32'd8149: dataIn1 = 32'd553
; 
32'd8150: dataIn1 = 32'd589
; 
32'd8151: dataIn1 = 32'd608
; 
32'd8152: dataIn1 = 32'd613
; 
32'd8153: dataIn1 = 32'd678
; 
32'd8154: dataIn1 = 32'd686
; 
32'd8155: dataIn1 = 32'd697
; 
32'd8156: dataIn1 = 32'd717
; 
32'd8157: dataIn1 = 32'd724
; 
32'd8158: dataIn1 = 32'd734
; 
32'd8159: dataIn1 = 32'd785
; 
32'd8160: dataIn1 = 32'd28
; 
32'd8161: dataIn1 = 32'd47
; 
32'd8162: dataIn1 = 32'd54
; 
32'd8163: dataIn1 = 32'd55
; 
32'd8164: dataIn1 = 32'd109
; 
32'd8165: dataIn1 = 32'd123
; 
32'd8166: dataIn1 = 32'd127
; 
32'd8167: dataIn1 = 32'd140
; 
32'd8168: dataIn1 = 32'd171
; 
32'd8169: dataIn1 = 32'd197
; 
32'd8170: dataIn1 = 32'd233
; 
32'd8171: dataIn1 = 32'd240
; 
32'd8172: dataIn1 = 32'd242
; 
32'd8173: dataIn1 = 32'd244
; 
32'd8174: dataIn1 = 32'd247
; 
32'd8175: dataIn1 = 32'd253
; 
32'd8176: dataIn1 = 32'd261
; 
32'd8177: dataIn1 = 32'd272
; 
32'd8178: dataIn1 = 32'd278
; 
32'd8179: dataIn1 = 32'd296
; 
32'd8180: dataIn1 = 32'd355
; 
32'd8181: dataIn1 = 32'd359
; 
32'd8182: dataIn1 = 32'd361
; 
32'd8183: dataIn1 = 32'd399
; 
32'd8184: dataIn1 = 32'd429
; 
32'd8185: dataIn1 = 32'd433
; 
32'd8186: dataIn1 = 32'd434
; 
32'd8187: dataIn1 = 32'd440
; 
32'd8188: dataIn1 = 32'd441
; 
32'd8189: dataIn1 = 32'd442
; 
32'd8190: dataIn1 = 32'd466
; 
32'd8191: dataIn1 = 32'd474
; 
32'd8192: dataIn1 = 32'd490
; 
32'd8193: dataIn1 = 32'd493
; 
32'd8194: dataIn1 = 32'd495
; 
32'd8195: dataIn1 = 32'd506
; 
32'd8196: dataIn1 = 32'd516
; 
32'd8197: dataIn1 = 32'd529
; 
32'd8198: dataIn1 = 32'd531
; 
32'd8199: dataIn1 = 32'd535
; 
32'd8200: dataIn1 = 32'd537
; 
32'd8201: dataIn1 = 32'd546
; 
32'd8202: dataIn1 = 32'd557
; 
32'd8203: dataIn1 = 32'd574
; 
32'd8204: dataIn1 = 32'd576
; 
32'd8205: dataIn1 = 32'd577
; 
32'd8206: dataIn1 = 32'd580
; 
32'd8207: dataIn1 = 32'd587
; 
32'd8208: dataIn1 = 32'd603
; 
32'd8209: dataIn1 = 32'd604
; 
32'd8210: dataIn1 = 32'd612
; 
32'd8211: dataIn1 = 32'd624
; 
32'd8212: dataIn1 = 32'd641
; 
32'd8213: dataIn1 = 32'd643
; 
32'd8214: dataIn1 = 32'd669
; 
32'd8215: dataIn1 = 32'd671
; 
32'd8216: dataIn1 = 32'd672
; 
32'd8217: dataIn1 = 32'd709
; 
32'd8218: dataIn1 = 32'd719
; 
32'd8219: dataIn1 = 32'd722
; 
32'd8220: dataIn1 = 32'd725
; 
32'd8221: dataIn1 = 32'd740
; 
32'd8222: dataIn1 = 32'd748
; 
32'd8223: dataIn1 = 32'd752
; 
32'd8224: dataIn1 = 32'd769
; 
32'd8225: dataIn1 = 32'd773
; 
32'd8226: dataIn1 = 32'd13
; 
32'd8227: dataIn1 = 32'd18
; 
32'd8228: dataIn1 = 32'd25
; 
32'd8229: dataIn1 = 32'd37
; 
32'd8230: dataIn1 = 32'd41
; 
32'd8231: dataIn1 = 32'd48
; 
32'd8232: dataIn1 = 32'd103
; 
32'd8233: dataIn1 = 32'd124
; 
32'd8234: dataIn1 = 32'd133
; 
32'd8235: dataIn1 = 32'd163
; 
32'd8236: dataIn1 = 32'd175
; 
32'd8237: dataIn1 = 32'd191
; 
32'd8238: dataIn1 = 32'd201
; 
32'd8239: dataIn1 = 32'd221
; 
32'd8240: dataIn1 = 32'd244
; 
32'd8241: dataIn1 = 32'd287
; 
32'd8242: dataIn1 = 32'd289
; 
32'd8243: dataIn1 = 32'd294
; 
32'd8244: dataIn1 = 32'd296
; 
32'd8245: dataIn1 = 32'd300
; 
32'd8246: dataIn1 = 32'd313
; 
32'd8247: dataIn1 = 32'd328
; 
32'd8248: dataIn1 = 32'd337
; 
32'd8249: dataIn1 = 32'd344
; 
32'd8250: dataIn1 = 32'd354
; 
32'd8251: dataIn1 = 32'd356
; 
32'd8252: dataIn1 = 32'd367
; 
32'd8253: dataIn1 = 32'd378
; 
32'd8254: dataIn1 = 32'd382
; 
32'd8255: dataIn1 = 32'd388
; 
32'd8256: dataIn1 = 32'd425
; 
32'd8257: dataIn1 = 32'd453
; 
32'd8258: dataIn1 = 32'd455
; 
32'd8259: dataIn1 = 32'd458
; 
32'd8260: dataIn1 = 32'd463
; 
32'd8261: dataIn1 = 32'd469
; 
32'd8262: dataIn1 = 32'd501
; 
32'd8263: dataIn1 = 32'd510
; 
32'd8264: dataIn1 = 32'd519
; 
32'd8265: dataIn1 = 32'd540
; 
32'd8266: dataIn1 = 32'd542
; 
32'd8267: dataIn1 = 32'd543
; 
32'd8268: dataIn1 = 32'd556
; 
32'd8269: dataIn1 = 32'd623
; 
32'd8270: dataIn1 = 32'd654
; 
32'd8271: dataIn1 = 32'd689
; 
32'd8272: dataIn1 = 32'd694
; 
32'd8273: dataIn1 = 32'd708
; 
32'd8274: dataIn1 = 32'd760
; 
32'd8275: dataIn1 = 32'd781
; 
32'd8276: dataIn1 = 32'd21
; 
32'd8277: dataIn1 = 32'd41
; 
32'd8278: dataIn1 = 32'd53
; 
32'd8279: dataIn1 = 32'd68
; 
32'd8280: dataIn1 = 32'd85
; 
32'd8281: dataIn1 = 32'd96
; 
32'd8282: dataIn1 = 32'd97
; 
32'd8283: dataIn1 = 32'd104
; 
32'd8284: dataIn1 = 32'd113
; 
32'd8285: dataIn1 = 32'd115
; 
32'd8286: dataIn1 = 32'd121
; 
32'd8287: dataIn1 = 32'd146
; 
32'd8288: dataIn1 = 32'd158
; 
32'd8289: dataIn1 = 32'd181
; 
32'd8290: dataIn1 = 32'd185
; 
32'd8291: dataIn1 = 32'd191
; 
32'd8292: dataIn1 = 32'd193
; 
32'd8293: dataIn1 = 32'd253
; 
32'd8294: dataIn1 = 32'd256
; 
32'd8295: dataIn1 = 32'd298
; 
32'd8296: dataIn1 = 32'd352
; 
32'd8297: dataIn1 = 32'd411
; 
32'd8298: dataIn1 = 32'd422
; 
32'd8299: dataIn1 = 32'd449
; 
32'd8300: dataIn1 = 32'd452
; 
32'd8301: dataIn1 = 32'd458
; 
32'd8302: dataIn1 = 32'd487
; 
32'd8303: dataIn1 = 32'd510
; 
32'd8304: dataIn1 = 32'd525
; 
32'd8305: dataIn1 = 32'd538
; 
32'd8306: dataIn1 = 32'd551
; 
32'd8307: dataIn1 = 32'd568
; 
32'd8308: dataIn1 = 32'd571
; 
32'd8309: dataIn1 = 32'd618
; 
32'd8310: dataIn1 = 32'd630
; 
32'd8311: dataIn1 = 32'd652
; 
32'd8312: dataIn1 = 32'd680
; 
32'd8313: dataIn1 = 32'd684
; 
32'd8314: dataIn1 = 32'd695
; 
32'd8315: dataIn1 = 32'd717
; 
32'd8316: dataIn1 = 32'd727
; 
32'd8317: dataIn1 = 32'd746
; 
32'd8318: dataIn1 = 32'd769
; 
32'd8319: dataIn1 = 32'd23
; 
32'd8320: dataIn1 = 32'd25
; 
32'd8321: dataIn1 = 32'd44
; 
32'd8322: dataIn1 = 32'd51
; 
32'd8323: dataIn1 = 32'd55
; 
32'd8324: dataIn1 = 32'd75
; 
32'd8325: dataIn1 = 32'd107
; 
32'd8326: dataIn1 = 32'd112
; 
32'd8327: dataIn1 = 32'd135
; 
32'd8328: dataIn1 = 32'd169
; 
32'd8329: dataIn1 = 32'd171
; 
32'd8330: dataIn1 = 32'd184
; 
32'd8331: dataIn1 = 32'd190
; 
32'd8332: dataIn1 = 32'd195
; 
32'd8333: dataIn1 = 32'd203
; 
32'd8334: dataIn1 = 32'd222
; 
32'd8335: dataIn1 = 32'd225
; 
32'd8336: dataIn1 = 32'd236
; 
32'd8337: dataIn1 = 32'd263
; 
32'd8338: dataIn1 = 32'd280
; 
32'd8339: dataIn1 = 32'd285
; 
32'd8340: dataIn1 = 32'd294
; 
32'd8341: dataIn1 = 32'd296
; 
32'd8342: dataIn1 = 32'd323
; 
32'd8343: dataIn1 = 32'd332
; 
32'd8344: dataIn1 = 32'd336
; 
32'd8345: dataIn1 = 32'd358
; 
32'd8346: dataIn1 = 32'd363
; 
32'd8347: dataIn1 = 32'd374
; 
32'd8348: dataIn1 = 32'd386
; 
32'd8349: dataIn1 = 32'd387
; 
32'd8350: dataIn1 = 32'd426
; 
32'd8351: dataIn1 = 32'd432
; 
32'd8352: dataIn1 = 32'd440
; 
32'd8353: dataIn1 = 32'd456
; 
32'd8354: dataIn1 = 32'd479
; 
32'd8355: dataIn1 = 32'd527
; 
32'd8356: dataIn1 = 32'd538
; 
32'd8357: dataIn1 = 32'd539
; 
32'd8358: dataIn1 = 32'd544
; 
32'd8359: dataIn1 = 32'd547
; 
32'd8360: dataIn1 = 32'd564
; 
32'd8361: dataIn1 = 32'd589
; 
32'd8362: dataIn1 = 32'd599
; 
32'd8363: dataIn1 = 32'd607
; 
32'd8364: dataIn1 = 32'd620
; 
32'd8365: dataIn1 = 32'd627
; 
32'd8366: dataIn1 = 32'd630
; 
32'd8367: dataIn1 = 32'd673
; 
32'd8368: dataIn1 = 32'd736
; 
32'd8369: dataIn1 = 32'd743
; 
32'd8370: dataIn1 = 32'd759
; 
32'd8371: dataIn1 = 32'd781
; 
32'd8372: dataIn1 = 32'd789
; 
32'd8373: dataIn1 = 32'd47
; 
32'd8374: dataIn1 = 32'd65
; 
32'd8375: dataIn1 = 32'd69
; 
32'd8376: dataIn1 = 32'd141
; 
32'd8377: dataIn1 = 32'd143
; 
32'd8378: dataIn1 = 32'd145
; 
32'd8379: dataIn1 = 32'd176
; 
32'd8380: dataIn1 = 32'd214
; 
32'd8381: dataIn1 = 32'd217
; 
32'd8382: dataIn1 = 32'd225
; 
32'd8383: dataIn1 = 32'd253
; 
32'd8384: dataIn1 = 32'd330
; 
32'd8385: dataIn1 = 32'd337
; 
32'd8386: dataIn1 = 32'd344
; 
32'd8387: dataIn1 = 32'd347
; 
32'd8388: dataIn1 = 32'd360
; 
32'd8389: dataIn1 = 32'd365
; 
32'd8390: dataIn1 = 32'd367
; 
32'd8391: dataIn1 = 32'd369
; 
32'd8392: dataIn1 = 32'd394
; 
32'd8393: dataIn1 = 32'd419
; 
32'd8394: dataIn1 = 32'd421
; 
32'd8395: dataIn1 = 32'd450
; 
32'd8396: dataIn1 = 32'd465
; 
32'd8397: dataIn1 = 32'd468
; 
32'd8398: dataIn1 = 32'd476
; 
32'd8399: dataIn1 = 32'd509
; 
32'd8400: dataIn1 = 32'd510
; 
32'd8401: dataIn1 = 32'd514
; 
32'd8402: dataIn1 = 32'd515
; 
32'd8403: dataIn1 = 32'd516
; 
32'd8404: dataIn1 = 32'd531
; 
32'd8405: dataIn1 = 32'd577
; 
32'd8406: dataIn1 = 32'd592
; 
32'd8407: dataIn1 = 32'd660
; 
32'd8408: dataIn1 = 32'd688
; 
32'd8409: dataIn1 = 32'd697
; 
32'd8410: dataIn1 = 32'd721
; 
32'd8411: dataIn1 = 32'd747
; 
32'd8412: dataIn1 = 32'd749
; 
32'd8413: dataIn1 = 32'd795
; 
32'd8414: dataIn1 = 32'd800
; 
32'd8415: dataIn1 = 32'd31
; 
32'd8416: dataIn1 = 32'd39
; 
32'd8417: dataIn1 = 32'd40
; 
32'd8418: dataIn1 = 32'd43
; 
32'd8419: dataIn1 = 32'd55
; 
32'd8420: dataIn1 = 32'd71
; 
32'd8421: dataIn1 = 32'd91
; 
32'd8422: dataIn1 = 32'd114
; 
32'd8423: dataIn1 = 32'd139
; 
32'd8424: dataIn1 = 32'd157
; 
32'd8425: dataIn1 = 32'd174
; 
32'd8426: dataIn1 = 32'd199
; 
32'd8427: dataIn1 = 32'd204
; 
32'd8428: dataIn1 = 32'd216
; 
32'd8429: dataIn1 = 32'd218
; 
32'd8430: dataIn1 = 32'd251
; 
32'd8431: dataIn1 = 32'd291
; 
32'd8432: dataIn1 = 32'd308
; 
32'd8433: dataIn1 = 32'd313
; 
32'd8434: dataIn1 = 32'd318
; 
32'd8435: dataIn1 = 32'd353
; 
32'd8436: dataIn1 = 32'd361
; 
32'd8437: dataIn1 = 32'd387
; 
32'd8438: dataIn1 = 32'd401
; 
32'd8439: dataIn1 = 32'd410
; 
32'd8440: dataIn1 = 32'd419
; 
32'd8441: dataIn1 = 32'd424
; 
32'd8442: dataIn1 = 32'd461
; 
32'd8443: dataIn1 = 32'd468
; 
32'd8444: dataIn1 = 32'd470
; 
32'd8445: dataIn1 = 32'd483
; 
32'd8446: dataIn1 = 32'd484
; 
32'd8447: dataIn1 = 32'd501
; 
32'd8448: dataIn1 = 32'd530
; 
32'd8449: dataIn1 = 32'd550
; 
32'd8450: dataIn1 = 32'd560
; 
32'd8451: dataIn1 = 32'd614
; 
32'd8452: dataIn1 = 32'd631
; 
32'd8453: dataIn1 = 32'd651
; 
32'd8454: dataIn1 = 32'd655
; 
32'd8455: dataIn1 = 32'd668
; 
32'd8456: dataIn1 = 32'd684
; 
32'd8457: dataIn1 = 32'd714
; 
32'd8458: dataIn1 = 32'd748
; 
32'd8459: dataIn1 = 32'd769
; 
32'd8460: dataIn1 = 32'd771
; 
32'd8461: dataIn1 = 32'd13
; 
32'd8462: dataIn1 = 32'd19
; 
32'd8463: dataIn1 = 32'd25
; 
32'd8464: dataIn1 = 32'd49
; 
32'd8465: dataIn1 = 32'd57
; 
32'd8466: dataIn1 = 32'd67
; 
32'd8467: dataIn1 = 32'd105
; 
32'd8468: dataIn1 = 32'd116
; 
32'd8469: dataIn1 = 32'd144
; 
32'd8470: dataIn1 = 32'd145
; 
32'd8471: dataIn1 = 32'd152
; 
32'd8472: dataIn1 = 32'd158
; 
32'd8473: dataIn1 = 32'd184
; 
32'd8474: dataIn1 = 32'd194
; 
32'd8475: dataIn1 = 32'd200
; 
32'd8476: dataIn1 = 32'd204
; 
32'd8477: dataIn1 = 32'd213
; 
32'd8478: dataIn1 = 32'd222
; 
32'd8479: dataIn1 = 32'd234
; 
32'd8480: dataIn1 = 32'd240
; 
32'd8481: dataIn1 = 32'd241
; 
32'd8482: dataIn1 = 32'd243
; 
32'd8483: dataIn1 = 32'd253
; 
32'd8484: dataIn1 = 32'd254
; 
32'd8485: dataIn1 = 32'd384
; 
32'd8486: dataIn1 = 32'd392
; 
32'd8487: dataIn1 = 32'd421
; 
32'd8488: dataIn1 = 32'd432
; 
32'd8489: dataIn1 = 32'd441
; 
32'd8490: dataIn1 = 32'd471
; 
32'd8491: dataIn1 = 32'd486
; 
32'd8492: dataIn1 = 32'd530
; 
32'd8493: dataIn1 = 32'd568
; 
32'd8494: dataIn1 = 32'd617
; 
32'd8495: dataIn1 = 32'd679
; 
32'd8496: dataIn1 = 32'd688
; 
32'd8497: dataIn1 = 32'd695
; 
32'd8498: dataIn1 = 32'd697
; 
32'd8499: dataIn1 = 32'd793
; 
32'd8500: dataIn1 = 32'd26
; 
32'd8501: dataIn1 = 32'd27
; 
32'd8502: dataIn1 = 32'd44
; 
32'd8503: dataIn1 = 32'd49
; 
32'd8504: dataIn1 = 32'd78
; 
32'd8505: dataIn1 = 32'd86
; 
32'd8506: dataIn1 = 32'd97
; 
32'd8507: dataIn1 = 32'd124
; 
32'd8508: dataIn1 = 32'd156
; 
32'd8509: dataIn1 = 32'd182
; 
32'd8510: dataIn1 = 32'd234
; 
32'd8511: dataIn1 = 32'd260
; 
32'd8512: dataIn1 = 32'd279
; 
32'd8513: dataIn1 = 32'd281
; 
32'd8514: dataIn1 = 32'd296
; 
32'd8515: dataIn1 = 32'd335
; 
32'd8516: dataIn1 = 32'd352
; 
32'd8517: dataIn1 = 32'd366
; 
32'd8518: dataIn1 = 32'd368
; 
32'd8519: dataIn1 = 32'd376
; 
32'd8520: dataIn1 = 32'd390
; 
32'd8521: dataIn1 = 32'd406
; 
32'd8522: dataIn1 = 32'd416
; 
32'd8523: dataIn1 = 32'd440
; 
32'd8524: dataIn1 = 32'd465
; 
32'd8525: dataIn1 = 32'd471
; 
32'd8526: dataIn1 = 32'd472
; 
32'd8527: dataIn1 = 32'd486
; 
32'd8528: dataIn1 = 32'd489
; 
32'd8529: dataIn1 = 32'd531
; 
32'd8530: dataIn1 = 32'd550
; 
32'd8531: dataIn1 = 32'd576
; 
32'd8532: dataIn1 = 32'd579
; 
32'd8533: dataIn1 = 32'd590
; 
32'd8534: dataIn1 = 32'd633
; 
32'd8535: dataIn1 = 32'd674
; 
32'd8536: dataIn1 = 32'd701
; 
32'd8537: dataIn1 = 32'd720
; 
32'd8538: dataIn1 = 32'd748
; 
32'd8539: dataIn1 = 32'd773
; 
32'd8540: dataIn1 = 32'd777
; 
32'd8541: dataIn1 = 32'd785
; 
32'd8542: dataIn1 = 32'd792
; 
32'd8543: dataIn1 = 32'd16
; 
32'd8544: dataIn1 = 32'd18
; 
32'd8545: dataIn1 = 32'd59
; 
32'd8546: dataIn1 = 32'd64
; 
32'd8547: dataIn1 = 32'd76
; 
32'd8548: dataIn1 = 32'd101
; 
32'd8549: dataIn1 = 32'd105
; 
32'd8550: dataIn1 = 32'd126
; 
32'd8551: dataIn1 = 32'd143
; 
32'd8552: dataIn1 = 32'd145
; 
32'd8553: dataIn1 = 32'd207
; 
32'd8554: dataIn1 = 32'd212
; 
32'd8555: dataIn1 = 32'd229
; 
32'd8556: dataIn1 = 32'd251
; 
32'd8557: dataIn1 = 32'd261
; 
32'd8558: dataIn1 = 32'd262
; 
32'd8559: dataIn1 = 32'd268
; 
32'd8560: dataIn1 = 32'd283
; 
32'd8561: dataIn1 = 32'd307
; 
32'd8562: dataIn1 = 32'd337
; 
32'd8563: dataIn1 = 32'd338
; 
32'd8564: dataIn1 = 32'd349
; 
32'd8565: dataIn1 = 32'd357
; 
32'd8566: dataIn1 = 32'd396
; 
32'd8567: dataIn1 = 32'd397
; 
32'd8568: dataIn1 = 32'd408
; 
32'd8569: dataIn1 = 32'd417
; 
32'd8570: dataIn1 = 32'd432
; 
32'd8571: dataIn1 = 32'd439
; 
32'd8572: dataIn1 = 32'd459
; 
32'd8573: dataIn1 = 32'd464
; 
32'd8574: dataIn1 = 32'd491
; 
32'd8575: dataIn1 = 32'd493
; 
32'd8576: dataIn1 = 32'd515
; 
32'd8577: dataIn1 = 32'd554
; 
32'd8578: dataIn1 = 32'd586
; 
32'd8579: dataIn1 = 32'd601
; 
32'd8580: dataIn1 = 32'd662
; 
32'd8581: dataIn1 = 32'd664
; 
32'd8582: dataIn1 = 32'd694
; 
32'd8583: dataIn1 = 32'd706
; 
32'd8584: dataIn1 = 32'd743
; 
32'd8585: dataIn1 = 32'd748
; 
32'd8586: dataIn1 = 32'd754
; 
32'd8587: dataIn1 = 32'd771
; 
32'd8588: dataIn1 = 32'd781
; 
32'd8589: dataIn1 = 32'd792
; 
32'd8590: dataIn1 = 32'd61
; 
32'd8591: dataIn1 = 32'd62
; 
32'd8592: dataIn1 = 32'd75
; 
32'd8593: dataIn1 = 32'd111
; 
32'd8594: dataIn1 = 32'd118
; 
32'd8595: dataIn1 = 32'd142
; 
32'd8596: dataIn1 = 32'd148
; 
32'd8597: dataIn1 = 32'd159
; 
32'd8598: dataIn1 = 32'd176
; 
32'd8599: dataIn1 = 32'd198
; 
32'd8600: dataIn1 = 32'd202
; 
32'd8601: dataIn1 = 32'd223
; 
32'd8602: dataIn1 = 32'd226
; 
32'd8603: dataIn1 = 32'd227
; 
32'd8604: dataIn1 = 32'd279
; 
32'd8605: dataIn1 = 32'd280
; 
32'd8606: dataIn1 = 32'd316
; 
32'd8607: dataIn1 = 32'd343
; 
32'd8608: dataIn1 = 32'd361
; 
32'd8609: dataIn1 = 32'd392
; 
32'd8610: dataIn1 = 32'd396
; 
32'd8611: dataIn1 = 32'd423
; 
32'd8612: dataIn1 = 32'd428
; 
32'd8613: dataIn1 = 32'd440
; 
32'd8614: dataIn1 = 32'd450
; 
32'd8615: dataIn1 = 32'd451
; 
32'd8616: dataIn1 = 32'd469
; 
32'd8617: dataIn1 = 32'd499
; 
32'd8618: dataIn1 = 32'd557
; 
32'd8619: dataIn1 = 32'd574
; 
32'd8620: dataIn1 = 32'd577
; 
32'd8621: dataIn1 = 32'd600
; 
32'd8622: dataIn1 = 32'd606
; 
32'd8623: dataIn1 = 32'd653
; 
32'd8624: dataIn1 = 32'd658
; 
32'd8625: dataIn1 = 32'd685
; 
32'd8626: dataIn1 = 32'd689
; 
32'd8627: dataIn1 = 32'd693
; 
32'd8628: dataIn1 = 32'd697
; 
32'd8629: dataIn1 = 32'd753
; 
32'd8630: dataIn1 = 32'd765
; 
32'd8631: dataIn1 = 32'd771
; 
32'd8632: dataIn1 = 32'd779
; 
32'd8633: dataIn1 = 32'd785
; 
32'd8634: dataIn1 = 32'd793
; 
32'd8635: dataIn1 = 32'd19
; 
32'd8636: dataIn1 = 32'd42
; 
32'd8637: dataIn1 = 32'd49
; 
32'd8638: dataIn1 = 32'd57
; 
32'd8639: dataIn1 = 32'd67
; 
32'd8640: dataIn1 = 32'd96
; 
32'd8641: dataIn1 = 32'd97
; 
32'd8642: dataIn1 = 32'd99
; 
32'd8643: dataIn1 = 32'd135
; 
32'd8644: dataIn1 = 32'd160
; 
32'd8645: dataIn1 = 32'd184
; 
32'd8646: dataIn1 = 32'd206
; 
32'd8647: dataIn1 = 32'd207
; 
32'd8648: dataIn1 = 32'd215
; 
32'd8649: dataIn1 = 32'd225
; 
32'd8650: dataIn1 = 32'd242
; 
32'd8651: dataIn1 = 32'd289
; 
32'd8652: dataIn1 = 32'd303
; 
32'd8653: dataIn1 = 32'd314
; 
32'd8654: dataIn1 = 32'd340
; 
32'd8655: dataIn1 = 32'd346
; 
32'd8656: dataIn1 = 32'd351
; 
32'd8657: dataIn1 = 32'd353
; 
32'd8658: dataIn1 = 32'd356
; 
32'd8659: dataIn1 = 32'd364
; 
32'd8660: dataIn1 = 32'd366
; 
32'd8661: dataIn1 = 32'd386
; 
32'd8662: dataIn1 = 32'd396
; 
32'd8663: dataIn1 = 32'd444
; 
32'd8664: dataIn1 = 32'd466
; 
32'd8665: dataIn1 = 32'd472
; 
32'd8666: dataIn1 = 32'd488
; 
32'd8667: dataIn1 = 32'd491
; 
32'd8668: dataIn1 = 32'd550
; 
32'd8669: dataIn1 = 32'd565
; 
32'd8670: dataIn1 = 32'd580
; 
32'd8671: dataIn1 = 32'd595
; 
32'd8672: dataIn1 = 32'd600
; 
32'd8673: dataIn1 = 32'd604
; 
32'd8674: dataIn1 = 32'd607
; 
32'd8675: dataIn1 = 32'd653
; 
32'd8676: dataIn1 = 32'd658
; 
32'd8677: dataIn1 = 32'd677
; 
32'd8678: dataIn1 = 32'd723
; 
32'd8679: dataIn1 = 32'd725
; 
32'd8680: dataIn1 = 32'd732
; 
32'd8681: dataIn1 = 32'd733
; 
32'd8682: dataIn1 = 32'd741
; 
32'd8683: dataIn1 = 32'd742
; 
32'd8684: dataIn1 = 32'd750
; 
32'd8685: dataIn1 = 32'd759
; 
32'd8686: dataIn1 = 32'd34
; 
32'd8687: dataIn1 = 32'd69
; 
32'd8688: dataIn1 = 32'd81
; 
32'd8689: dataIn1 = 32'd83
; 
32'd8690: dataIn1 = 32'd85
; 
32'd8691: dataIn1 = 32'd89
; 
32'd8692: dataIn1 = 32'd98
; 
32'd8693: dataIn1 = 32'd109
; 
32'd8694: dataIn1 = 32'd111
; 
32'd8695: dataIn1 = 32'd130
; 
32'd8696: dataIn1 = 32'd154
; 
32'd8697: dataIn1 = 32'd155
; 
32'd8698: dataIn1 = 32'd156
; 
32'd8699: dataIn1 = 32'd162
; 
32'd8700: dataIn1 = 32'd182
; 
32'd8701: dataIn1 = 32'd190
; 
32'd8702: dataIn1 = 32'd191
; 
32'd8703: dataIn1 = 32'd194
; 
32'd8704: dataIn1 = 32'd207
; 
32'd8705: dataIn1 = 32'd285
; 
32'd8706: dataIn1 = 32'd315
; 
32'd8707: dataIn1 = 32'd353
; 
32'd8708: dataIn1 = 32'd371
; 
32'd8709: dataIn1 = 32'd397
; 
32'd8710: dataIn1 = 32'd432
; 
32'd8711: dataIn1 = 32'd468
; 
32'd8712: dataIn1 = 32'd500
; 
32'd8713: dataIn1 = 32'd511
; 
32'd8714: dataIn1 = 32'd513
; 
32'd8715: dataIn1 = 32'd535
; 
32'd8716: dataIn1 = 32'd559
; 
32'd8717: dataIn1 = 32'd576
; 
32'd8718: dataIn1 = 32'd603
; 
32'd8719: dataIn1 = 32'd615
; 
32'd8720: dataIn1 = 32'd616
; 
32'd8721: dataIn1 = 32'd648
; 
32'd8722: dataIn1 = 32'd650
; 
32'd8723: dataIn1 = 32'd660
; 
32'd8724: dataIn1 = 32'd683
; 
32'd8725: dataIn1 = 32'd692
; 
32'd8726: dataIn1 = 32'd727
; 
32'd8727: dataIn1 = 32'd731
; 
32'd8728: dataIn1 = 32'd737
; 
32'd8729: dataIn1 = 32'd740
; 
32'd8730: dataIn1 = 32'd744
; 
32'd8731: dataIn1 = 32'd751
; 
32'd8732: dataIn1 = 32'd784
; 
32'd8733: dataIn1 = 32'd786
; 
32'd8734: dataIn1 = 32'd794
; 
32'd8735: dataIn1 = 32'd70
; 
32'd8736: dataIn1 = 32'd73
; 
32'd8737: dataIn1 = 32'd76
; 
32'd8738: dataIn1 = 32'd84
; 
32'd8739: dataIn1 = 32'd97
; 
32'd8740: dataIn1 = 32'd102
; 
32'd8741: dataIn1 = 32'd107
; 
32'd8742: dataIn1 = 32'd118
; 
32'd8743: dataIn1 = 32'd120
; 
32'd8744: dataIn1 = 32'd153
; 
32'd8745: dataIn1 = 32'd191
; 
32'd8746: dataIn1 = 32'd216
; 
32'd8747: dataIn1 = 32'd228
; 
32'd8748: dataIn1 = 32'd234
; 
32'd8749: dataIn1 = 32'd235
; 
32'd8750: dataIn1 = 32'd269
; 
32'd8751: dataIn1 = 32'd276
; 
32'd8752: dataIn1 = 32'd330
; 
32'd8753: dataIn1 = 32'd360
; 
32'd8754: dataIn1 = 32'd364
; 
32'd8755: dataIn1 = 32'd380
; 
32'd8756: dataIn1 = 32'd389
; 
32'd8757: dataIn1 = 32'd400
; 
32'd8758: dataIn1 = 32'd412
; 
32'd8759: dataIn1 = 32'd426
; 
32'd8760: dataIn1 = 32'd428
; 
32'd8761: dataIn1 = 32'd454
; 
32'd8762: dataIn1 = 32'd461
; 
32'd8763: dataIn1 = 32'd481
; 
32'd8764: dataIn1 = 32'd515
; 
32'd8765: dataIn1 = 32'd558
; 
32'd8766: dataIn1 = 32'd607
; 
32'd8767: dataIn1 = 32'd613
; 
32'd8768: dataIn1 = 32'd616
; 
32'd8769: dataIn1 = 32'd619
; 
32'd8770: dataIn1 = 32'd621
; 
32'd8771: dataIn1 = 32'd626
; 
32'd8772: dataIn1 = 32'd637
; 
32'd8773: dataIn1 = 32'd690
; 
32'd8774: dataIn1 = 32'd699
; 
32'd8775: dataIn1 = 32'd704
; 
32'd8776: dataIn1 = 32'd707
; 
32'd8777: dataIn1 = 32'd760
; 
32'd8778: dataIn1 = 32'd781
; 
32'd8779: dataIn1 = 32'd784
; 
32'd8780: dataIn1 = 32'd29
; 
32'd8781: dataIn1 = 32'd30
; 
32'd8782: dataIn1 = 32'd33
; 
32'd8783: dataIn1 = 32'd54
; 
32'd8784: dataIn1 = 32'd83
; 
32'd8785: dataIn1 = 32'd85
; 
32'd8786: dataIn1 = 32'd139
; 
32'd8787: dataIn1 = 32'd213
; 
32'd8788: dataIn1 = 32'd225
; 
32'd8789: dataIn1 = 32'd248
; 
32'd8790: dataIn1 = 32'd277
; 
32'd8791: dataIn1 = 32'd305
; 
32'd8792: dataIn1 = 32'd319
; 
32'd8793: dataIn1 = 32'd336
; 
32'd8794: dataIn1 = 32'd355
; 
32'd8795: dataIn1 = 32'd363
; 
32'd8796: dataIn1 = 32'd408
; 
32'd8797: dataIn1 = 32'd412
; 
32'd8798: dataIn1 = 32'd427
; 
32'd8799: dataIn1 = 32'd485
; 
32'd8800: dataIn1 = 32'd491
; 
32'd8801: dataIn1 = 32'd494
; 
32'd8802: dataIn1 = 32'd554
; 
32'd8803: dataIn1 = 32'd585
; 
32'd8804: dataIn1 = 32'd635
; 
32'd8805: dataIn1 = 32'd638
; 
32'd8806: dataIn1 = 32'd655
; 
32'd8807: dataIn1 = 32'd665
; 
32'd8808: dataIn1 = 32'd667
; 
32'd8809: dataIn1 = 32'd679
; 
32'd8810: dataIn1 = 32'd696
; 
32'd8811: dataIn1 = 32'd716
; 
32'd8812: dataIn1 = 32'd738
; 
32'd8813: dataIn1 = 32'd762
; 
32'd8814: dataIn1 = 32'd786
; 
32'd8815: dataIn1 = 32'd800
; 
32'd8816: dataIn1 = 32'd21
; 
32'd8817: dataIn1 = 32'd30
; 
32'd8818: dataIn1 = 32'd58
; 
32'd8819: dataIn1 = 32'd78
; 
32'd8820: dataIn1 = 32'd86
; 
32'd8821: dataIn1 = 32'd94
; 
32'd8822: dataIn1 = 32'd113
; 
32'd8823: dataIn1 = 32'd121
; 
32'd8824: dataIn1 = 32'd185
; 
32'd8825: dataIn1 = 32'd232
; 
32'd8826: dataIn1 = 32'd238
; 
32'd8827: dataIn1 = 32'd291
; 
32'd8828: dataIn1 = 32'd333
; 
32'd8829: dataIn1 = 32'd336
; 
32'd8830: dataIn1 = 32'd363
; 
32'd8831: dataIn1 = 32'd373
; 
32'd8832: dataIn1 = 32'd415
; 
32'd8833: dataIn1 = 32'd427
; 
32'd8834: dataIn1 = 32'd476
; 
32'd8835: dataIn1 = 32'd477
; 
32'd8836: dataIn1 = 32'd494
; 
32'd8837: dataIn1 = 32'd510
; 
32'd8838: dataIn1 = 32'd533
; 
32'd8839: dataIn1 = 32'd534
; 
32'd8840: dataIn1 = 32'd547
; 
32'd8841: dataIn1 = 32'd552
; 
32'd8842: dataIn1 = 32'd573
; 
32'd8843: dataIn1 = 32'd592
; 
32'd8844: dataIn1 = 32'd607
; 
32'd8845: dataIn1 = 32'd620
; 
32'd8846: dataIn1 = 32'd635
; 
32'd8847: dataIn1 = 32'd641
; 
32'd8848: dataIn1 = 32'd642
; 
32'd8849: dataIn1 = 32'd664
; 
32'd8850: dataIn1 = 32'd667
; 
32'd8851: dataIn1 = 32'd668
; 
32'd8852: dataIn1 = 32'd715
; 
32'd8853: dataIn1 = 32'd734
; 
32'd8854: dataIn1 = 32'd736
; 
32'd8855: dataIn1 = 32'd784
; 
32'd8856: dataIn1 = 32'd793
; 
32'd8857: dataIn1 = 32'd800
; 
32'd8858: dataIn1 = 32'd29
; 
32'd8859: dataIn1 = 32'd35
; 
32'd8860: dataIn1 = 32'd39
; 
32'd8861: dataIn1 = 32'd42
; 
32'd8862: dataIn1 = 32'd84
; 
32'd8863: dataIn1 = 32'd96
; 
32'd8864: dataIn1 = 32'd108
; 
32'd8865: dataIn1 = 32'd162
; 
32'd8866: dataIn1 = 32'd202
; 
32'd8867: dataIn1 = 32'd235
; 
32'd8868: dataIn1 = 32'd249
; 
32'd8869: dataIn1 = 32'd250
; 
32'd8870: dataIn1 = 32'd281
; 
32'd8871: dataIn1 = 32'd324
; 
32'd8872: dataIn1 = 32'd342
; 
32'd8873: dataIn1 = 32'd349
; 
32'd8874: dataIn1 = 32'd351
; 
32'd8875: dataIn1 = 32'd363
; 
32'd8876: dataIn1 = 32'd395
; 
32'd8877: dataIn1 = 32'd400
; 
32'd8878: dataIn1 = 32'd439
; 
32'd8879: dataIn1 = 32'd445
; 
32'd8880: dataIn1 = 32'd478
; 
32'd8881: dataIn1 = 32'd484
; 
32'd8882: dataIn1 = 32'd500
; 
32'd8883: dataIn1 = 32'd510
; 
32'd8884: dataIn1 = 32'd522
; 
32'd8885: dataIn1 = 32'd538
; 
32'd8886: dataIn1 = 32'd541
; 
32'd8887: dataIn1 = 32'd548
; 
32'd8888: dataIn1 = 32'd552
; 
32'd8889: dataIn1 = 32'd556
; 
32'd8890: dataIn1 = 32'd618
; 
32'd8891: dataIn1 = 32'd654
; 
32'd8892: dataIn1 = 32'd655
; 
32'd8893: dataIn1 = 32'd670
; 
32'd8894: dataIn1 = 32'd699
; 
32'd8895: dataIn1 = 32'd772
; 
32'd8896: dataIn1 = 32'd777
; 
32'd8897: dataIn1 = 32'd799
; 
32'd8898: dataIn1 = 32'd41
; 
32'd8899: dataIn1 = 32'd86
; 
32'd8900: dataIn1 = 32'd128
; 
32'd8901: dataIn1 = 32'd199
; 
32'd8902: dataIn1 = 32'd205
; 
32'd8903: dataIn1 = 32'd215
; 
32'd8904: dataIn1 = 32'd236
; 
32'd8905: dataIn1 = 32'd249
; 
32'd8906: dataIn1 = 32'd270
; 
32'd8907: dataIn1 = 32'd274
; 
32'd8908: dataIn1 = 32'd289
; 
32'd8909: dataIn1 = 32'd455
; 
32'd8910: dataIn1 = 32'd458
; 
32'd8911: dataIn1 = 32'd492
; 
32'd8912: dataIn1 = 32'd502
; 
32'd8913: dataIn1 = 32'd539
; 
32'd8914: dataIn1 = 32'd550
; 
32'd8915: dataIn1 = 32'd568
; 
32'd8916: dataIn1 = 32'd569
; 
32'd8917: dataIn1 = 32'd586
; 
32'd8918: dataIn1 = 32'd594
; 
32'd8919: dataIn1 = 32'd601
; 
32'd8920: dataIn1 = 32'd636
; 
32'd8921: dataIn1 = 32'd649
; 
32'd8922: dataIn1 = 32'd650
; 
32'd8923: dataIn1 = 32'd653
; 
32'd8924: dataIn1 = 32'd660
; 
32'd8925: dataIn1 = 32'd709
; 
32'd8926: dataIn1 = 32'd712
; 
32'd8927: dataIn1 = 32'd741
; 
32'd8928: dataIn1 = 32'd751
; 
32'd8929: dataIn1 = 32'd760
; 
32'd8930: dataIn1 = 32'd763
; 
32'd8931: dataIn1 = 32'd34
; 
32'd8932: dataIn1 = 32'd62
; 
32'd8933: dataIn1 = 32'd74
; 
32'd8934: dataIn1 = 32'd76
; 
32'd8935: dataIn1 = 32'd82
; 
32'd8936: dataIn1 = 32'd83
; 
32'd8937: dataIn1 = 32'd139
; 
32'd8938: dataIn1 = 32'd141
; 
32'd8939: dataIn1 = 32'd142
; 
32'd8940: dataIn1 = 32'd149
; 
32'd8941: dataIn1 = 32'd196
; 
32'd8942: dataIn1 = 32'd220
; 
32'd8943: dataIn1 = 32'd235
; 
32'd8944: dataIn1 = 32'd242
; 
32'd8945: dataIn1 = 32'd246
; 
32'd8946: dataIn1 = 32'd263
; 
32'd8947: dataIn1 = 32'd288
; 
32'd8948: dataIn1 = 32'd290
; 
32'd8949: dataIn1 = 32'd293
; 
32'd8950: dataIn1 = 32'd294
; 
32'd8951: dataIn1 = 32'd320
; 
32'd8952: dataIn1 = 32'd338
; 
32'd8953: dataIn1 = 32'd370
; 
32'd8954: dataIn1 = 32'd376
; 
32'd8955: dataIn1 = 32'd382
; 
32'd8956: dataIn1 = 32'd397
; 
32'd8957: dataIn1 = 32'd402
; 
32'd8958: dataIn1 = 32'd421
; 
32'd8959: dataIn1 = 32'd424
; 
32'd8960: dataIn1 = 32'd448
; 
32'd8961: dataIn1 = 32'd452
; 
32'd8962: dataIn1 = 32'd472
; 
32'd8963: dataIn1 = 32'd478
; 
32'd8964: dataIn1 = 32'd489
; 
32'd8965: dataIn1 = 32'd494
; 
32'd8966: dataIn1 = 32'd544
; 
32'd8967: dataIn1 = 32'd549
; 
32'd8968: dataIn1 = 32'd560
; 
32'd8969: dataIn1 = 32'd603
; 
32'd8970: dataIn1 = 32'd635
; 
32'd8971: dataIn1 = 32'd683
; 
32'd8972: dataIn1 = 32'd703
; 
32'd8973: dataIn1 = 32'd714
; 
32'd8974: dataIn1 = 32'd728
; 
32'd8975: dataIn1 = 32'd731
; 
32'd8976: dataIn1 = 32'd759
; 
32'd8977: dataIn1 = 32'd776
; 
32'd8978: dataIn1 = 32'd40
; 
32'd8979: dataIn1 = 32'd41
; 
32'd8980: dataIn1 = 32'd45
; 
32'd8981: dataIn1 = 32'd61
; 
32'd8982: dataIn1 = 32'd63
; 
32'd8983: dataIn1 = 32'd98
; 
32'd8984: dataIn1 = 32'd99
; 
32'd8985: dataIn1 = 32'd111
; 
32'd8986: dataIn1 = 32'd116
; 
32'd8987: dataIn1 = 32'd120
; 
32'd8988: dataIn1 = 32'd123
; 
32'd8989: dataIn1 = 32'd136
; 
32'd8990: dataIn1 = 32'd139
; 
32'd8991: dataIn1 = 32'd157
; 
32'd8992: dataIn1 = 32'd161
; 
32'd8993: dataIn1 = 32'd175
; 
32'd8994: dataIn1 = 32'd196
; 
32'd8995: dataIn1 = 32'd202
; 
32'd8996: dataIn1 = 32'd231
; 
32'd8997: dataIn1 = 32'd247
; 
32'd8998: dataIn1 = 32'd303
; 
32'd8999: dataIn1 = 32'd316
; 
32'd9000: dataIn1 = 32'd317
; 
32'd9001: dataIn1 = 32'd327
; 
32'd9002: dataIn1 = 32'd368
; 
32'd9003: dataIn1 = 32'd421
; 
32'd9004: dataIn1 = 32'd444
; 
32'd9005: dataIn1 = 32'd447
; 
32'd9006: dataIn1 = 32'd463
; 
32'd9007: dataIn1 = 32'd464
; 
32'd9008: dataIn1 = 32'd465
; 
32'd9009: dataIn1 = 32'd472
; 
32'd9010: dataIn1 = 32'd485
; 
32'd9011: dataIn1 = 32'd491
; 
32'd9012: dataIn1 = 32'd492
; 
32'd9013: dataIn1 = 32'd524
; 
32'd9014: dataIn1 = 32'd530
; 
32'd9015: dataIn1 = 32'd554
; 
32'd9016: dataIn1 = 32'd571
; 
32'd9017: dataIn1 = 32'd581
; 
32'd9018: dataIn1 = 32'd610
; 
32'd9019: dataIn1 = 32'd611
; 
32'd9020: dataIn1 = 32'd633
; 
32'd9021: dataIn1 = 32'd692
; 
32'd9022: dataIn1 = 32'd747
; 
32'd9023: dataIn1 = 32'd29
; 
32'd9024: dataIn1 = 32'd79
; 
32'd9025: dataIn1 = 32'd111
; 
32'd9026: dataIn1 = 32'd133
; 
32'd9027: dataIn1 = 32'd154
; 
32'd9028: dataIn1 = 32'd179
; 
32'd9029: dataIn1 = 32'd202
; 
32'd9030: dataIn1 = 32'd274
; 
32'd9031: dataIn1 = 32'd286
; 
32'd9032: dataIn1 = 32'd298
; 
32'd9033: dataIn1 = 32'd307
; 
32'd9034: dataIn1 = 32'd337
; 
32'd9035: dataIn1 = 32'd344
; 
32'd9036: dataIn1 = 32'd383
; 
32'd9037: dataIn1 = 32'd387
; 
32'd9038: dataIn1 = 32'd407
; 
32'd9039: dataIn1 = 32'd417
; 
32'd9040: dataIn1 = 32'd427
; 
32'd9041: dataIn1 = 32'd457
; 
32'd9042: dataIn1 = 32'd487
; 
32'd9043: dataIn1 = 32'd489
; 
32'd9044: dataIn1 = 32'd497
; 
32'd9045: dataIn1 = 32'd514
; 
32'd9046: dataIn1 = 32'd525
; 
32'd9047: dataIn1 = 32'd528
; 
32'd9048: dataIn1 = 32'd536
; 
32'd9049: dataIn1 = 32'd567
; 
32'd9050: dataIn1 = 32'd588
; 
32'd9051: dataIn1 = 32'd622
; 
32'd9052: dataIn1 = 32'd630
; 
32'd9053: dataIn1 = 32'd645
; 
32'd9054: dataIn1 = 32'd670
; 
32'd9055: dataIn1 = 32'd682
; 
32'd9056: dataIn1 = 32'd739
; 
32'd9057: dataIn1 = 32'd748
; 
32'd9058: dataIn1 = 32'd776
; 
32'd9059: dataIn1 = 32'd777
; 
32'd9060: dataIn1 = 32'd782
; 
32'd9061: dataIn1 = 32'd795
; 
32'd9062: dataIn1 = 32'd34
; 
32'd9063: dataIn1 = 32'd53
; 
32'd9064: dataIn1 = 32'd93
; 
32'd9065: dataIn1 = 32'd95
; 
32'd9066: dataIn1 = 32'd100
; 
32'd9067: dataIn1 = 32'd116
; 
32'd9068: dataIn1 = 32'd122
; 
32'd9069: dataIn1 = 32'd150
; 
32'd9070: dataIn1 = 32'd171
; 
32'd9071: dataIn1 = 32'd174
; 
32'd9072: dataIn1 = 32'd178
; 
32'd9073: dataIn1 = 32'd192
; 
32'd9074: dataIn1 = 32'd223
; 
32'd9075: dataIn1 = 32'd246
; 
32'd9076: dataIn1 = 32'd249
; 
32'd9077: dataIn1 = 32'd271
; 
32'd9078: dataIn1 = 32'd285
; 
32'd9079: dataIn1 = 32'd295
; 
32'd9080: dataIn1 = 32'd308
; 
32'd9081: dataIn1 = 32'd317
; 
32'd9082: dataIn1 = 32'd348
; 
32'd9083: dataIn1 = 32'd349
; 
32'd9084: dataIn1 = 32'd396
; 
32'd9085: dataIn1 = 32'd400
; 
32'd9086: dataIn1 = 32'd412
; 
32'd9087: dataIn1 = 32'd487
; 
32'd9088: dataIn1 = 32'd490
; 
32'd9089: dataIn1 = 32'd505
; 
32'd9090: dataIn1 = 32'd509
; 
32'd9091: dataIn1 = 32'd537
; 
32'd9092: dataIn1 = 32'd550
; 
32'd9093: dataIn1 = 32'd591
; 
32'd9094: dataIn1 = 32'd615
; 
32'd9095: dataIn1 = 32'd627
; 
32'd9096: dataIn1 = 32'd632
; 
32'd9097: dataIn1 = 32'd676
; 
32'd9098: dataIn1 = 32'd685
; 
32'd9099: dataIn1 = 32'd706
; 
32'd9100: dataIn1 = 32'd729
; 
32'd9101: dataIn1 = 32'd730
; 
32'd9102: dataIn1 = 32'd737
; 
32'd9103: dataIn1 = 32'd754
; 
32'd9104: dataIn1 = 32'd766
; 
32'd9105: dataIn1 = 32'd27
; 
32'd9106: dataIn1 = 32'd35
; 
32'd9107: dataIn1 = 32'd41
; 
32'd9108: dataIn1 = 32'd57
; 
32'd9109: dataIn1 = 32'd98
; 
32'd9110: dataIn1 = 32'd141
; 
32'd9111: dataIn1 = 32'd151
; 
32'd9112: dataIn1 = 32'd152
; 
32'd9113: dataIn1 = 32'd161
; 
32'd9114: dataIn1 = 32'd168
; 
32'd9115: dataIn1 = 32'd185
; 
32'd9116: dataIn1 = 32'd217
; 
32'd9117: dataIn1 = 32'd221
; 
32'd9118: dataIn1 = 32'd247
; 
32'd9119: dataIn1 = 32'd279
; 
32'd9120: dataIn1 = 32'd287
; 
32'd9121: dataIn1 = 32'd298
; 
32'd9122: dataIn1 = 32'd306
; 
32'd9123: dataIn1 = 32'd314
; 
32'd9124: dataIn1 = 32'd338
; 
32'd9125: dataIn1 = 32'd339
; 
32'd9126: dataIn1 = 32'd347
; 
32'd9127: dataIn1 = 32'd379
; 
32'd9128: dataIn1 = 32'd395
; 
32'd9129: dataIn1 = 32'd401
; 
32'd9130: dataIn1 = 32'd402
; 
32'd9131: dataIn1 = 32'd421
; 
32'd9132: dataIn1 = 32'd427
; 
32'd9133: dataIn1 = 32'd428
; 
32'd9134: dataIn1 = 32'd448
; 
32'd9135: dataIn1 = 32'd468
; 
32'd9136: dataIn1 = 32'd475
; 
32'd9137: dataIn1 = 32'd478
; 
32'd9138: dataIn1 = 32'd485
; 
32'd9139: dataIn1 = 32'd508
; 
32'd9140: dataIn1 = 32'd513
; 
32'd9141: dataIn1 = 32'd547
; 
32'd9142: dataIn1 = 32'd571
; 
32'd9143: dataIn1 = 32'd572
; 
32'd9144: dataIn1 = 32'd605
; 
32'd9145: dataIn1 = 32'd615
; 
32'd9146: dataIn1 = 32'd620
; 
32'd9147: dataIn1 = 32'd658
; 
32'd9148: dataIn1 = 32'd670
; 
32'd9149: dataIn1 = 32'd689
; 
32'd9150: dataIn1 = 32'd710
; 
32'd9151: dataIn1 = 32'd728
; 
32'd9152: dataIn1 = 32'd739
; 
32'd9153: dataIn1 = 32'd755
; 
32'd9154: dataIn1 = 32'd758
; 
32'd9155: dataIn1 = 32'd779
; 
32'd9156: dataIn1 = 32'd796
; 
32'd9157: dataIn1 = 32'd47
; 
32'd9158: dataIn1 = 32'd65
; 
32'd9159: dataIn1 = 32'd73
; 
32'd9160: dataIn1 = 32'd105
; 
32'd9161: dataIn1 = 32'd111
; 
32'd9162: dataIn1 = 32'd112
; 
32'd9163: dataIn1 = 32'd114
; 
32'd9164: dataIn1 = 32'd150
; 
32'd9165: dataIn1 = 32'd169
; 
32'd9166: dataIn1 = 32'd202
; 
32'd9167: dataIn1 = 32'd217
; 
32'd9168: dataIn1 = 32'd234
; 
32'd9169: dataIn1 = 32'd242
; 
32'd9170: dataIn1 = 32'd249
; 
32'd9171: dataIn1 = 32'd251
; 
32'd9172: dataIn1 = 32'd252
; 
32'd9173: dataIn1 = 32'd334
; 
32'd9174: dataIn1 = 32'd342
; 
32'd9175: dataIn1 = 32'd347
; 
32'd9176: dataIn1 = 32'd363
; 
32'd9177: dataIn1 = 32'd377
; 
32'd9178: dataIn1 = 32'd385
; 
32'd9179: dataIn1 = 32'd394
; 
32'd9180: dataIn1 = 32'd408
; 
32'd9181: dataIn1 = 32'd437
; 
32'd9182: dataIn1 = 32'd447
; 
32'd9183: dataIn1 = 32'd448
; 
32'd9184: dataIn1 = 32'd483
; 
32'd9185: dataIn1 = 32'd485
; 
32'd9186: dataIn1 = 32'd503
; 
32'd9187: dataIn1 = 32'd508
; 
32'd9188: dataIn1 = 32'd516
; 
32'd9189: dataIn1 = 32'd560
; 
32'd9190: dataIn1 = 32'd562
; 
32'd9191: dataIn1 = 32'd617
; 
32'd9192: dataIn1 = 32'd621
; 
32'd9193: dataIn1 = 32'd670
; 
32'd9194: dataIn1 = 32'd686
; 
32'd9195: dataIn1 = 32'd692
; 
32'd9196: dataIn1 = 32'd695
; 
32'd9197: dataIn1 = 32'd723
; 
32'd9198: dataIn1 = 32'd726
; 
32'd9199: dataIn1 = 32'd732
; 
32'd9200: dataIn1 = 32'd751
; 
32'd9201: dataIn1 = 32'd759
; 
32'd9202: dataIn1 = 32'd762
; 
32'd9203: dataIn1 = 32'd62
; 
32'd9204: dataIn1 = 32'd66
; 
32'd9205: dataIn1 = 32'd104
; 
32'd9206: dataIn1 = 32'd129
; 
32'd9207: dataIn1 = 32'd131
; 
32'd9208: dataIn1 = 32'd134
; 
32'd9209: dataIn1 = 32'd143
; 
32'd9210: dataIn1 = 32'd176
; 
32'd9211: dataIn1 = 32'd191
; 
32'd9212: dataIn1 = 32'd206
; 
32'd9213: dataIn1 = 32'd220
; 
32'd9214: dataIn1 = 32'd229
; 
32'd9215: dataIn1 = 32'd324
; 
32'd9216: dataIn1 = 32'd358
; 
32'd9217: dataIn1 = 32'd363
; 
32'd9218: dataIn1 = 32'd397
; 
32'd9219: dataIn1 = 32'd398
; 
32'd9220: dataIn1 = 32'd408
; 
32'd9221: dataIn1 = 32'd412
; 
32'd9222: dataIn1 = 32'd422
; 
32'd9223: dataIn1 = 32'd443
; 
32'd9224: dataIn1 = 32'd452
; 
32'd9225: dataIn1 = 32'd458
; 
32'd9226: dataIn1 = 32'd467
; 
32'd9227: dataIn1 = 32'd481
; 
32'd9228: dataIn1 = 32'd499
; 
32'd9229: dataIn1 = 32'd506
; 
32'd9230: dataIn1 = 32'd528
; 
32'd9231: dataIn1 = 32'd532
; 
32'd9232: dataIn1 = 32'd547
; 
32'd9233: dataIn1 = 32'd571
; 
32'd9234: dataIn1 = 32'd583
; 
32'd9235: dataIn1 = 32'd603
; 
32'd9236: dataIn1 = 32'd605
; 
32'd9237: dataIn1 = 32'd607
; 
32'd9238: dataIn1 = 32'd624
; 
32'd9239: dataIn1 = 32'd626
; 
32'd9240: dataIn1 = 32'd646
; 
32'd9241: dataIn1 = 32'd647
; 
32'd9242: dataIn1 = 32'd675
; 
32'd9243: dataIn1 = 32'd677
; 
32'd9244: dataIn1 = 32'd684
; 
32'd9245: dataIn1 = 32'd685
; 
32'd9246: dataIn1 = 32'd723
; 
32'd9247: dataIn1 = 32'd731
; 
32'd9248: dataIn1 = 32'd760
; 
32'd9249: dataIn1 = 32'd772
; 
32'd9250: dataIn1 = 32'd786
; 
32'd9251: dataIn1 = 32'd792
; 
32'd9252: dataIn1 = 32'd34
; 
32'd9253: dataIn1 = 32'd35
; 
32'd9254: dataIn1 = 32'd36
; 
32'd9255: dataIn1 = 32'd41
; 
32'd9256: dataIn1 = 32'd58
; 
32'd9257: dataIn1 = 32'd60
; 
32'd9258: dataIn1 = 32'd92
; 
32'd9259: dataIn1 = 32'd105
; 
32'd9260: dataIn1 = 32'd135
; 
32'd9261: dataIn1 = 32'd152
; 
32'd9262: dataIn1 = 32'd153
; 
32'd9263: dataIn1 = 32'd159
; 
32'd9264: dataIn1 = 32'd160
; 
32'd9265: dataIn1 = 32'd177
; 
32'd9266: dataIn1 = 32'd204
; 
32'd9267: dataIn1 = 32'd210
; 
32'd9268: dataIn1 = 32'd246
; 
32'd9269: dataIn1 = 32'd284
; 
32'd9270: dataIn1 = 32'd300
; 
32'd9271: dataIn1 = 32'd372
; 
32'd9272: dataIn1 = 32'd379
; 
32'd9273: dataIn1 = 32'd393
; 
32'd9274: dataIn1 = 32'd435
; 
32'd9275: dataIn1 = 32'd437
; 
32'd9276: dataIn1 = 32'd470
; 
32'd9277: dataIn1 = 32'd485
; 
32'd9278: dataIn1 = 32'd501
; 
32'd9279: dataIn1 = 32'd506
; 
32'd9280: dataIn1 = 32'd513
; 
32'd9281: dataIn1 = 32'd531
; 
32'd9282: dataIn1 = 32'd532
; 
32'd9283: dataIn1 = 32'd539
; 
32'd9284: dataIn1 = 32'd541
; 
32'd9285: dataIn1 = 32'd563
; 
32'd9286: dataIn1 = 32'd587
; 
32'd9287: dataIn1 = 32'd614
; 
32'd9288: dataIn1 = 32'd616
; 
32'd9289: dataIn1 = 32'd688
; 
32'd9290: dataIn1 = 32'd718
; 
32'd9291: dataIn1 = 32'd735
; 
32'd9292: dataIn1 = 32'd737
; 
32'd9293: dataIn1 = 32'd758
; 
32'd9294: dataIn1 = 32'd771
; 
32'd9295: dataIn1 = 32'd48
; 
32'd9296: dataIn1 = 32'd52
; 
32'd9297: dataIn1 = 32'd58
; 
32'd9298: dataIn1 = 32'd65
; 
32'd9299: dataIn1 = 32'd67
; 
32'd9300: dataIn1 = 32'd78
; 
32'd9301: dataIn1 = 32'd112
; 
32'd9302: dataIn1 = 32'd119
; 
32'd9303: dataIn1 = 32'd142
; 
32'd9304: dataIn1 = 32'd200
; 
32'd9305: dataIn1 = 32'd217
; 
32'd9306: dataIn1 = 32'd237
; 
32'd9307: dataIn1 = 32'd249
; 
32'd9308: dataIn1 = 32'd273
; 
32'd9309: dataIn1 = 32'd288
; 
32'd9310: dataIn1 = 32'd309
; 
32'd9311: dataIn1 = 32'd313
; 
32'd9312: dataIn1 = 32'd322
; 
32'd9313: dataIn1 = 32'd325
; 
32'd9314: dataIn1 = 32'd332
; 
32'd9315: dataIn1 = 32'd351
; 
32'd9316: dataIn1 = 32'd355
; 
32'd9317: dataIn1 = 32'd359
; 
32'd9318: dataIn1 = 32'd382
; 
32'd9319: dataIn1 = 32'd390
; 
32'd9320: dataIn1 = 32'd397
; 
32'd9321: dataIn1 = 32'd418
; 
32'd9322: dataIn1 = 32'd422
; 
32'd9323: dataIn1 = 32'd437
; 
32'd9324: dataIn1 = 32'd455
; 
32'd9325: dataIn1 = 32'd459
; 
32'd9326: dataIn1 = 32'd467
; 
32'd9327: dataIn1 = 32'd474
; 
32'd9328: dataIn1 = 32'd486
; 
32'd9329: dataIn1 = 32'd508
; 
32'd9330: dataIn1 = 32'd561
; 
32'd9331: dataIn1 = 32'd575
; 
32'd9332: dataIn1 = 32'd582
; 
32'd9333: dataIn1 = 32'd617
; 
32'd9334: dataIn1 = 32'd619
; 
32'd9335: dataIn1 = 32'd629
; 
32'd9336: dataIn1 = 32'd640
; 
32'd9337: dataIn1 = 32'd644
; 
32'd9338: dataIn1 = 32'd661
; 
32'd9339: dataIn1 = 32'd684
; 
32'd9340: dataIn1 = 32'd698
; 
32'd9341: dataIn1 = 32'd732
; 
32'd9342: dataIn1 = 32'd739
; 
32'd9343: dataIn1 = 32'd788
; 
32'd9344: dataIn1 = 32'd43
; 
32'd9345: dataIn1 = 32'd53
; 
32'd9346: dataIn1 = 32'd54
; 
32'd9347: dataIn1 = 32'd83
; 
32'd9348: dataIn1 = 32'd101
; 
32'd9349: dataIn1 = 32'd146
; 
32'd9350: dataIn1 = 32'd147
; 
32'd9351: dataIn1 = 32'd148
; 
32'd9352: dataIn1 = 32'd152
; 
32'd9353: dataIn1 = 32'd177
; 
32'd9354: dataIn1 = 32'd205
; 
32'd9355: dataIn1 = 32'd212
; 
32'd9356: dataIn1 = 32'd225
; 
32'd9357: dataIn1 = 32'd231
; 
32'd9358: dataIn1 = 32'd234
; 
32'd9359: dataIn1 = 32'd251
; 
32'd9360: dataIn1 = 32'd252
; 
32'd9361: dataIn1 = 32'd255
; 
32'd9362: dataIn1 = 32'd260
; 
32'd9363: dataIn1 = 32'd267
; 
32'd9364: dataIn1 = 32'd288
; 
32'd9365: dataIn1 = 32'd301
; 
32'd9366: dataIn1 = 32'd320
; 
32'd9367: dataIn1 = 32'd323
; 
32'd9368: dataIn1 = 32'd343
; 
32'd9369: dataIn1 = 32'd348
; 
32'd9370: dataIn1 = 32'd362
; 
32'd9371: dataIn1 = 32'd386
; 
32'd9372: dataIn1 = 32'd410
; 
32'd9373: dataIn1 = 32'd415
; 
32'd9374: dataIn1 = 32'd421
; 
32'd9375: dataIn1 = 32'd451
; 
32'd9376: dataIn1 = 32'd484
; 
32'd9377: dataIn1 = 32'd519
; 
32'd9378: dataIn1 = 32'd535
; 
32'd9379: dataIn1 = 32'd570
; 
32'd9380: dataIn1 = 32'd581
; 
32'd9381: dataIn1 = 32'd587
; 
32'd9382: dataIn1 = 32'd589
; 
32'd9383: dataIn1 = 32'd627
; 
32'd9384: dataIn1 = 32'd633
; 
32'd9385: dataIn1 = 32'd680
; 
32'd9386: dataIn1 = 32'd731
; 
32'd9387: dataIn1 = 32'd743
; 
32'd9388: dataIn1 = 32'd755
; 
32'd9389: dataIn1 = 32'd762
; 
32'd9390: dataIn1 = 32'd763
; 
32'd9391: dataIn1 = 32'd765
; 
32'd9392: dataIn1 = 32'd35
; 
32'd9393: dataIn1 = 32'd41
; 
32'd9394: dataIn1 = 32'd84
; 
32'd9395: dataIn1 = 32'd87
; 
32'd9396: dataIn1 = 32'd102
; 
32'd9397: dataIn1 = 32'd112
; 
32'd9398: dataIn1 = 32'd117
; 
32'd9399: dataIn1 = 32'd141
; 
32'd9400: dataIn1 = 32'd146
; 
32'd9401: dataIn1 = 32'd158
; 
32'd9402: dataIn1 = 32'd163
; 
32'd9403: dataIn1 = 32'd175
; 
32'd9404: dataIn1 = 32'd179
; 
32'd9405: dataIn1 = 32'd200
; 
32'd9406: dataIn1 = 32'd203
; 
32'd9407: dataIn1 = 32'd210
; 
32'd9408: dataIn1 = 32'd213
; 
32'd9409: dataIn1 = 32'd255
; 
32'd9410: dataIn1 = 32'd268
; 
32'd9411: dataIn1 = 32'd269
; 
32'd9412: dataIn1 = 32'd308
; 
32'd9413: dataIn1 = 32'd319
; 
32'd9414: dataIn1 = 32'd332
; 
32'd9415: dataIn1 = 32'd340
; 
32'd9416: dataIn1 = 32'd353
; 
32'd9417: dataIn1 = 32'd366
; 
32'd9418: dataIn1 = 32'd384
; 
32'd9419: dataIn1 = 32'd397
; 
32'd9420: dataIn1 = 32'd414
; 
32'd9421: dataIn1 = 32'd427
; 
32'd9422: dataIn1 = 32'd453
; 
32'd9423: dataIn1 = 32'd470
; 
32'd9424: dataIn1 = 32'd531
; 
32'd9425: dataIn1 = 32'd539
; 
32'd9426: dataIn1 = 32'd572
; 
32'd9427: dataIn1 = 32'd603
; 
32'd9428: dataIn1 = 32'd606
; 
32'd9429: dataIn1 = 32'd655
; 
32'd9430: dataIn1 = 32'd659
; 
32'd9431: dataIn1 = 32'd666
; 
32'd9432: dataIn1 = 32'd697
; 
32'd9433: dataIn1 = 32'd699
; 
32'd9434: dataIn1 = 32'd714
; 
32'd9435: dataIn1 = 32'd719
; 
32'd9436: dataIn1 = 32'd740
; 
32'd9437: dataIn1 = 32'd759
; 
32'd9438: dataIn1 = 32'd794
; 
32'd9439: dataIn1 = 32'd34
; 
32'd9440: dataIn1 = 32'd87
; 
32'd9441: dataIn1 = 32'd136
; 
32'd9442: dataIn1 = 32'd149
; 
32'd9443: dataIn1 = 32'd234
; 
32'd9444: dataIn1 = 32'd255
; 
32'd9445: dataIn1 = 32'd263
; 
32'd9446: dataIn1 = 32'd269
; 
32'd9447: dataIn1 = 32'd288
; 
32'd9448: dataIn1 = 32'd289
; 
32'd9449: dataIn1 = 32'd343
; 
32'd9450: dataIn1 = 32'd356
; 
32'd9451: dataIn1 = 32'd370
; 
32'd9452: dataIn1 = 32'd411
; 
32'd9453: dataIn1 = 32'd423
; 
32'd9454: dataIn1 = 32'd426
; 
32'd9455: dataIn1 = 32'd435
; 
32'd9456: dataIn1 = 32'd493
; 
32'd9457: dataIn1 = 32'd507
; 
32'd9458: dataIn1 = 32'd515
; 
32'd9459: dataIn1 = 32'd519
; 
32'd9460: dataIn1 = 32'd520
; 
32'd9461: dataIn1 = 32'd535
; 
32'd9462: dataIn1 = 32'd537
; 
32'd9463: dataIn1 = 32'd558
; 
32'd9464: dataIn1 = 32'd576
; 
32'd9465: dataIn1 = 32'd600
; 
32'd9466: dataIn1 = 32'd616
; 
32'd9467: dataIn1 = 32'd622
; 
32'd9468: dataIn1 = 32'd630
; 
32'd9469: dataIn1 = 32'd650
; 
32'd9470: dataIn1 = 32'd674
; 
32'd9471: dataIn1 = 32'd684
; 
32'd9472: dataIn1 = 32'd688
; 
32'd9473: dataIn1 = 32'd704
; 
32'd9474: dataIn1 = 32'd713
; 
32'd9475: dataIn1 = 32'd722
; 
32'd9476: dataIn1 = 32'd732
; 
32'd9477: dataIn1 = 32'd762
; 
32'd9478: dataIn1 = 32'd773
; 
32'd9479: dataIn1 = 32'd783
; 
32'd9480: dataIn1 = 32'd793
; 
32'd9481: dataIn1 = 32'd798
; 
32'd9482: dataIn1 = 32'd44
; 
32'd9483: dataIn1 = 32'd54
; 
32'd9484: dataIn1 = 32'd61
; 
32'd9485: dataIn1 = 32'd76
; 
32'd9486: dataIn1 = 32'd98
; 
32'd9487: dataIn1 = 32'd121
; 
32'd9488: dataIn1 = 32'd123
; 
32'd9489: dataIn1 = 32'd130
; 
32'd9490: dataIn1 = 32'd132
; 
32'd9491: dataIn1 = 32'd151
; 
32'd9492: dataIn1 = 32'd162
; 
32'd9493: dataIn1 = 32'd175
; 
32'd9494: dataIn1 = 32'd189
; 
32'd9495: dataIn1 = 32'd211
; 
32'd9496: dataIn1 = 32'd219
; 
32'd9497: dataIn1 = 32'd221
; 
32'd9498: dataIn1 = 32'd247
; 
32'd9499: dataIn1 = 32'd248
; 
32'd9500: dataIn1 = 32'd269
; 
32'd9501: dataIn1 = 32'd281
; 
32'd9502: dataIn1 = 32'd345
; 
32'd9503: dataIn1 = 32'd349
; 
32'd9504: dataIn1 = 32'd360
; 
32'd9505: dataIn1 = 32'd368
; 
32'd9506: dataIn1 = 32'd383
; 
32'd9507: dataIn1 = 32'd403
; 
32'd9508: dataIn1 = 32'd413
; 
32'd9509: dataIn1 = 32'd448
; 
32'd9510: dataIn1 = 32'd456
; 
32'd9511: dataIn1 = 32'd483
; 
32'd9512: dataIn1 = 32'd493
; 
32'd9513: dataIn1 = 32'd567
; 
32'd9514: dataIn1 = 32'd590
; 
32'd9515: dataIn1 = 32'd599
; 
32'd9516: dataIn1 = 32'd613
; 
32'd9517: dataIn1 = 32'd632
; 
32'd9518: dataIn1 = 32'd645
; 
32'd9519: dataIn1 = 32'd688
; 
32'd9520: dataIn1 = 32'd702
; 
32'd9521: dataIn1 = 32'd775
; 
32'd9522: dataIn1 = 32'd50
; 
32'd9523: dataIn1 = 32'd69
; 
32'd9524: dataIn1 = 32'd82
; 
32'd9525: dataIn1 = 32'd93
; 
32'd9526: dataIn1 = 32'd96
; 
32'd9527: dataIn1 = 32'd133
; 
32'd9528: dataIn1 = 32'd143
; 
32'd9529: dataIn1 = 32'd162
; 
32'd9530: dataIn1 = 32'd178
; 
32'd9531: dataIn1 = 32'd181
; 
32'd9532: dataIn1 = 32'd197
; 
32'd9533: dataIn1 = 32'd200
; 
32'd9534: dataIn1 = 32'd210
; 
32'd9535: dataIn1 = 32'd221
; 
32'd9536: dataIn1 = 32'd264
; 
32'd9537: dataIn1 = 32'd276
; 
32'd9538: dataIn1 = 32'd293
; 
32'd9539: dataIn1 = 32'd340
; 
32'd9540: dataIn1 = 32'd373
; 
32'd9541: dataIn1 = 32'd383
; 
32'd9542: dataIn1 = 32'd402
; 
32'd9543: dataIn1 = 32'd483
; 
32'd9544: dataIn1 = 32'd504
; 
32'd9545: dataIn1 = 32'd505
; 
32'd9546: dataIn1 = 32'd518
; 
32'd9547: dataIn1 = 32'd554
; 
32'd9548: dataIn1 = 32'd565
; 
32'd9549: dataIn1 = 32'd568
; 
32'd9550: dataIn1 = 32'd569
; 
32'd9551: dataIn1 = 32'd571
; 
32'd9552: dataIn1 = 32'd572
; 
32'd9553: dataIn1 = 32'd584
; 
32'd9554: dataIn1 = 32'd588
; 
32'd9555: dataIn1 = 32'd593
; 
32'd9556: dataIn1 = 32'd600
; 
32'd9557: dataIn1 = 32'd665
; 
32'd9558: dataIn1 = 32'd684
; 
32'd9559: dataIn1 = 32'd699
; 
32'd9560: dataIn1 = 32'd762
; 
32'd9561: dataIn1 = 32'd769
; 
32'd9562: dataIn1 = 32'd772
; 
32'd9563: dataIn1 = 32'd774
; 
32'd9564: dataIn1 = 32'd775
; 
32'd9565: dataIn1 = 32'd789
; 
32'd9566: dataIn1 = 32'd39
; 
32'd9567: dataIn1 = 32'd76
; 
32'd9568: dataIn1 = 32'd98
; 
32'd9569: dataIn1 = 32'd116
; 
32'd9570: dataIn1 = 32'd120
; 
32'd9571: dataIn1 = 32'd134
; 
32'd9572: dataIn1 = 32'd171
; 
32'd9573: dataIn1 = 32'd175
; 
32'd9574: dataIn1 = 32'd184
; 
32'd9575: dataIn1 = 32'd185
; 
32'd9576: dataIn1 = 32'd204
; 
32'd9577: dataIn1 = 32'd216
; 
32'd9578: dataIn1 = 32'd221
; 
32'd9579: dataIn1 = 32'd224
; 
32'd9580: dataIn1 = 32'd225
; 
32'd9581: dataIn1 = 32'd237
; 
32'd9582: dataIn1 = 32'd239
; 
32'd9583: dataIn1 = 32'd252
; 
32'd9584: dataIn1 = 32'd259
; 
32'd9585: dataIn1 = 32'd268
; 
32'd9586: dataIn1 = 32'd295
; 
32'd9587: dataIn1 = 32'd297
; 
32'd9588: dataIn1 = 32'd333
; 
32'd9589: dataIn1 = 32'd359
; 
32'd9590: dataIn1 = 32'd377
; 
32'd9591: dataIn1 = 32'd388
; 
32'd9592: dataIn1 = 32'd407
; 
32'd9593: dataIn1 = 32'd414
; 
32'd9594: dataIn1 = 32'd419
; 
32'd9595: dataIn1 = 32'd433
; 
32'd9596: dataIn1 = 32'd442
; 
32'd9597: dataIn1 = 32'd445
; 
32'd9598: dataIn1 = 32'd453
; 
32'd9599: dataIn1 = 32'd465
; 
32'd9600: dataIn1 = 32'd470
; 
32'd9601: dataIn1 = 32'd484
; 
32'd9602: dataIn1 = 32'd489
; 
32'd9603: dataIn1 = 32'd507
; 
32'd9604: dataIn1 = 32'd513
; 
32'd9605: dataIn1 = 32'd539
; 
32'd9606: dataIn1 = 32'd547
; 
32'd9607: dataIn1 = 32'd550
; 
32'd9608: dataIn1 = 32'd559
; 
32'd9609: dataIn1 = 32'd561
; 
32'd9610: dataIn1 = 32'd583
; 
32'd9611: dataIn1 = 32'd585
; 
32'd9612: dataIn1 = 32'd598
; 
32'd9613: dataIn1 = 32'd611
; 
32'd9614: dataIn1 = 32'd620
; 
32'd9615: dataIn1 = 32'd623
; 
32'd9616: dataIn1 = 32'd624
; 
32'd9617: dataIn1 = 32'd631
; 
32'd9618: dataIn1 = 32'd660
; 
32'd9619: dataIn1 = 32'd666
; 
32'd9620: dataIn1 = 32'd688
; 
32'd9621: dataIn1 = 32'd699
; 
32'd9622: dataIn1 = 32'd738
; 
32'd9623: dataIn1 = 32'd762
; 
32'd9624: dataIn1 = 32'd799
; 
32'd9625: dataIn1 = 32'd50
; 
32'd9626: dataIn1 = 32'd64
; 
32'd9627: dataIn1 = 32'd96
; 
32'd9628: dataIn1 = 32'd113
; 
32'd9629: dataIn1 = 32'd123
; 
32'd9630: dataIn1 = 32'd132
; 
32'd9631: dataIn1 = 32'd150
; 
32'd9632: dataIn1 = 32'd192
; 
32'd9633: dataIn1 = 32'd197
; 
32'd9634: dataIn1 = 32'd212
; 
32'd9635: dataIn1 = 32'd223
; 
32'd9636: dataIn1 = 32'd256
; 
32'd9637: dataIn1 = 32'd260
; 
32'd9638: dataIn1 = 32'd294
; 
32'd9639: dataIn1 = 32'd304
; 
32'd9640: dataIn1 = 32'd321
; 
32'd9641: dataIn1 = 32'd323
; 
32'd9642: dataIn1 = 32'd332
; 
32'd9643: dataIn1 = 32'd335
; 
32'd9644: dataIn1 = 32'd340
; 
32'd9645: dataIn1 = 32'd416
; 
32'd9646: dataIn1 = 32'd423
; 
32'd9647: dataIn1 = 32'd428
; 
32'd9648: dataIn1 = 32'd481
; 
32'd9649: dataIn1 = 32'd484
; 
32'd9650: dataIn1 = 32'd497
; 
32'd9651: dataIn1 = 32'd596
; 
32'd9652: dataIn1 = 32'd666
; 
32'd9653: dataIn1 = 32'd670
; 
32'd9654: dataIn1 = 32'd738
; 
32'd9655: dataIn1 = 32'd739
; 
32'd9656: dataIn1 = 32'd741
; 
32'd9657: dataIn1 = 32'd748
; 
32'd9658: dataIn1 = 32'd754
; 
32'd9659: dataIn1 = 32'd755
; 
32'd9660: dataIn1 = 32'd758
; 
32'd9661: dataIn1 = 32'd778
; 
32'd9662: dataIn1 = 32'd781
; 
32'd9663: dataIn1 = 32'd39
; 
32'd9664: dataIn1 = 32'd79
; 
32'd9665: dataIn1 = 32'd132
; 
32'd9666: dataIn1 = 32'd137
; 
32'd9667: dataIn1 = 32'd156
; 
32'd9668: dataIn1 = 32'd162
; 
32'd9669: dataIn1 = 32'd179
; 
32'd9670: dataIn1 = 32'd264
; 
32'd9671: dataIn1 = 32'd286
; 
32'd9672: dataIn1 = 32'd318
; 
32'd9673: dataIn1 = 32'd350
; 
32'd9674: dataIn1 = 32'd355
; 
32'd9675: dataIn1 = 32'd382
; 
32'd9676: dataIn1 = 32'd384
; 
32'd9677: dataIn1 = 32'd397
; 
32'd9678: dataIn1 = 32'd416
; 
32'd9679: dataIn1 = 32'd453
; 
32'd9680: dataIn1 = 32'd470
; 
32'd9681: dataIn1 = 32'd481
; 
32'd9682: dataIn1 = 32'd505
; 
32'd9683: dataIn1 = 32'd511
; 
32'd9684: dataIn1 = 32'd513
; 
32'd9685: dataIn1 = 32'd515
; 
32'd9686: dataIn1 = 32'd520
; 
32'd9687: dataIn1 = 32'd521
; 
32'd9688: dataIn1 = 32'd523
; 
32'd9689: dataIn1 = 32'd533
; 
32'd9690: dataIn1 = 32'd601
; 
32'd9691: dataIn1 = 32'd621
; 
32'd9692: dataIn1 = 32'd623
; 
32'd9693: dataIn1 = 32'd647
; 
32'd9694: dataIn1 = 32'd674
; 
32'd9695: dataIn1 = 32'd682
; 
32'd9696: dataIn1 = 32'd685
; 
32'd9697: dataIn1 = 32'd689
; 
32'd9698: dataIn1 = 32'd712
; 
32'd9699: dataIn1 = 32'd748
; 
32'd9700: dataIn1 = 32'd752
; 
32'd9701: dataIn1 = 32'd765
; 
32'd9702: dataIn1 = 32'd97
; 
32'd9703: dataIn1 = 32'd190
; 
32'd9704: dataIn1 = 32'd192
; 
32'd9705: dataIn1 = 32'd202
; 
32'd9706: dataIn1 = 32'd203
; 
32'd9707: dataIn1 = 32'd272
; 
32'd9708: dataIn1 = 32'd274
; 
32'd9709: dataIn1 = 32'd283
; 
32'd9710: dataIn1 = 32'd285
; 
32'd9711: dataIn1 = 32'd289
; 
32'd9712: dataIn1 = 32'd315
; 
32'd9713: dataIn1 = 32'd329
; 
32'd9714: dataIn1 = 32'd333
; 
32'd9715: dataIn1 = 32'd356
; 
32'd9716: dataIn1 = 32'd365
; 
32'd9717: dataIn1 = 32'd375
; 
32'd9718: dataIn1 = 32'd396
; 
32'd9719: dataIn1 = 32'd411
; 
32'd9720: dataIn1 = 32'd419
; 
32'd9721: dataIn1 = 32'd428
; 
32'd9722: dataIn1 = 32'd434
; 
32'd9723: dataIn1 = 32'd448
; 
32'd9724: dataIn1 = 32'd450
; 
32'd9725: dataIn1 = 32'd485
; 
32'd9726: dataIn1 = 32'd505
; 
32'd9727: dataIn1 = 32'd526
; 
32'd9728: dataIn1 = 32'd547
; 
32'd9729: dataIn1 = 32'd598
; 
32'd9730: dataIn1 = 32'd644
; 
32'd9731: dataIn1 = 32'd645
; 
32'd9732: dataIn1 = 32'd668
; 
32'd9733: dataIn1 = 32'd697
; 
32'd9734: dataIn1 = 32'd711
; 
32'd9735: dataIn1 = 32'd758
; 
32'd9736: dataIn1 = 32'd779
; 
32'd9737: dataIn1 = 32'd60
; 
32'd9738: dataIn1 = 32'd91
; 
32'd9739: dataIn1 = 32'd111
; 
32'd9740: dataIn1 = 32'd182
; 
32'd9741: dataIn1 = 32'd188
; 
32'd9742: dataIn1 = 32'd203
; 
32'd9743: dataIn1 = 32'd223
; 
32'd9744: dataIn1 = 32'd225
; 
32'd9745: dataIn1 = 32'd231
; 
32'd9746: dataIn1 = 32'd235
; 
32'd9747: dataIn1 = 32'd241
; 
32'd9748: dataIn1 = 32'd278
; 
32'd9749: dataIn1 = 32'd283
; 
32'd9750: dataIn1 = 32'd288
; 
32'd9751: dataIn1 = 32'd303
; 
32'd9752: dataIn1 = 32'd370
; 
32'd9753: dataIn1 = 32'd372
; 
32'd9754: dataIn1 = 32'd377
; 
32'd9755: dataIn1 = 32'd381
; 
32'd9756: dataIn1 = 32'd393
; 
32'd9757: dataIn1 = 32'd395
; 
32'd9758: dataIn1 = 32'd420
; 
32'd9759: dataIn1 = 32'd446
; 
32'd9760: dataIn1 = 32'd451
; 
32'd9761: dataIn1 = 32'd453
; 
32'd9762: dataIn1 = 32'd459
; 
32'd9763: dataIn1 = 32'd463
; 
32'd9764: dataIn1 = 32'd500
; 
32'd9765: dataIn1 = 32'd514
; 
32'd9766: dataIn1 = 32'd525
; 
32'd9767: dataIn1 = 32'd538
; 
32'd9768: dataIn1 = 32'd552
; 
32'd9769: dataIn1 = 32'd554
; 
32'd9770: dataIn1 = 32'd606
; 
32'd9771: dataIn1 = 32'd640
; 
32'd9772: dataIn1 = 32'd644
; 
32'd9773: dataIn1 = 32'd685
; 
32'd9774: dataIn1 = 32'd695
; 
32'd9775: dataIn1 = 32'd708
; 
32'd9776: dataIn1 = 32'd712
; 
32'd9777: dataIn1 = 32'd722
; 
32'd9778: dataIn1 = 32'd728
; 
32'd9779: dataIn1 = 32'd751
; 
32'd9780: dataIn1 = 32'd772
; 
32'd9781: dataIn1 = 32'd778
; 
32'd9782: dataIn1 = 32'd797
; 
32'd9783: dataIn1 = 32'd798
; 
32'd9784: dataIn1 = 32'd800
; 
32'd9785: dataIn1 = 32'd68
; 
32'd9786: dataIn1 = 32'd71
; 
32'd9787: dataIn1 = 32'd76
; 
32'd9788: dataIn1 = 32'd87
; 
32'd9789: dataIn1 = 32'd100
; 
32'd9790: dataIn1 = 32'd119
; 
32'd9791: dataIn1 = 32'd121
; 
32'd9792: dataIn1 = 32'd124
; 
32'd9793: dataIn1 = 32'd132
; 
32'd9794: dataIn1 = 32'd144
; 
32'd9795: dataIn1 = 32'd185
; 
32'd9796: dataIn1 = 32'd239
; 
32'd9797: dataIn1 = 32'd247
; 
32'd9798: dataIn1 = 32'd253
; 
32'd9799: dataIn1 = 32'd287
; 
32'd9800: dataIn1 = 32'd313
; 
32'd9801: dataIn1 = 32'd332
; 
32'd9802: dataIn1 = 32'd338
; 
32'd9803: dataIn1 = 32'd356
; 
32'd9804: dataIn1 = 32'd362
; 
32'd9805: dataIn1 = 32'd384
; 
32'd9806: dataIn1 = 32'd386
; 
32'd9807: dataIn1 = 32'd390
; 
32'd9808: dataIn1 = 32'd423
; 
32'd9809: dataIn1 = 32'd450
; 
32'd9810: dataIn1 = 32'd451
; 
32'd9811: dataIn1 = 32'd461
; 
32'd9812: dataIn1 = 32'd489
; 
32'd9813: dataIn1 = 32'd495
; 
32'd9814: dataIn1 = 32'd496
; 
32'd9815: dataIn1 = 32'd520
; 
32'd9816: dataIn1 = 32'd533
; 
32'd9817: dataIn1 = 32'd546
; 
32'd9818: dataIn1 = 32'd547
; 
32'd9819: dataIn1 = 32'd555
; 
32'd9820: dataIn1 = 32'd588
; 
32'd9821: dataIn1 = 32'd591
; 
32'd9822: dataIn1 = 32'd639
; 
32'd9823: dataIn1 = 32'd651
; 
32'd9824: dataIn1 = 32'd655
; 
32'd9825: dataIn1 = 32'd687
; 
32'd9826: dataIn1 = 32'd696
; 
32'd9827: dataIn1 = 32'd697
; 
32'd9828: dataIn1 = 32'd768
; 
32'd9829: dataIn1 = 32'd779
; 
32'd9830: dataIn1 = 32'd787
; 
32'd9831: dataIn1 = 32'd794
; 
32'd9832: dataIn1 = 32'd68
; 
32'd9833: dataIn1 = 32'd73
; 
32'd9834: dataIn1 = 32'd77
; 
32'd9835: dataIn1 = 32'd84
; 
32'd9836: dataIn1 = 32'd94
; 
32'd9837: dataIn1 = 32'd138
; 
32'd9838: dataIn1 = 32'd154
; 
32'd9839: dataIn1 = 32'd163
; 
32'd9840: dataIn1 = 32'd186
; 
32'd9841: dataIn1 = 32'd210
; 
32'd9842: dataIn1 = 32'd211
; 
32'd9843: dataIn1 = 32'd223
; 
32'd9844: dataIn1 = 32'd243
; 
32'd9845: dataIn1 = 32'd253
; 
32'd9846: dataIn1 = 32'd268
; 
32'd9847: dataIn1 = 32'd271
; 
32'd9848: dataIn1 = 32'd306
; 
32'd9849: dataIn1 = 32'd332
; 
32'd9850: dataIn1 = 32'd342
; 
32'd9851: dataIn1 = 32'd350
; 
32'd9852: dataIn1 = 32'd355
; 
32'd9853: dataIn1 = 32'd374
; 
32'd9854: dataIn1 = 32'd392
; 
32'd9855: dataIn1 = 32'd402
; 
32'd9856: dataIn1 = 32'd423
; 
32'd9857: dataIn1 = 32'd457
; 
32'd9858: dataIn1 = 32'd465
; 
32'd9859: dataIn1 = 32'd492
; 
32'd9860: dataIn1 = 32'd500
; 
32'd9861: dataIn1 = 32'd502
; 
32'd9862: dataIn1 = 32'd510
; 
32'd9863: dataIn1 = 32'd518
; 
32'd9864: dataIn1 = 32'd526
; 
32'd9865: dataIn1 = 32'd561
; 
32'd9866: dataIn1 = 32'd578
; 
32'd9867: dataIn1 = 32'd597
; 
32'd9868: dataIn1 = 32'd619
; 
32'd9869: dataIn1 = 32'd664
; 
32'd9870: dataIn1 = 32'd665
; 
32'd9871: dataIn1 = 32'd692
; 
32'd9872: dataIn1 = 32'd695
; 
32'd9873: dataIn1 = 32'd712
; 
32'd9874: dataIn1 = 32'd744
; 
32'd9875: dataIn1 = 32'd765
; 
32'd9876: dataIn1 = 32'd796
; 
32'd9877: dataIn1 = 32'd58
; 
32'd9878: dataIn1 = 32'd77
; 
32'd9879: dataIn1 = 32'd131
; 
32'd9880: dataIn1 = 32'd148
; 
32'd9881: dataIn1 = 32'd164
; 
32'd9882: dataIn1 = 32'd180
; 
32'd9883: dataIn1 = 32'd192
; 
32'd9884: dataIn1 = 32'd229
; 
32'd9885: dataIn1 = 32'd235
; 
32'd9886: dataIn1 = 32'd238
; 
32'd9887: dataIn1 = 32'd240
; 
32'd9888: dataIn1 = 32'd243
; 
32'd9889: dataIn1 = 32'd244
; 
32'd9890: dataIn1 = 32'd251
; 
32'd9891: dataIn1 = 32'd252
; 
32'd9892: dataIn1 = 32'd255
; 
32'd9893: dataIn1 = 32'd261
; 
32'd9894: dataIn1 = 32'd276
; 
32'd9895: dataIn1 = 32'd289
; 
32'd9896: dataIn1 = 32'd327
; 
32'd9897: dataIn1 = 32'd341
; 
32'd9898: dataIn1 = 32'd343
; 
32'd9899: dataIn1 = 32'd369
; 
32'd9900: dataIn1 = 32'd406
; 
32'd9901: dataIn1 = 32'd421
; 
32'd9902: dataIn1 = 32'd438
; 
32'd9903: dataIn1 = 32'd442
; 
32'd9904: dataIn1 = 32'd443
; 
32'd9905: dataIn1 = 32'd456
; 
32'd9906: dataIn1 = 32'd467
; 
32'd9907: dataIn1 = 32'd476
; 
32'd9908: dataIn1 = 32'd486
; 
32'd9909: dataIn1 = 32'd491
; 
32'd9910: dataIn1 = 32'd504
; 
32'd9911: dataIn1 = 32'd518
; 
32'd9912: dataIn1 = 32'd524
; 
32'd9913: dataIn1 = 32'd532
; 
32'd9914: dataIn1 = 32'd542
; 
32'd9915: dataIn1 = 32'd569
; 
32'd9916: dataIn1 = 32'd579
; 
32'd9917: dataIn1 = 32'd606
; 
32'd9918: dataIn1 = 32'd607
; 
32'd9919: dataIn1 = 32'd608
; 
32'd9920: dataIn1 = 32'd615
; 
32'd9921: dataIn1 = 32'd643
; 
32'd9922: dataIn1 = 32'd672
; 
32'd9923: dataIn1 = 32'd692
; 
32'd9924: dataIn1 = 32'd702
; 
32'd9925: dataIn1 = 32'd713
; 
32'd9926: dataIn1 = 32'd722
; 
32'd9927: dataIn1 = 32'd739
; 
32'd9928: dataIn1 = 32'd755
; 
32'd9929: dataIn1 = 32'd777
; 
32'd9930: dataIn1 = 32'd786
; 
32'd9931: dataIn1 = 32'd788
; 
32'd9932: dataIn1 = 32'd789
; 
32'd9933: dataIn1 = 32'd57
; 
32'd9934: dataIn1 = 32'd83
; 
32'd9935: dataIn1 = 32'd91
; 
32'd9936: dataIn1 = 32'd117
; 
32'd9937: dataIn1 = 32'd128
; 
32'd9938: dataIn1 = 32'd133
; 
32'd9939: dataIn1 = 32'd166
; 
32'd9940: dataIn1 = 32'd210
; 
32'd9941: dataIn1 = 32'd214
; 
32'd9942: dataIn1 = 32'd218
; 
32'd9943: dataIn1 = 32'd230
; 
32'd9944: dataIn1 = 32'd238
; 
32'd9945: dataIn1 = 32'd245
; 
32'd9946: dataIn1 = 32'd248
; 
32'd9947: dataIn1 = 32'd251
; 
32'd9948: dataIn1 = 32'd256
; 
32'd9949: dataIn1 = 32'd257
; 
32'd9950: dataIn1 = 32'd268
; 
32'd9951: dataIn1 = 32'd277
; 
32'd9952: dataIn1 = 32'd312
; 
32'd9953: dataIn1 = 32'd326
; 
32'd9954: dataIn1 = 32'd332
; 
32'd9955: dataIn1 = 32'd344
; 
32'd9956: dataIn1 = 32'd357
; 
32'd9957: dataIn1 = 32'd365
; 
32'd9958: dataIn1 = 32'd403
; 
32'd9959: dataIn1 = 32'd410
; 
32'd9960: dataIn1 = 32'd411
; 
32'd9961: dataIn1 = 32'd416
; 
32'd9962: dataIn1 = 32'd450
; 
32'd9963: dataIn1 = 32'd451
; 
32'd9964: dataIn1 = 32'd468
; 
32'd9965: dataIn1 = 32'd473
; 
32'd9966: dataIn1 = 32'd475
; 
32'd9967: dataIn1 = 32'd482
; 
32'd9968: dataIn1 = 32'd497
; 
32'd9969: dataIn1 = 32'd498
; 
32'd9970: dataIn1 = 32'd518
; 
32'd9971: dataIn1 = 32'd531
; 
32'd9972: dataIn1 = 32'd533
; 
32'd9973: dataIn1 = 32'd539
; 
32'd9974: dataIn1 = 32'd544
; 
32'd9975: dataIn1 = 32'd581
; 
32'd9976: dataIn1 = 32'd651
; 
32'd9977: dataIn1 = 32'd657
; 
32'd9978: dataIn1 = 32'd662
; 
32'd9979: dataIn1 = 32'd673
; 
32'd9980: dataIn1 = 32'd692
; 
32'd9981: dataIn1 = 32'd712
; 
32'd9982: dataIn1 = 32'd736
; 
32'd9983: dataIn1 = 32'd739
; 
32'd9984: dataIn1 = 32'd742
; 
32'd9985: dataIn1 = 32'd779
; 
32'd9986: dataIn1 = 32'd788
; 
32'd9987: dataIn1 = 32'd790
; 
32'd9988: dataIn1 = 32'd58
; 
32'd9989: dataIn1 = 32'd69
; 
32'd9990: dataIn1 = 32'd86
; 
32'd9991: dataIn1 = 32'd94
; 
32'd9992: dataIn1 = 32'd96
; 
32'd9993: dataIn1 = 32'd123
; 
32'd9994: dataIn1 = 32'd160
; 
32'd9995: dataIn1 = 32'd170
; 
32'd9996: dataIn1 = 32'd172
; 
32'd9997: dataIn1 = 32'd201
; 
32'd9998: dataIn1 = 32'd229
; 
32'd9999: dataIn1 = 32'd237
; 
32'd10000: dataIn1 = 32'd255
; 
32'd10001: dataIn1 = 32'd279
; 
32'd10002: dataIn1 = 32'd284
; 
32'd10003: dataIn1 = 32'd286
; 
32'd10004: dataIn1 = 32'd298
; 
32'd10005: dataIn1 = 32'd334
; 
32'd10006: dataIn1 = 32'd336
; 
32'd10007: dataIn1 = 32'd370
; 
32'd10008: dataIn1 = 32'd376
; 
32'd10009: dataIn1 = 32'd379
; 
32'd10010: dataIn1 = 32'd380
; 
32'd10011: dataIn1 = 32'd430
; 
32'd10012: dataIn1 = 32'd448
; 
32'd10013: dataIn1 = 32'd453
; 
32'd10014: dataIn1 = 32'd471
; 
32'd10015: dataIn1 = 32'd479
; 
32'd10016: dataIn1 = 32'd490
; 
32'd10017: dataIn1 = 32'd525
; 
32'd10018: dataIn1 = 32'd539
; 
32'd10019: dataIn1 = 32'd595
; 
32'd10020: dataIn1 = 32'd606
; 
32'd10021: dataIn1 = 32'd667
; 
32'd10022: dataIn1 = 32'd676
; 
32'd10023: dataIn1 = 32'd712
; 
32'd10024: dataIn1 = 32'd729
; 
32'd10025: dataIn1 = 32'd773
; 
32'd10026: dataIn1 = 32'd800
; 
32'd10027: dataIn1 = 32'd52
; 
32'd10028: dataIn1 = 32'd55
; 
32'd10029: dataIn1 = 32'd83
; 
32'd10030: dataIn1 = 32'd112
; 
32'd10031: dataIn1 = 32'd121
; 
32'd10032: dataIn1 = 32'd139
; 
32'd10033: dataIn1 = 32'd151
; 
32'd10034: dataIn1 = 32'd163
; 
32'd10035: dataIn1 = 32'd198
; 
32'd10036: dataIn1 = 32'd200
; 
32'd10037: dataIn1 = 32'd202
; 
32'd10038: dataIn1 = 32'd213
; 
32'd10039: dataIn1 = 32'd219
; 
32'd10040: dataIn1 = 32'd234
; 
32'd10041: dataIn1 = 32'd247
; 
32'd10042: dataIn1 = 32'd272
; 
32'd10043: dataIn1 = 32'd287
; 
32'd10044: dataIn1 = 32'd307
; 
32'd10045: dataIn1 = 32'd320
; 
32'd10046: dataIn1 = 32'd324
; 
32'd10047: dataIn1 = 32'd342
; 
32'd10048: dataIn1 = 32'd350
; 
32'd10049: dataIn1 = 32'd359
; 
32'd10050: dataIn1 = 32'd371
; 
32'd10051: dataIn1 = 32'd388
; 
32'd10052: dataIn1 = 32'd396
; 
32'd10053: dataIn1 = 32'd409
; 
32'd10054: dataIn1 = 32'd449
; 
32'd10055: dataIn1 = 32'd454
; 
32'd10056: dataIn1 = 32'd459
; 
32'd10057: dataIn1 = 32'd461
; 
32'd10058: dataIn1 = 32'd493
; 
32'd10059: dataIn1 = 32'd508
; 
32'd10060: dataIn1 = 32'd549
; 
32'd10061: dataIn1 = 32'd573
; 
32'd10062: dataIn1 = 32'd589
; 
32'd10063: dataIn1 = 32'd596
; 
32'd10064: dataIn1 = 32'd601
; 
32'd10065: dataIn1 = 32'd617
; 
32'd10066: dataIn1 = 32'd618
; 
32'd10067: dataIn1 = 32'd620
; 
32'd10068: dataIn1 = 32'd639
; 
32'd10069: dataIn1 = 32'd668
; 
32'd10070: dataIn1 = 32'd673
; 
32'd10071: dataIn1 = 32'd679
; 
32'd10072: dataIn1 = 32'd689
; 
32'd10073: dataIn1 = 32'd692
; 
32'd10074: dataIn1 = 32'd704
; 
32'd10075: dataIn1 = 32'd759
; 
32'd10076: dataIn1 = 32'd775
; 
32'd10077: dataIn1 = 32'd785
; 
32'd10078: dataIn1 = 32'd797
; 
32'd10079: dataIn1 = 32'd77
; 
32'd10080: dataIn1 = 32'd85
; 
32'd10081: dataIn1 = 32'd89
; 
32'd10082: dataIn1 = 32'd92
; 
32'd10083: dataIn1 = 32'd97
; 
32'd10084: dataIn1 = 32'd99
; 
32'd10085: dataIn1 = 32'd143
; 
32'd10086: dataIn1 = 32'd169
; 
32'd10087: dataIn1 = 32'd170
; 
32'd10088: dataIn1 = 32'd177
; 
32'd10089: dataIn1 = 32'd195
; 
32'd10090: dataIn1 = 32'd235
; 
32'd10091: dataIn1 = 32'd242
; 
32'd10092: dataIn1 = 32'd250
; 
32'd10093: dataIn1 = 32'd288
; 
32'd10094: dataIn1 = 32'd309
; 
32'd10095: dataIn1 = 32'd318
; 
32'd10096: dataIn1 = 32'd358
; 
32'd10097: dataIn1 = 32'd369
; 
32'd10098: dataIn1 = 32'd377
; 
32'd10099: dataIn1 = 32'd386
; 
32'd10100: dataIn1 = 32'd388
; 
32'd10101: dataIn1 = 32'd401
; 
32'd10102: dataIn1 = 32'd412
; 
32'd10103: dataIn1 = 32'd438
; 
32'd10104: dataIn1 = 32'd442
; 
32'd10105: dataIn1 = 32'd444
; 
32'd10106: dataIn1 = 32'd457
; 
32'd10107: dataIn1 = 32'd459
; 
32'd10108: dataIn1 = 32'd460
; 
32'd10109: dataIn1 = 32'd467
; 
32'd10110: dataIn1 = 32'd507
; 
32'd10111: dataIn1 = 32'd521
; 
32'd10112: dataIn1 = 32'd532
; 
32'd10113: dataIn1 = 32'd550
; 
32'd10114: dataIn1 = 32'd569
; 
32'd10115: dataIn1 = 32'd589
; 
32'd10116: dataIn1 = 32'd657
; 
32'd10117: dataIn1 = 32'd706
; 
32'd10118: dataIn1 = 32'd709
; 
32'd10119: dataIn1 = 32'd725
; 
32'd10120: dataIn1 = 32'd746
; 
32'd10121: dataIn1 = 32'd758
; 
32'd10122: dataIn1 = 32'd769
; 
32'd10123: dataIn1 = 32'd779
; 
32'd10124: dataIn1 = 32'd783
; 
32'd10125: dataIn1 = 32'd784
; 
32'd10126: dataIn1 = 32'd792
; 
32'd10127: dataIn1 = 32'd60
; 
32'd10128: dataIn1 = 32'd61
; 
32'd10129: dataIn1 = 32'd62
; 
32'd10130: dataIn1 = 32'd63
; 
32'd10131: dataIn1 = 32'd80
; 
32'd10132: dataIn1 = 32'd139
; 
32'd10133: dataIn1 = 32'd141
; 
32'd10134: dataIn1 = 32'd168
; 
32'd10135: dataIn1 = 32'd171
; 
32'd10136: dataIn1 = 32'd201
; 
32'd10137: dataIn1 = 32'd231
; 
32'd10138: dataIn1 = 32'd233
; 
32'd10139: dataIn1 = 32'd240
; 
32'd10140: dataIn1 = 32'd267
; 
32'd10141: dataIn1 = 32'd270
; 
32'd10142: dataIn1 = 32'd277
; 
32'd10143: dataIn1 = 32'd311
; 
32'd10144: dataIn1 = 32'd313
; 
32'd10145: dataIn1 = 32'd323
; 
32'd10146: dataIn1 = 32'd341
; 
32'd10147: dataIn1 = 32'd352
; 
32'd10148: dataIn1 = 32'd357
; 
32'd10149: dataIn1 = 32'd379
; 
32'd10150: dataIn1 = 32'd390
; 
32'd10151: dataIn1 = 32'd399
; 
32'd10152: dataIn1 = 32'd406
; 
32'd10153: dataIn1 = 32'd408
; 
32'd10154: dataIn1 = 32'd476
; 
32'd10155: dataIn1 = 32'd484
; 
32'd10156: dataIn1 = 32'd502
; 
32'd10157: dataIn1 = 32'd504
; 
32'd10158: dataIn1 = 32'd517
; 
32'd10159: dataIn1 = 32'd528
; 
32'd10160: dataIn1 = 32'd534
; 
32'd10161: dataIn1 = 32'd537
; 
32'd10162: dataIn1 = 32'd541
; 
32'd10163: dataIn1 = 32'd542
; 
32'd10164: dataIn1 = 32'd553
; 
32'd10165: dataIn1 = 32'd566
; 
32'd10166: dataIn1 = 32'd586
; 
32'd10167: dataIn1 = 32'd603
; 
32'd10168: dataIn1 = 32'd628
; 
32'd10169: dataIn1 = 32'd630
; 
32'd10170: dataIn1 = 32'd641
; 
32'd10171: dataIn1 = 32'd642
; 
32'd10172: dataIn1 = 32'd651
; 
32'd10173: dataIn1 = 32'd681
; 
32'd10174: dataIn1 = 32'd693
; 
32'd10175: dataIn1 = 32'd700
; 
32'd10176: dataIn1 = 32'd705
; 
32'd10177: dataIn1 = 32'd710
; 
32'd10178: dataIn1 = 32'd732
; 
32'd10179: dataIn1 = 32'd733
; 
32'd10180: dataIn1 = 32'd734
; 
32'd10181: dataIn1 = 32'd747
; 
32'd10182: dataIn1 = 32'd768
; 
32'd10183: dataIn1 = 32'd776
; 
32'd10184: dataIn1 = 32'd799
; 
32'd10185: dataIn1 = 32'd50
; 
32'd10186: dataIn1 = 32'd58
; 
32'd10187: dataIn1 = 32'd86
; 
32'd10188: dataIn1 = 32'd100
; 
32'd10189: dataIn1 = 32'd107
; 
32'd10190: dataIn1 = 32'd109
; 
32'd10191: dataIn1 = 32'd116
; 
32'd10192: dataIn1 = 32'd119
; 
32'd10193: dataIn1 = 32'd120
; 
32'd10194: dataIn1 = 32'd155
; 
32'd10195: dataIn1 = 32'd162
; 
32'd10196: dataIn1 = 32'd168
; 
32'd10197: dataIn1 = 32'd178
; 
32'd10198: dataIn1 = 32'd193
; 
32'd10199: dataIn1 = 32'd246
; 
32'd10200: dataIn1 = 32'd252
; 
32'd10201: dataIn1 = 32'd267
; 
32'd10202: dataIn1 = 32'd292
; 
32'd10203: dataIn1 = 32'd313
; 
32'd10204: dataIn1 = 32'd314
; 
32'd10205: dataIn1 = 32'd337
; 
32'd10206: dataIn1 = 32'd355
; 
32'd10207: dataIn1 = 32'd365
; 
32'd10208: dataIn1 = 32'd401
; 
32'd10209: dataIn1 = 32'd402
; 
32'd10210: dataIn1 = 32'd421
; 
32'd10211: dataIn1 = 32'd453
; 
32'd10212: dataIn1 = 32'd483
; 
32'd10213: dataIn1 = 32'd485
; 
32'd10214: dataIn1 = 32'd505
; 
32'd10215: dataIn1 = 32'd538
; 
32'd10216: dataIn1 = 32'd557
; 
32'd10217: dataIn1 = 32'd587
; 
32'd10218: dataIn1 = 32'd613
; 
32'd10219: dataIn1 = 32'd701
; 
32'd10220: dataIn1 = 32'd720
; 
32'd10221: dataIn1 = 32'd721
; 
32'd10222: dataIn1 = 32'd735
; 
32'd10223: dataIn1 = 32'd742
; 
32'd10224: dataIn1 = 32'd772
; 
32'd10225: dataIn1 = 32'd777
; 
32'd10226: dataIn1 = 32'd779
; 
32'd10227: dataIn1 = 32'd99
; 
32'd10228: dataIn1 = 32'd100
; 
32'd10229: dataIn1 = 32'd153
; 
32'd10230: dataIn1 = 32'd166
; 
32'd10231: dataIn1 = 32'd182
; 
32'd10232: dataIn1 = 32'd206
; 
32'd10233: dataIn1 = 32'd209
; 
32'd10234: dataIn1 = 32'd216
; 
32'd10235: dataIn1 = 32'd221
; 
32'd10236: dataIn1 = 32'd230
; 
32'd10237: dataIn1 = 32'd234
; 
32'd10238: dataIn1 = 32'd278
; 
32'd10239: dataIn1 = 32'd279
; 
32'd10240: dataIn1 = 32'd316
; 
32'd10241: dataIn1 = 32'd318
; 
32'd10242: dataIn1 = 32'd335
; 
32'd10243: dataIn1 = 32'd357
; 
32'd10244: dataIn1 = 32'd371
; 
32'd10245: dataIn1 = 32'd413
; 
32'd10246: dataIn1 = 32'd416
; 
32'd10247: dataIn1 = 32'd445
; 
32'd10248: dataIn1 = 32'd446
; 
32'd10249: dataIn1 = 32'd468
; 
32'd10250: dataIn1 = 32'd478
; 
32'd10251: dataIn1 = 32'd481
; 
32'd10252: dataIn1 = 32'd512
; 
32'd10253: dataIn1 = 32'd531
; 
32'd10254: dataIn1 = 32'd535
; 
32'd10255: dataIn1 = 32'd538
; 
32'd10256: dataIn1 = 32'd564
; 
32'd10257: dataIn1 = 32'd588
; 
32'd10258: dataIn1 = 32'd599
; 
32'd10259: dataIn1 = 32'd613
; 
32'd10260: dataIn1 = 32'd627
; 
32'd10261: dataIn1 = 32'd636
; 
32'd10262: dataIn1 = 32'd665
; 
32'd10263: dataIn1 = 32'd670
; 
32'd10264: dataIn1 = 32'd707
; 
32'd10265: dataIn1 = 32'd759
; 
32'd10266: dataIn1 = 32'd790
; 
32'd10267: dataIn1 = 32'd795
; 
32'd10268: dataIn1 = 32'd93
; 
32'd10269: dataIn1 = 32'd127
; 
32'd10270: dataIn1 = 32'd189
; 
32'd10271: dataIn1 = 32'd207
; 
32'd10272: dataIn1 = 32'd211
; 
32'd10273: dataIn1 = 32'd236
; 
32'd10274: dataIn1 = 32'd258
; 
32'd10275: dataIn1 = 32'd262
; 
32'd10276: dataIn1 = 32'd302
; 
32'd10277: dataIn1 = 32'd330
; 
32'd10278: dataIn1 = 32'd348
; 
32'd10279: dataIn1 = 32'd426
; 
32'd10280: dataIn1 = 32'd469
; 
32'd10281: dataIn1 = 32'd471
; 
32'd10282: dataIn1 = 32'd521
; 
32'd10283: dataIn1 = 32'd523
; 
32'd10284: dataIn1 = 32'd533
; 
32'd10285: dataIn1 = 32'd557
; 
32'd10286: dataIn1 = 32'd563
; 
32'd10287: dataIn1 = 32'd586
; 
32'd10288: dataIn1 = 32'd587
; 
32'd10289: dataIn1 = 32'd596
; 
32'd10290: dataIn1 = 32'd597
; 
32'd10291: dataIn1 = 32'd633
; 
32'd10292: dataIn1 = 32'd674
; 
32'd10293: dataIn1 = 32'd706
; 
32'd10294: dataIn1 = 32'd707
; 
32'd10295: dataIn1 = 32'd749
; 
32'd10296: dataIn1 = 32'd750
; 
32'd10297: dataIn1 = 32'd793
; 
32'd10298: dataIn1 = 32'd798
; 
32'd10299: dataIn1 = 32'd799
; 
32'd10300: dataIn1 = 32'd58
; 
32'd10301: dataIn1 = 32'd78
; 
32'd10302: dataIn1 = 32'd81
; 
32'd10303: dataIn1 = 32'd99
; 
32'd10304: dataIn1 = 32'd130
; 
32'd10305: dataIn1 = 32'd151
; 
32'd10306: dataIn1 = 32'd169
; 
32'd10307: dataIn1 = 32'd171
; 
32'd10308: dataIn1 = 32'd172
; 
32'd10309: dataIn1 = 32'd173
; 
32'd10310: dataIn1 = 32'd179
; 
32'd10311: dataIn1 = 32'd222
; 
32'd10312: dataIn1 = 32'd226
; 
32'd10313: dataIn1 = 32'd230
; 
32'd10314: dataIn1 = 32'd246
; 
32'd10315: dataIn1 = 32'd248
; 
32'd10316: dataIn1 = 32'd321
; 
32'd10317: dataIn1 = 32'd328
; 
32'd10318: dataIn1 = 32'd337
; 
32'd10319: dataIn1 = 32'd340
; 
32'd10320: dataIn1 = 32'd378
; 
32'd10321: dataIn1 = 32'd441
; 
32'd10322: dataIn1 = 32'd448
; 
32'd10323: dataIn1 = 32'd463
; 
32'd10324: dataIn1 = 32'd474
; 
32'd10325: dataIn1 = 32'd484
; 
32'd10326: dataIn1 = 32'd488
; 
32'd10327: dataIn1 = 32'd490
; 
32'd10328: dataIn1 = 32'd492
; 
32'd10329: dataIn1 = 32'd519
; 
32'd10330: dataIn1 = 32'd520
; 
32'd10331: dataIn1 = 32'd552
; 
32'd10332: dataIn1 = 32'd566
; 
32'd10333: dataIn1 = 32'd584
; 
32'd10334: dataIn1 = 32'd617
; 
32'd10335: dataIn1 = 32'd627
; 
32'd10336: dataIn1 = 32'd632
; 
32'd10337: dataIn1 = 32'd637
; 
32'd10338: dataIn1 = 32'd642
; 
32'd10339: dataIn1 = 32'd649
; 
32'd10340: dataIn1 = 32'd655
; 
32'd10341: dataIn1 = 32'd665
; 
32'd10342: dataIn1 = 32'd678
; 
32'd10343: dataIn1 = 32'd680
; 
32'd10344: dataIn1 = 32'd740
; 
32'd10345: dataIn1 = 32'd753
; 
32'd10346: dataIn1 = 32'd775
; 
32'd10347: dataIn1 = 32'd781
; 
32'd10348: dataIn1 = 32'd783
; 
32'd10349: dataIn1 = 32'd789
; 
32'd10350: dataIn1 = 32'd71
; 
32'd10351: dataIn1 = 32'd80
; 
32'd10352: dataIn1 = 32'd92
; 
32'd10353: dataIn1 = 32'd104
; 
32'd10354: dataIn1 = 32'd116
; 
32'd10355: dataIn1 = 32'd118
; 
32'd10356: dataIn1 = 32'd135
; 
32'd10357: dataIn1 = 32'd139
; 
32'd10358: dataIn1 = 32'd170
; 
32'd10359: dataIn1 = 32'd219
; 
32'd10360: dataIn1 = 32'd229
; 
32'd10361: dataIn1 = 32'd242
; 
32'd10362: dataIn1 = 32'd247
; 
32'd10363: dataIn1 = 32'd310
; 
32'd10364: dataIn1 = 32'd324
; 
32'd10365: dataIn1 = 32'd339
; 
32'd10366: dataIn1 = 32'd342
; 
32'd10367: dataIn1 = 32'd354
; 
32'd10368: dataIn1 = 32'd389
; 
32'd10369: dataIn1 = 32'd393
; 
32'd10370: dataIn1 = 32'd404
; 
32'd10371: dataIn1 = 32'd407
; 
32'd10372: dataIn1 = 32'd415
; 
32'd10373: dataIn1 = 32'd422
; 
32'd10374: dataIn1 = 32'd448
; 
32'd10375: dataIn1 = 32'd455
; 
32'd10376: dataIn1 = 32'd476
; 
32'd10377: dataIn1 = 32'd485
; 
32'd10378: dataIn1 = 32'd498
; 
32'd10379: dataIn1 = 32'd528
; 
32'd10380: dataIn1 = 32'd541
; 
32'd10381: dataIn1 = 32'd596
; 
32'd10382: dataIn1 = 32'd605
; 
32'd10383: dataIn1 = 32'd647
; 
32'd10384: dataIn1 = 32'd659
; 
32'd10385: dataIn1 = 32'd683
; 
32'd10386: dataIn1 = 32'd696
; 
32'd10387: dataIn1 = 32'd706
; 
32'd10388: dataIn1 = 32'd715
; 
32'd10389: dataIn1 = 32'd733
; 
32'd10390: dataIn1 = 32'd736
; 
32'd10391: dataIn1 = 32'd751
; 
32'd10392: dataIn1 = 32'd776
; 
32'd10393: dataIn1 = 32'd783
; 
32'd10394: dataIn1 = 32'd791
; 
32'd10395: dataIn1 = 32'd792
; 
32'd10396: dataIn1 = 32'd795
; 
32'd10397: dataIn1 = 32'd800
; 
32'd10398: dataIn1 = 32'd61
; 
32'd10399: dataIn1 = 32'd83
; 
32'd10400: dataIn1 = 32'd125
; 
32'd10401: dataIn1 = 32'd135
; 
32'd10402: dataIn1 = 32'd181
; 
32'd10403: dataIn1 = 32'd208
; 
32'd10404: dataIn1 = 32'd221
; 
32'd10405: dataIn1 = 32'd239
; 
32'd10406: dataIn1 = 32'd262
; 
32'd10407: dataIn1 = 32'd267
; 
32'd10408: dataIn1 = 32'd276
; 
32'd10409: dataIn1 = 32'd278
; 
32'd10410: dataIn1 = 32'd361
; 
32'd10411: dataIn1 = 32'd367
; 
32'd10412: dataIn1 = 32'd452
; 
32'd10413: dataIn1 = 32'd457
; 
32'd10414: dataIn1 = 32'd458
; 
32'd10415: dataIn1 = 32'd463
; 
32'd10416: dataIn1 = 32'd510
; 
32'd10417: dataIn1 = 32'd530
; 
32'd10418: dataIn1 = 32'd559
; 
32'd10419: dataIn1 = 32'd564
; 
32'd10420: dataIn1 = 32'd592
; 
32'd10421: dataIn1 = 32'd595
; 
32'd10422: dataIn1 = 32'd604
; 
32'd10423: dataIn1 = 32'd605
; 
32'd10424: dataIn1 = 32'd612
; 
32'd10425: dataIn1 = 32'd625
; 
32'd10426: dataIn1 = 32'd626
; 
32'd10427: dataIn1 = 32'd652
; 
32'd10428: dataIn1 = 32'd672
; 
32'd10429: dataIn1 = 32'd677
; 
32'd10430: dataIn1 = 32'd688
; 
32'd10431: dataIn1 = 32'd689
; 
32'd10432: dataIn1 = 32'd708
; 
32'd10433: dataIn1 = 32'd717
; 
32'd10434: dataIn1 = 32'd743
; 
32'd10435: dataIn1 = 32'd748
; 
32'd10436: dataIn1 = 32'd768
; 
32'd10437: dataIn1 = 32'd772
; 
32'd10438: dataIn1 = 32'd55
; 
32'd10439: dataIn1 = 32'd81
; 
32'd10440: dataIn1 = 32'd82
; 
32'd10441: dataIn1 = 32'd85
; 
32'd10442: dataIn1 = 32'd108
; 
32'd10443: dataIn1 = 32'd134
; 
32'd10444: dataIn1 = 32'd141
; 
32'd10445: dataIn1 = 32'd161
; 
32'd10446: dataIn1 = 32'd182
; 
32'd10447: dataIn1 = 32'd192
; 
32'd10448: dataIn1 = 32'd244
; 
32'd10449: dataIn1 = 32'd245
; 
32'd10450: dataIn1 = 32'd261
; 
32'd10451: dataIn1 = 32'd266
; 
32'd10452: dataIn1 = 32'd269
; 
32'd10453: dataIn1 = 32'd302
; 
32'd10454: dataIn1 = 32'd332
; 
32'd10455: dataIn1 = 32'd333
; 
32'd10456: dataIn1 = 32'd341
; 
32'd10457: dataIn1 = 32'd347
; 
32'd10458: dataIn1 = 32'd362
; 
32'd10459: dataIn1 = 32'd394
; 
32'd10460: dataIn1 = 32'd454
; 
32'd10461: dataIn1 = 32'd455
; 
32'd10462: dataIn1 = 32'd461
; 
32'd10463: dataIn1 = 32'd482
; 
32'd10464: dataIn1 = 32'd487
; 
32'd10465: dataIn1 = 32'd491
; 
32'd10466: dataIn1 = 32'd530
; 
32'd10467: dataIn1 = 32'd550
; 
32'd10468: dataIn1 = 32'd558
; 
32'd10469: dataIn1 = 32'd575
; 
32'd10470: dataIn1 = 32'd648
; 
32'd10471: dataIn1 = 32'd660
; 
32'd10472: dataIn1 = 32'd662
; 
32'd10473: dataIn1 = 32'd670
; 
32'd10474: dataIn1 = 32'd687
; 
32'd10475: dataIn1 = 32'd697
; 
32'd10476: dataIn1 = 32'd699
; 
32'd10477: dataIn1 = 32'd738
; 
32'd10478: dataIn1 = 32'd764
; 
32'd10479: dataIn1 = 32'd780
; 
32'd10480: dataIn1 = 32'd62
; 
32'd10481: dataIn1 = 32'd68
; 
32'd10482: dataIn1 = 32'd77
; 
32'd10483: dataIn1 = 32'd83
; 
32'd10484: dataIn1 = 32'd101
; 
32'd10485: dataIn1 = 32'd124
; 
32'd10486: dataIn1 = 32'd127
; 
32'd10487: dataIn1 = 32'd139
; 
32'd10488: dataIn1 = 32'd147
; 
32'd10489: dataIn1 = 32'd148
; 
32'd10490: dataIn1 = 32'd151
; 
32'd10491: dataIn1 = 32'd157
; 
32'd10492: dataIn1 = 32'd177
; 
32'd10493: dataIn1 = 32'd181
; 
32'd10494: dataIn1 = 32'd206
; 
32'd10495: dataIn1 = 32'd211
; 
32'd10496: dataIn1 = 32'd217
; 
32'd10497: dataIn1 = 32'd223
; 
32'd10498: dataIn1 = 32'd226
; 
32'd10499: dataIn1 = 32'd245
; 
32'd10500: dataIn1 = 32'd246
; 
32'd10501: dataIn1 = 32'd254
; 
32'd10502: dataIn1 = 32'd261
; 
32'd10503: dataIn1 = 32'd265
; 
32'd10504: dataIn1 = 32'd282
; 
32'd10505: dataIn1 = 32'd333
; 
32'd10506: dataIn1 = 32'd337
; 
32'd10507: dataIn1 = 32'd357
; 
32'd10508: dataIn1 = 32'd407
; 
32'd10509: dataIn1 = 32'd426
; 
32'd10510: dataIn1 = 32'd428
; 
32'd10511: dataIn1 = 32'd437
; 
32'd10512: dataIn1 = 32'd452
; 
32'd10513: dataIn1 = 32'd461
; 
32'd10514: dataIn1 = 32'd471
; 
32'd10515: dataIn1 = 32'd475
; 
32'd10516: dataIn1 = 32'd545
; 
32'd10517: dataIn1 = 32'd549
; 
32'd10518: dataIn1 = 32'd552
; 
32'd10519: dataIn1 = 32'd569
; 
32'd10520: dataIn1 = 32'd570
; 
32'd10521: dataIn1 = 32'd573
; 
32'd10522: dataIn1 = 32'd586
; 
32'd10523: dataIn1 = 32'd604
; 
32'd10524: dataIn1 = 32'd608
; 
32'd10525: dataIn1 = 32'd631
; 
32'd10526: dataIn1 = 32'd635
; 
32'd10527: dataIn1 = 32'd641
; 
32'd10528: dataIn1 = 32'd642
; 
32'd10529: dataIn1 = 32'd649
; 
32'd10530: dataIn1 = 32'd664
; 
32'd10531: dataIn1 = 32'd676
; 
32'd10532: dataIn1 = 32'd683
; 
32'd10533: dataIn1 = 32'd685
; 
32'd10534: dataIn1 = 32'd708
; 
32'd10535: dataIn1 = 32'd747
; 
32'd10536: dataIn1 = 32'd750
; 
32'd10537: dataIn1 = 32'd782
; 
32'd10538: dataIn1 = 32'd800
; 
32'd10539: dataIn1 = 32'd75
; 
32'd10540: dataIn1 = 32'd91
; 
32'd10541: dataIn1 = 32'd112
; 
32'd10542: dataIn1 = 32'd120
; 
32'd10543: dataIn1 = 32'd203
; 
32'd10544: dataIn1 = 32'd211
; 
32'd10545: dataIn1 = 32'd212
; 
32'd10546: dataIn1 = 32'd234
; 
32'd10547: dataIn1 = 32'd251
; 
32'd10548: dataIn1 = 32'd272
; 
32'd10549: dataIn1 = 32'd285
; 
32'd10550: dataIn1 = 32'd296
; 
32'd10551: dataIn1 = 32'd305
; 
32'd10552: dataIn1 = 32'd316
; 
32'd10553: dataIn1 = 32'd340
; 
32'd10554: dataIn1 = 32'd347
; 
32'd10555: dataIn1 = 32'd355
; 
32'd10556: dataIn1 = 32'd366
; 
32'd10557: dataIn1 = 32'd378
; 
32'd10558: dataIn1 = 32'd419
; 
32'd10559: dataIn1 = 32'd434
; 
32'd10560: dataIn1 = 32'd435
; 
32'd10561: dataIn1 = 32'd450
; 
32'd10562: dataIn1 = 32'd457
; 
32'd10563: dataIn1 = 32'd464
; 
32'd10564: dataIn1 = 32'd491
; 
32'd10565: dataIn1 = 32'd496
; 
32'd10566: dataIn1 = 32'd518
; 
32'd10567: dataIn1 = 32'd528
; 
32'd10568: dataIn1 = 32'd540
; 
32'd10569: dataIn1 = 32'd547
; 
32'd10570: dataIn1 = 32'd581
; 
32'd10571: dataIn1 = 32'd586
; 
32'd10572: dataIn1 = 32'd602
; 
32'd10573: dataIn1 = 32'd668
; 
32'd10574: dataIn1 = 32'd690
; 
32'd10575: dataIn1 = 32'd709
; 
32'd10576: dataIn1 = 32'd720
; 
32'd10577: dataIn1 = 32'd735
; 
32'd10578: dataIn1 = 32'd738
; 
32'd10579: dataIn1 = 32'd764
; 
32'd10580: dataIn1 = 32'd776
; 
32'd10581: dataIn1 = 32'd58
; 
32'd10582: dataIn1 = 32'd72
; 
32'd10583: dataIn1 = 32'd89
; 
32'd10584: dataIn1 = 32'd138
; 
32'd10585: dataIn1 = 32'd153
; 
32'd10586: dataIn1 = 32'd167
; 
32'd10587: dataIn1 = 32'd174
; 
32'd10588: dataIn1 = 32'd175
; 
32'd10589: dataIn1 = 32'd201
; 
32'd10590: dataIn1 = 32'd272
; 
32'd10591: dataIn1 = 32'd286
; 
32'd10592: dataIn1 = 32'd314
; 
32'd10593: dataIn1 = 32'd374
; 
32'd10594: dataIn1 = 32'd402
; 
32'd10595: dataIn1 = 32'd409
; 
32'd10596: dataIn1 = 32'd466
; 
32'd10597: dataIn1 = 32'd478
; 
32'd10598: dataIn1 = 32'd486
; 
32'd10599: dataIn1 = 32'd503
; 
32'd10600: dataIn1 = 32'd509
; 
32'd10601: dataIn1 = 32'd517
; 
32'd10602: dataIn1 = 32'd530
; 
32'd10603: dataIn1 = 32'd550
; 
32'd10604: dataIn1 = 32'd561
; 
32'd10605: dataIn1 = 32'd574
; 
32'd10606: dataIn1 = 32'd592
; 
32'd10607: dataIn1 = 32'd603
; 
32'd10608: dataIn1 = 32'd656
; 
32'd10609: dataIn1 = 32'd668
; 
32'd10610: dataIn1 = 32'd745
; 
32'd10611: dataIn1 = 32'd750
; 
32'd10612: dataIn1 = 32'd769
; 
32'd10613: dataIn1 = 32'd772
; 
32'd10614: dataIn1 = 32'd788
; 
32'd10615: dataIn1 = 32'd140
; 
32'd10616: dataIn1 = 32'd145
; 
32'd10617: dataIn1 = 32'd153
; 
32'd10618: dataIn1 = 32'd158
; 
32'd10619: dataIn1 = 32'd169
; 
32'd10620: dataIn1 = 32'd178
; 
32'd10621: dataIn1 = 32'd208
; 
32'd10622: dataIn1 = 32'd213
; 
32'd10623: dataIn1 = 32'd259
; 
32'd10624: dataIn1 = 32'd309
; 
32'd10625: dataIn1 = 32'd344
; 
32'd10626: dataIn1 = 32'd355
; 
32'd10627: dataIn1 = 32'd379
; 
32'd10628: dataIn1 = 32'd415
; 
32'd10629: dataIn1 = 32'd464
; 
32'd10630: dataIn1 = 32'd493
; 
32'd10631: dataIn1 = 32'd520
; 
32'd10632: dataIn1 = 32'd544
; 
32'd10633: dataIn1 = 32'd556
; 
32'd10634: dataIn1 = 32'd577
; 
32'd10635: dataIn1 = 32'd588
; 
32'd10636: dataIn1 = 32'd590
; 
32'd10637: dataIn1 = 32'd612
; 
32'd10638: dataIn1 = 32'd646
; 
32'd10639: dataIn1 = 32'd688
; 
32'd10640: dataIn1 = 32'd689
; 
32'd10641: dataIn1 = 32'd698
; 
32'd10642: dataIn1 = 32'd707
; 
32'd10643: dataIn1 = 32'd715
; 
32'd10644: dataIn1 = 32'd717
; 
32'd10645: dataIn1 = 32'd719
; 
32'd10646: dataIn1 = 32'd743
; 
32'd10647: dataIn1 = 32'd756
; 
32'd10648: dataIn1 = 32'd77
; 
32'd10649: dataIn1 = 32'd109
; 
32'd10650: dataIn1 = 32'd117
; 
32'd10651: dataIn1 = 32'd121
; 
32'd10652: dataIn1 = 32'd146
; 
32'd10653: dataIn1 = 32'd149
; 
32'd10654: dataIn1 = 32'd175
; 
32'd10655: dataIn1 = 32'd188
; 
32'd10656: dataIn1 = 32'd189
; 
32'd10657: dataIn1 = 32'd198
; 
32'd10658: dataIn1 = 32'd203
; 
32'd10659: dataIn1 = 32'd243
; 
32'd10660: dataIn1 = 32'd246
; 
32'd10661: dataIn1 = 32'd258
; 
32'd10662: dataIn1 = 32'd263
; 
32'd10663: dataIn1 = 32'd283
; 
32'd10664: dataIn1 = 32'd285
; 
32'd10665: dataIn1 = 32'd295
; 
32'd10666: dataIn1 = 32'd299
; 
32'd10667: dataIn1 = 32'd309
; 
32'd10668: dataIn1 = 32'd353
; 
32'd10669: dataIn1 = 32'd378
; 
32'd10670: dataIn1 = 32'd382
; 
32'd10671: dataIn1 = 32'd395
; 
32'd10672: dataIn1 = 32'd398
; 
32'd10673: dataIn1 = 32'd406
; 
32'd10674: dataIn1 = 32'd422
; 
32'd10675: dataIn1 = 32'd456
; 
32'd10676: dataIn1 = 32'd479
; 
32'd10677: dataIn1 = 32'd489
; 
32'd10678: dataIn1 = 32'd521
; 
32'd10679: dataIn1 = 32'd541
; 
32'd10680: dataIn1 = 32'd567
; 
32'd10681: dataIn1 = 32'd595
; 
32'd10682: dataIn1 = 32'd596
; 
32'd10683: dataIn1 = 32'd605
; 
32'd10684: dataIn1 = 32'd633
; 
32'd10685: dataIn1 = 32'd643
; 
32'd10686: dataIn1 = 32'd679
; 
32'd10687: dataIn1 = 32'd730
; 
32'd10688: dataIn1 = 32'd742
; 
32'd10689: dataIn1 = 32'd745
; 
32'd10690: dataIn1 = 32'd756
; 
32'd10691: dataIn1 = 32'd790
; 
32'd10692: dataIn1 = 32'd61
; 
32'd10693: dataIn1 = 32'd82
; 
32'd10694: dataIn1 = 32'd101
; 
32'd10695: dataIn1 = 32'd129
; 
32'd10696: dataIn1 = 32'd141
; 
32'd10697: dataIn1 = 32'd175
; 
32'd10698: dataIn1 = 32'd199
; 
32'd10699: dataIn1 = 32'd202
; 
32'd10700: dataIn1 = 32'd206
; 
32'd10701: dataIn1 = 32'd235
; 
32'd10702: dataIn1 = 32'd259
; 
32'd10703: dataIn1 = 32'd285
; 
32'd10704: dataIn1 = 32'd319
; 
32'd10705: dataIn1 = 32'd359
; 
32'd10706: dataIn1 = 32'd380
; 
32'd10707: dataIn1 = 32'd394
; 
32'd10708: dataIn1 = 32'd402
; 
32'd10709: dataIn1 = 32'd404
; 
32'd10710: dataIn1 = 32'd431
; 
32'd10711: dataIn1 = 32'd439
; 
32'd10712: dataIn1 = 32'd440
; 
32'd10713: dataIn1 = 32'd458
; 
32'd10714: dataIn1 = 32'd466
; 
32'd10715: dataIn1 = 32'd491
; 
32'd10716: dataIn1 = 32'd495
; 
32'd10717: dataIn1 = 32'd559
; 
32'd10718: dataIn1 = 32'd561
; 
32'd10719: dataIn1 = 32'd566
; 
32'd10720: dataIn1 = 32'd575
; 
32'd10721: dataIn1 = 32'd617
; 
32'd10722: dataIn1 = 32'd678
; 
32'd10723: dataIn1 = 32'd679
; 
32'd10724: dataIn1 = 32'd685
; 
32'd10725: dataIn1 = 32'd698
; 
32'd10726: dataIn1 = 32'd702
; 
32'd10727: dataIn1 = 32'd721
; 
32'd10728: dataIn1 = 32'd785
; 
32'd10729: dataIn1 = 32'd63
; 
32'd10730: dataIn1 = 32'd78
; 
32'd10731: dataIn1 = 32'd85
; 
32'd10732: dataIn1 = 32'd93
; 
32'd10733: dataIn1 = 32'd108
; 
32'd10734: dataIn1 = 32'd134
; 
32'd10735: dataIn1 = 32'd183
; 
32'd10736: dataIn1 = 32'd196
; 
32'd10737: dataIn1 = 32'd210
; 
32'd10738: dataIn1 = 32'd211
; 
32'd10739: dataIn1 = 32'd312
; 
32'd10740: dataIn1 = 32'd327
; 
32'd10741: dataIn1 = 32'd348
; 
32'd10742: dataIn1 = 32'd353
; 
32'd10743: dataIn1 = 32'd358
; 
32'd10744: dataIn1 = 32'd394
; 
32'd10745: dataIn1 = 32'd441
; 
32'd10746: dataIn1 = 32'd474
; 
32'd10747: dataIn1 = 32'd489
; 
32'd10748: dataIn1 = 32'd498
; 
32'd10749: dataIn1 = 32'd503
; 
32'd10750: dataIn1 = 32'd519
; 
32'd10751: dataIn1 = 32'd525
; 
32'd10752: dataIn1 = 32'd527
; 
32'd10753: dataIn1 = 32'd556
; 
32'd10754: dataIn1 = 32'd573
; 
32'd10755: dataIn1 = 32'd612
; 
32'd10756: dataIn1 = 32'd617
; 
32'd10757: dataIn1 = 32'd632
; 
32'd10758: dataIn1 = 32'd635
; 
32'd10759: dataIn1 = 32'd670
; 
32'd10760: dataIn1 = 32'd676
; 
32'd10761: dataIn1 = 32'd681
; 
32'd10762: dataIn1 = 32'd698
; 
32'd10763: dataIn1 = 32'd702
; 
32'd10764: dataIn1 = 32'd707
; 
32'd10765: dataIn1 = 32'd725
; 
32'd10766: dataIn1 = 32'd767
; 
32'd10767: dataIn1 = 32'd775
; 
32'd10768: dataIn1 = 32'd783
; 
32'd10769: dataIn1 = 32'd795
; 
32'd10770: dataIn1 = 32'd72
; 
32'd10771: dataIn1 = 32'd89
; 
32'd10772: dataIn1 = 32'd144
; 
32'd10773: dataIn1 = 32'd167
; 
32'd10774: dataIn1 = 32'd195
; 
32'd10775: dataIn1 = 32'd199
; 
32'd10776: dataIn1 = 32'd221
; 
32'd10777: dataIn1 = 32'd266
; 
32'd10778: dataIn1 = 32'd273
; 
32'd10779: dataIn1 = 32'd287
; 
32'd10780: dataIn1 = 32'd303
; 
32'd10781: dataIn1 = 32'd343
; 
32'd10782: dataIn1 = 32'd378
; 
32'd10783: dataIn1 = 32'd383
; 
32'd10784: dataIn1 = 32'd388
; 
32'd10785: dataIn1 = 32'd406
; 
32'd10786: dataIn1 = 32'd409
; 
32'd10787: dataIn1 = 32'd425
; 
32'd10788: dataIn1 = 32'd428
; 
32'd10789: dataIn1 = 32'd433
; 
32'd10790: dataIn1 = 32'd437
; 
32'd10791: dataIn1 = 32'd470
; 
32'd10792: dataIn1 = 32'd518
; 
32'd10793: dataIn1 = 32'd537
; 
32'd10794: dataIn1 = 32'd560
; 
32'd10795: dataIn1 = 32'd566
; 
32'd10796: dataIn1 = 32'd612
; 
32'd10797: dataIn1 = 32'd626
; 
32'd10798: dataIn1 = 32'd636
; 
32'd10799: dataIn1 = 32'd637
; 
32'd10800: dataIn1 = 32'd641
; 
32'd10801: dataIn1 = 32'd684
; 
32'd10802: dataIn1 = 32'd693
; 
32'd10803: dataIn1 = 32'd717
; 
32'd10804: dataIn1 = 32'd789
; 
32'd10805: dataIn1 = 32'd797
; 
32'd10806: dataIn1 = 32'd800
; 
32'd10807: dataIn1 = 32'd72
; 
32'd10808: dataIn1 = 32'd107
; 
32'd10809: dataIn1 = 32'd127
; 
32'd10810: dataIn1 = 32'd142
; 
32'd10811: dataIn1 = 32'd181
; 
32'd10812: dataIn1 = 32'd184
; 
32'd10813: dataIn1 = 32'd190
; 
32'd10814: dataIn1 = 32'd209
; 
32'd10815: dataIn1 = 32'd210
; 
32'd10816: dataIn1 = 32'd240
; 
32'd10817: dataIn1 = 32'd286
; 
32'd10818: dataIn1 = 32'd307
; 
32'd10819: dataIn1 = 32'd312
; 
32'd10820: dataIn1 = 32'd335
; 
32'd10821: dataIn1 = 32'd341
; 
32'd10822: dataIn1 = 32'd346
; 
32'd10823: dataIn1 = 32'd354
; 
32'd10824: dataIn1 = 32'd382
; 
32'd10825: dataIn1 = 32'd430
; 
32'd10826: dataIn1 = 32'd440
; 
32'd10827: dataIn1 = 32'd506
; 
32'd10828: dataIn1 = 32'd541
; 
32'd10829: dataIn1 = 32'd562
; 
32'd10830: dataIn1 = 32'd577
; 
32'd10831: dataIn1 = 32'd580
; 
32'd10832: dataIn1 = 32'd587
; 
32'd10833: dataIn1 = 32'd589
; 
32'd10834: dataIn1 = 32'd596
; 
32'd10835: dataIn1 = 32'd611
; 
32'd10836: dataIn1 = 32'd613
; 
32'd10837: dataIn1 = 32'd614
; 
32'd10838: dataIn1 = 32'd617
; 
32'd10839: dataIn1 = 32'd627
; 
32'd10840: dataIn1 = 32'd633
; 
32'd10841: dataIn1 = 32'd635
; 
32'd10842: dataIn1 = 32'd650
; 
32'd10843: dataIn1 = 32'd662
; 
32'd10844: dataIn1 = 32'd671
; 
32'd10845: dataIn1 = 32'd674
; 
32'd10846: dataIn1 = 32'd687
; 
32'd10847: dataIn1 = 32'd701
; 
32'd10848: dataIn1 = 32'd702
; 
32'd10849: dataIn1 = 32'd724
; 
32'd10850: dataIn1 = 32'd736
; 
32'd10851: dataIn1 = 32'd740
; 
32'd10852: dataIn1 = 32'd744
; 
32'd10853: dataIn1 = 32'd750
; 
32'd10854: dataIn1 = 32'd784
; 
32'd10855: dataIn1 = 32'd82
; 
32'd10856: dataIn1 = 32'd88
; 
32'd10857: dataIn1 = 32'd93
; 
32'd10858: dataIn1 = 32'd112
; 
32'd10859: dataIn1 = 32'd182
; 
32'd10860: dataIn1 = 32'd208
; 
32'd10861: dataIn1 = 32'd229
; 
32'd10862: dataIn1 = 32'd240
; 
32'd10863: dataIn1 = 32'd258
; 
32'd10864: dataIn1 = 32'd263
; 
32'd10865: dataIn1 = 32'd281
; 
32'd10866: dataIn1 = 32'd289
; 
32'd10867: dataIn1 = 32'd304
; 
32'd10868: dataIn1 = 32'd320
; 
32'd10869: dataIn1 = 32'd326
; 
32'd10870: dataIn1 = 32'd328
; 
32'd10871: dataIn1 = 32'd331
; 
32'd10872: dataIn1 = 32'd337
; 
32'd10873: dataIn1 = 32'd364
; 
32'd10874: dataIn1 = 32'd368
; 
32'd10875: dataIn1 = 32'd382
; 
32'd10876: dataIn1 = 32'd390
; 
32'd10877: dataIn1 = 32'd396
; 
32'd10878: dataIn1 = 32'd400
; 
32'd10879: dataIn1 = 32'd419
; 
32'd10880: dataIn1 = 32'd446
; 
32'd10881: dataIn1 = 32'd467
; 
32'd10882: dataIn1 = 32'd474
; 
32'd10883: dataIn1 = 32'd501
; 
32'd10884: dataIn1 = 32'd509
; 
32'd10885: dataIn1 = 32'd530
; 
32'd10886: dataIn1 = 32'd571
; 
32'd10887: dataIn1 = 32'd581
; 
32'd10888: dataIn1 = 32'd592
; 
32'd10889: dataIn1 = 32'd629
; 
32'd10890: dataIn1 = 32'd646
; 
32'd10891: dataIn1 = 32'd669
; 
32'd10892: dataIn1 = 32'd671
; 
32'd10893: dataIn1 = 32'd684
; 
32'd10894: dataIn1 = 32'd701
; 
32'd10895: dataIn1 = 32'd738
; 
32'd10896: dataIn1 = 32'd775
; 
32'd10897: dataIn1 = 32'd779
; 
32'd10898: dataIn1 = 32'd72
; 
32'd10899: dataIn1 = 32'd77
; 
32'd10900: dataIn1 = 32'd79
; 
32'd10901: dataIn1 = 32'd84
; 
32'd10902: dataIn1 = 32'd102
; 
32'd10903: dataIn1 = 32'd147
; 
32'd10904: dataIn1 = 32'd169
; 
32'd10905: dataIn1 = 32'd192
; 
32'd10906: dataIn1 = 32'd194
; 
32'd10907: dataIn1 = 32'd195
; 
32'd10908: dataIn1 = 32'd199
; 
32'd10909: dataIn1 = 32'd212
; 
32'd10910: dataIn1 = 32'd238
; 
32'd10911: dataIn1 = 32'd268
; 
32'd10912: dataIn1 = 32'd290
; 
32'd10913: dataIn1 = 32'd292
; 
32'd10914: dataIn1 = 32'd299
; 
32'd10915: dataIn1 = 32'd307
; 
32'd10916: dataIn1 = 32'd308
; 
32'd10917: dataIn1 = 32'd327
; 
32'd10918: dataIn1 = 32'd364
; 
32'd10919: dataIn1 = 32'd378
; 
32'd10920: dataIn1 = 32'd431
; 
32'd10921: dataIn1 = 32'd437
; 
32'd10922: dataIn1 = 32'd443
; 
32'd10923: dataIn1 = 32'd446
; 
32'd10924: dataIn1 = 32'd455
; 
32'd10925: dataIn1 = 32'd465
; 
32'd10926: dataIn1 = 32'd474
; 
32'd10927: dataIn1 = 32'd479
; 
32'd10928: dataIn1 = 32'd508
; 
32'd10929: dataIn1 = 32'd510
; 
32'd10930: dataIn1 = 32'd523
; 
32'd10931: dataIn1 = 32'd544
; 
32'd10932: dataIn1 = 32'd547
; 
32'd10933: dataIn1 = 32'd553
; 
32'd10934: dataIn1 = 32'd577
; 
32'd10935: dataIn1 = 32'd588
; 
32'd10936: dataIn1 = 32'd597
; 
32'd10937: dataIn1 = 32'd617
; 
32'd10938: dataIn1 = 32'd633
; 
32'd10939: dataIn1 = 32'd644
; 
32'd10940: dataIn1 = 32'd698
; 
32'd10941: dataIn1 = 32'd706
; 
32'd10942: dataIn1 = 32'd729
; 
32'd10943: dataIn1 = 32'd734
; 
32'd10944: dataIn1 = 32'd768
; 
32'd10945: dataIn1 = 32'd783
; 
32'd10946: dataIn1 = 32'd786
; 
32'd10947: dataIn1 = 32'd791
; 
32'd10948: dataIn1 = 32'd799
; 
32'd10949: dataIn1 = 32'd67
; 
32'd10950: dataIn1 = 32'd70
; 
32'd10951: dataIn1 = 32'd75
; 
32'd10952: dataIn1 = 32'd93
; 
32'd10953: dataIn1 = 32'd127
; 
32'd10954: dataIn1 = 32'd141
; 
32'd10955: dataIn1 = 32'd195
; 
32'd10956: dataIn1 = 32'd216
; 
32'd10957: dataIn1 = 32'd239
; 
32'd10958: dataIn1 = 32'd250
; 
32'd10959: dataIn1 = 32'd268
; 
32'd10960: dataIn1 = 32'd278
; 
32'd10961: dataIn1 = 32'd281
; 
32'd10962: dataIn1 = 32'd285
; 
32'd10963: dataIn1 = 32'd309
; 
32'd10964: dataIn1 = 32'd312
; 
32'd10965: dataIn1 = 32'd323
; 
32'd10966: dataIn1 = 32'd382
; 
32'd10967: dataIn1 = 32'd384
; 
32'd10968: dataIn1 = 32'd395
; 
32'd10969: dataIn1 = 32'd414
; 
32'd10970: dataIn1 = 32'd422
; 
32'd10971: dataIn1 = 32'd438
; 
32'd10972: dataIn1 = 32'd440
; 
32'd10973: dataIn1 = 32'd462
; 
32'd10974: dataIn1 = 32'd465
; 
32'd10975: dataIn1 = 32'd519
; 
32'd10976: dataIn1 = 32'd521
; 
32'd10977: dataIn1 = 32'd525
; 
32'd10978: dataIn1 = 32'd536
; 
32'd10979: dataIn1 = 32'd555
; 
32'd10980: dataIn1 = 32'd590
; 
32'd10981: dataIn1 = 32'd601
; 
32'd10982: dataIn1 = 32'd603
; 
32'd10983: dataIn1 = 32'd645
; 
32'd10984: dataIn1 = 32'd656
; 
32'd10985: dataIn1 = 32'd660
; 
32'd10986: dataIn1 = 32'd665
; 
32'd10987: dataIn1 = 32'd687
; 
32'd10988: dataIn1 = 32'd703
; 
32'd10989: dataIn1 = 32'd735
; 
32'd10990: dataIn1 = 32'd760
; 
32'd10991: dataIn1 = 32'd774
; 
32'd10992: dataIn1 = 32'd785
; 
32'd10993: dataIn1 = 32'd797
; 
32'd10994: dataIn1 = 32'd96
; 
32'd10995: dataIn1 = 32'd99
; 
32'd10996: dataIn1 = 32'd109
; 
32'd10997: dataIn1 = 32'd139
; 
32'd10998: dataIn1 = 32'd163
; 
32'd10999: dataIn1 = 32'd171
; 
32'd11000: dataIn1 = 32'd172
; 
32'd11001: dataIn1 = 32'd196
; 
32'd11002: dataIn1 = 32'd198
; 
32'd11003: dataIn1 = 32'd257
; 
32'd11004: dataIn1 = 32'd270
; 
32'd11005: dataIn1 = 32'd284
; 
32'd11006: dataIn1 = 32'd316
; 
32'd11007: dataIn1 = 32'd332
; 
32'd11008: dataIn1 = 32'd359
; 
32'd11009: dataIn1 = 32'd372
; 
32'd11010: dataIn1 = 32'd379
; 
32'd11011: dataIn1 = 32'd389
; 
32'd11012: dataIn1 = 32'd392
; 
32'd11013: dataIn1 = 32'd418
; 
32'd11014: dataIn1 = 32'd429
; 
32'd11015: dataIn1 = 32'd430
; 
32'd11016: dataIn1 = 32'd434
; 
32'd11017: dataIn1 = 32'd441
; 
32'd11018: dataIn1 = 32'd453
; 
32'd11019: dataIn1 = 32'd466
; 
32'd11020: dataIn1 = 32'd473
; 
32'd11021: dataIn1 = 32'd479
; 
32'd11022: dataIn1 = 32'd482
; 
32'd11023: dataIn1 = 32'd507
; 
32'd11024: dataIn1 = 32'd574
; 
32'd11025: dataIn1 = 32'd603
; 
32'd11026: dataIn1 = 32'd621
; 
32'd11027: dataIn1 = 32'd622
; 
32'd11028: dataIn1 = 32'd661
; 
32'd11029: dataIn1 = 32'd693
; 
32'd11030: dataIn1 = 32'd706
; 
32'd11031: dataIn1 = 32'd723
; 
32'd11032: dataIn1 = 32'd725
; 
32'd11033: dataIn1 = 32'd735
; 
32'd11034: dataIn1 = 32'd763
; 
32'd11035: dataIn1 = 32'd779
; 
32'd11036: dataIn1 = 32'd781
; 
32'd11037: dataIn1 = 32'd69
; 
32'd11038: dataIn1 = 32'd124
; 
32'd11039: dataIn1 = 32'd134
; 
32'd11040: dataIn1 = 32'd164
; 
32'd11041: dataIn1 = 32'd182
; 
32'd11042: dataIn1 = 32'd196
; 
32'd11043: dataIn1 = 32'd206
; 
32'd11044: dataIn1 = 32'd222
; 
32'd11045: dataIn1 = 32'd305
; 
32'd11046: dataIn1 = 32'd316
; 
32'd11047: dataIn1 = 32'd329
; 
32'd11048: dataIn1 = 32'd339
; 
32'd11049: dataIn1 = 32'd348
; 
32'd11050: dataIn1 = 32'd396
; 
32'd11051: dataIn1 = 32'd414
; 
32'd11052: dataIn1 = 32'd442
; 
32'd11053: dataIn1 = 32'd444
; 
32'd11054: dataIn1 = 32'd455
; 
32'd11055: dataIn1 = 32'd506
; 
32'd11056: dataIn1 = 32'd519
; 
32'd11057: dataIn1 = 32'd522
; 
32'd11058: dataIn1 = 32'd545
; 
32'd11059: dataIn1 = 32'd628
; 
32'd11060: dataIn1 = 32'd641
; 
32'd11061: dataIn1 = 32'd656
; 
32'd11062: dataIn1 = 32'd658
; 
32'd11063: dataIn1 = 32'd690
; 
32'd11064: dataIn1 = 32'd700
; 
32'd11065: dataIn1 = 32'd739
; 
32'd11066: dataIn1 = 32'd754
; 
32'd11067: dataIn1 = 32'd762
; 
32'd11068: dataIn1 = 32'd789
; 
32'd11069: dataIn1 = 32'd796
; 
32'd11070: dataIn1 = 32'd86
; 
32'd11071: dataIn1 = 32'd88
; 
32'd11072: dataIn1 = 32'd170
; 
32'd11073: dataIn1 = 32'd198
; 
32'd11074: dataIn1 = 32'd213
; 
32'd11075: dataIn1 = 32'd232
; 
32'd11076: dataIn1 = 32'd240
; 
32'd11077: dataIn1 = 32'd259
; 
32'd11078: dataIn1 = 32'd288
; 
32'd11079: dataIn1 = 32'd348
; 
32'd11080: dataIn1 = 32'd367
; 
32'd11081: dataIn1 = 32'd376
; 
32'd11082: dataIn1 = 32'd378
; 
32'd11083: dataIn1 = 32'd379
; 
32'd11084: dataIn1 = 32'd383
; 
32'd11085: dataIn1 = 32'd393
; 
32'd11086: dataIn1 = 32'd406
; 
32'd11087: dataIn1 = 32'd431
; 
32'd11088: dataIn1 = 32'd432
; 
32'd11089: dataIn1 = 32'd445
; 
32'd11090: dataIn1 = 32'd508
; 
32'd11091: dataIn1 = 32'd511
; 
32'd11092: dataIn1 = 32'd518
; 
32'd11093: dataIn1 = 32'd524
; 
32'd11094: dataIn1 = 32'd549
; 
32'd11095: dataIn1 = 32'd555
; 
32'd11096: dataIn1 = 32'd556
; 
32'd11097: dataIn1 = 32'd561
; 
32'd11098: dataIn1 = 32'd594
; 
32'd11099: dataIn1 = 32'd598
; 
32'd11100: dataIn1 = 32'd619
; 
32'd11101: dataIn1 = 32'd625
; 
32'd11102: dataIn1 = 32'd626
; 
32'd11103: dataIn1 = 32'd666
; 
32'd11104: dataIn1 = 32'd680
; 
32'd11105: dataIn1 = 32'd692
; 
32'd11106: dataIn1 = 32'd753
; 
32'd11107: dataIn1 = 32'd761
; 
32'd11108: dataIn1 = 32'd84
; 
32'd11109: dataIn1 = 32'd97
; 
32'd11110: dataIn1 = 32'd104
; 
32'd11111: dataIn1 = 32'd139
; 
32'd11112: dataIn1 = 32'd144
; 
32'd11113: dataIn1 = 32'd161
; 
32'd11114: dataIn1 = 32'd189
; 
32'd11115: dataIn1 = 32'd199
; 
32'd11116: dataIn1 = 32'd200
; 
32'd11117: dataIn1 = 32'd216
; 
32'd11118: dataIn1 = 32'd272
; 
32'd11119: dataIn1 = 32'd326
; 
32'd11120: dataIn1 = 32'd344
; 
32'd11121: dataIn1 = 32'd353
; 
32'd11122: dataIn1 = 32'd355
; 
32'd11123: dataIn1 = 32'd381
; 
32'd11124: dataIn1 = 32'd391
; 
32'd11125: dataIn1 = 32'd401
; 
32'd11126: dataIn1 = 32'd477
; 
32'd11127: dataIn1 = 32'd490
; 
32'd11128: dataIn1 = 32'd491
; 
32'd11129: dataIn1 = 32'd547
; 
32'd11130: dataIn1 = 32'd554
; 
32'd11131: dataIn1 = 32'd561
; 
32'd11132: dataIn1 = 32'd576
; 
32'd11133: dataIn1 = 32'd595
; 
32'd11134: dataIn1 = 32'd601
; 
32'd11135: dataIn1 = 32'd611
; 
32'd11136: dataIn1 = 32'd624
; 
32'd11137: dataIn1 = 32'd643
; 
32'd11138: dataIn1 = 32'd646
; 
32'd11139: dataIn1 = 32'd655
; 
32'd11140: dataIn1 = 32'd699
; 
32'd11141: dataIn1 = 32'd716
; 
32'd11142: dataIn1 = 32'd718
; 
32'd11143: dataIn1 = 32'd719
; 
32'd11144: dataIn1 = 32'd723
; 
32'd11145: dataIn1 = 32'd734
; 
32'd11146: dataIn1 = 32'd748
; 
32'd11147: dataIn1 = 32'd759
; 
32'd11148: dataIn1 = 32'd773
; 
32'd11149: dataIn1 = 32'd78
; 
32'd11150: dataIn1 = 32'd88
; 
32'd11151: dataIn1 = 32'd99
; 
32'd11152: dataIn1 = 32'd103
; 
32'd11153: dataIn1 = 32'd106
; 
32'd11154: dataIn1 = 32'd124
; 
32'd11155: dataIn1 = 32'd164
; 
32'd11156: dataIn1 = 32'd214
; 
32'd11157: dataIn1 = 32'd224
; 
32'd11158: dataIn1 = 32'd226
; 
32'd11159: dataIn1 = 32'd231
; 
32'd11160: dataIn1 = 32'd240
; 
32'd11161: dataIn1 = 32'd243
; 
32'd11162: dataIn1 = 32'd252
; 
32'd11163: dataIn1 = 32'd263
; 
32'd11164: dataIn1 = 32'd328
; 
32'd11165: dataIn1 = 32'd356
; 
32'd11166: dataIn1 = 32'd386
; 
32'd11167: dataIn1 = 32'd388
; 
32'd11168: dataIn1 = 32'd389
; 
32'd11169: dataIn1 = 32'd391
; 
32'd11170: dataIn1 = 32'd419
; 
32'd11171: dataIn1 = 32'd436
; 
32'd11172: dataIn1 = 32'd447
; 
32'd11173: dataIn1 = 32'd464
; 
32'd11174: dataIn1 = 32'd481
; 
32'd11175: dataIn1 = 32'd485
; 
32'd11176: dataIn1 = 32'd494
; 
32'd11177: dataIn1 = 32'd579
; 
32'd11178: dataIn1 = 32'd583
; 
32'd11179: dataIn1 = 32'd586
; 
32'd11180: dataIn1 = 32'd589
; 
32'd11181: dataIn1 = 32'd613
; 
32'd11182: dataIn1 = 32'd619
; 
32'd11183: dataIn1 = 32'd636
; 
32'd11184: dataIn1 = 32'd664
; 
32'd11185: dataIn1 = 32'd739
; 
32'd11186: dataIn1 = 32'd751
; 
32'd11187: dataIn1 = 32'd757
; 
32'd11188: dataIn1 = 32'd776
; 
32'd11189: dataIn1 = 32'd787
; 
32'd11190: dataIn1 = 32'd790
; 
32'd11191: dataIn1 = 32'd792
; 
32'd11192: dataIn1 = 32'd795
; 
32'd11193: dataIn1 = 32'd79
; 
32'd11194: dataIn1 = 32'd83
; 
32'd11195: dataIn1 = 32'd87
; 
32'd11196: dataIn1 = 32'd106
; 
32'd11197: dataIn1 = 32'd109
; 
32'd11198: dataIn1 = 32'd125
; 
32'd11199: dataIn1 = 32'd149
; 
32'd11200: dataIn1 = 32'd159
; 
32'd11201: dataIn1 = 32'd188
; 
32'd11202: dataIn1 = 32'd216
; 
32'd11203: dataIn1 = 32'd225
; 
32'd11204: dataIn1 = 32'd249
; 
32'd11205: dataIn1 = 32'd252
; 
32'd11206: dataIn1 = 32'd266
; 
32'd11207: dataIn1 = 32'd275
; 
32'd11208: dataIn1 = 32'd276
; 
32'd11209: dataIn1 = 32'd296
; 
32'd11210: dataIn1 = 32'd323
; 
32'd11211: dataIn1 = 32'd355
; 
32'd11212: dataIn1 = 32'd364
; 
32'd11213: dataIn1 = 32'd392
; 
32'd11214: dataIn1 = 32'd460
; 
32'd11215: dataIn1 = 32'd463
; 
32'd11216: dataIn1 = 32'd474
; 
32'd11217: dataIn1 = 32'd488
; 
32'd11218: dataIn1 = 32'd492
; 
32'd11219: dataIn1 = 32'd514
; 
32'd11220: dataIn1 = 32'd529
; 
32'd11221: dataIn1 = 32'd532
; 
32'd11222: dataIn1 = 32'd559
; 
32'd11223: dataIn1 = 32'd569
; 
32'd11224: dataIn1 = 32'd602
; 
32'd11225: dataIn1 = 32'd615
; 
32'd11226: dataIn1 = 32'd633
; 
32'd11227: dataIn1 = 32'd648
; 
32'd11228: dataIn1 = 32'd656
; 
32'd11229: dataIn1 = 32'd695
; 
32'd11230: dataIn1 = 32'd715
; 
32'd11231: dataIn1 = 32'd734
; 
32'd11232: dataIn1 = 32'd780
; 
32'd11233: dataIn1 = 32'd784
; 
32'd11234: dataIn1 = 32'd790
; 
32'd11235: dataIn1 = 32'd795
; 
32'd11236: dataIn1 = 32'd96
; 
32'd11237: dataIn1 = 32'd101
; 
32'd11238: dataIn1 = 32'd103
; 
32'd11239: dataIn1 = 32'd104
; 
32'd11240: dataIn1 = 32'd116
; 
32'd11241: dataIn1 = 32'd143
; 
32'd11242: dataIn1 = 32'd148
; 
32'd11243: dataIn1 = 32'd162
; 
32'd11244: dataIn1 = 32'd190
; 
32'd11245: dataIn1 = 32'd191
; 
32'd11246: dataIn1 = 32'd230
; 
32'd11247: dataIn1 = 32'd241
; 
32'd11248: dataIn1 = 32'd245
; 
32'd11249: dataIn1 = 32'd249
; 
32'd11250: dataIn1 = 32'd252
; 
32'd11251: dataIn1 = 32'd266
; 
32'd11252: dataIn1 = 32'd291
; 
32'd11253: dataIn1 = 32'd363
; 
32'd11254: dataIn1 = 32'd364
; 
32'd11255: dataIn1 = 32'd366
; 
32'd11256: dataIn1 = 32'd380
; 
32'd11257: dataIn1 = 32'd419
; 
32'd11258: dataIn1 = 32'd429
; 
32'd11259: dataIn1 = 32'd464
; 
32'd11260: dataIn1 = 32'd477
; 
32'd11261: dataIn1 = 32'd500
; 
32'd11262: dataIn1 = 32'd510
; 
32'd11263: dataIn1 = 32'd625
; 
32'd11264: dataIn1 = 32'd626
; 
32'd11265: dataIn1 = 32'd661
; 
32'd11266: dataIn1 = 32'd675
; 
32'd11267: dataIn1 = 32'd696
; 
32'd11268: dataIn1 = 32'd715
; 
32'd11269: dataIn1 = 32'd777
; 
32'd11270: dataIn1 = 32'd787
; 
32'd11271: dataIn1 = 32'd131
; 
32'd11272: dataIn1 = 32'd142
; 
32'd11273: dataIn1 = 32'd156
; 
32'd11274: dataIn1 = 32'd162
; 
32'd11275: dataIn1 = 32'd207
; 
32'd11276: dataIn1 = 32'd220
; 
32'd11277: dataIn1 = 32'd232
; 
32'd11278: dataIn1 = 32'd234
; 
32'd11279: dataIn1 = 32'd251
; 
32'd11280: dataIn1 = 32'd275
; 
32'd11281: dataIn1 = 32'd291
; 
32'd11282: dataIn1 = 32'd293
; 
32'd11283: dataIn1 = 32'd300
; 
32'd11284: dataIn1 = 32'd339
; 
32'd11285: dataIn1 = 32'd344
; 
32'd11286: dataIn1 = 32'd365
; 
32'd11287: dataIn1 = 32'd369
; 
32'd11288: dataIn1 = 32'd398
; 
32'd11289: dataIn1 = 32'd428
; 
32'd11290: dataIn1 = 32'd441
; 
32'd11291: dataIn1 = 32'd447
; 
32'd11292: dataIn1 = 32'd463
; 
32'd11293: dataIn1 = 32'd475
; 
32'd11294: dataIn1 = 32'd504
; 
32'd11295: dataIn1 = 32'd514
; 
32'd11296: dataIn1 = 32'd529
; 
32'd11297: dataIn1 = 32'd553
; 
32'd11298: dataIn1 = 32'd557
; 
32'd11299: dataIn1 = 32'd566
; 
32'd11300: dataIn1 = 32'd585
; 
32'd11301: dataIn1 = 32'd603
; 
32'd11302: dataIn1 = 32'd625
; 
32'd11303: dataIn1 = 32'd671
; 
32'd11304: dataIn1 = 32'd681
; 
32'd11305: dataIn1 = 32'd725
; 
32'd11306: dataIn1 = 32'd745
; 
32'd11307: dataIn1 = 32'd777
; 
32'd11308: dataIn1 = 32'd782
; 
32'd11309: dataIn1 = 32'd145
; 
32'd11310: dataIn1 = 32'd158
; 
32'd11311: dataIn1 = 32'd164
; 
32'd11312: dataIn1 = 32'd167
; 
32'd11313: dataIn1 = 32'd186
; 
32'd11314: dataIn1 = 32'd191
; 
32'd11315: dataIn1 = 32'd227
; 
32'd11316: dataIn1 = 32'd249
; 
32'd11317: dataIn1 = 32'd259
; 
32'd11318: dataIn1 = 32'd282
; 
32'd11319: dataIn1 = 32'd286
; 
32'd11320: dataIn1 = 32'd336
; 
32'd11321: dataIn1 = 32'd342
; 
32'd11322: dataIn1 = 32'd392
; 
32'd11323: dataIn1 = 32'd428
; 
32'd11324: dataIn1 = 32'd447
; 
32'd11325: dataIn1 = 32'd455
; 
32'd11326: dataIn1 = 32'd492
; 
32'd11327: dataIn1 = 32'd507
; 
32'd11328: dataIn1 = 32'd538
; 
32'd11329: dataIn1 = 32'd571
; 
32'd11330: dataIn1 = 32'd620
; 
32'd11331: dataIn1 = 32'd629
; 
32'd11332: dataIn1 = 32'd632
; 
32'd11333: dataIn1 = 32'd643
; 
32'd11334: dataIn1 = 32'd659
; 
32'd11335: dataIn1 = 32'd697
; 
32'd11336: dataIn1 = 32'd733
; 
32'd11337: dataIn1 = 32'd736
; 
32'd11338: dataIn1 = 32'd787
; 
32'd11339: dataIn1 = 32'd111
; 
32'd11340: dataIn1 = 32'd143
; 
32'd11341: dataIn1 = 32'd150
; 
32'd11342: dataIn1 = 32'd156
; 
32'd11343: dataIn1 = 32'd181
; 
32'd11344: dataIn1 = 32'd206
; 
32'd11345: dataIn1 = 32'd247
; 
32'd11346: dataIn1 = 32'd253
; 
32'd11347: dataIn1 = 32'd262
; 
32'd11348: dataIn1 = 32'd275
; 
32'd11349: dataIn1 = 32'd277
; 
32'd11350: dataIn1 = 32'd286
; 
32'd11351: dataIn1 = 32'd289
; 
32'd11352: dataIn1 = 32'd334
; 
32'd11353: dataIn1 = 32'd383
; 
32'd11354: dataIn1 = 32'd456
; 
32'd11355: dataIn1 = 32'd476
; 
32'd11356: dataIn1 = 32'd538
; 
32'd11357: dataIn1 = 32'd554
; 
32'd11358: dataIn1 = 32'd560
; 
32'd11359: dataIn1 = 32'd567
; 
32'd11360: dataIn1 = 32'd577
; 
32'd11361: dataIn1 = 32'd582
; 
32'd11362: dataIn1 = 32'd584
; 
32'd11363: dataIn1 = 32'd587
; 
32'd11364: dataIn1 = 32'd612
; 
32'd11365: dataIn1 = 32'd625
; 
32'd11366: dataIn1 = 32'd640
; 
32'd11367: dataIn1 = 32'd657
; 
32'd11368: dataIn1 = 32'd703
; 
32'd11369: dataIn1 = 32'd708
; 
32'd11370: dataIn1 = 32'd714
; 
32'd11371: dataIn1 = 32'd719
; 
32'd11372: dataIn1 = 32'd721
; 
32'd11373: dataIn1 = 32'd722
; 
32'd11374: dataIn1 = 32'd724
; 
32'd11375: dataIn1 = 32'd727
; 
32'd11376: dataIn1 = 32'd757
; 
32'd11377: dataIn1 = 32'd790
; 
32'd11378: dataIn1 = 32'd800
; 
32'd11379: dataIn1 = 32'd86
; 
32'd11380: dataIn1 = 32'd110
; 
32'd11381: dataIn1 = 32'd119
; 
32'd11382: dataIn1 = 32'd124
; 
32'd11383: dataIn1 = 32'd178
; 
32'd11384: dataIn1 = 32'd201
; 
32'd11385: dataIn1 = 32'd217
; 
32'd11386: dataIn1 = 32'd222
; 
32'd11387: dataIn1 = 32'd238
; 
32'd11388: dataIn1 = 32'd249
; 
32'd11389: dataIn1 = 32'd255
; 
32'd11390: dataIn1 = 32'd269
; 
32'd11391: dataIn1 = 32'd276
; 
32'd11392: dataIn1 = 32'd286
; 
32'd11393: dataIn1 = 32'd322
; 
32'd11394: dataIn1 = 32'd336
; 
32'd11395: dataIn1 = 32'd351
; 
32'd11396: dataIn1 = 32'd357
; 
32'd11397: dataIn1 = 32'd368
; 
32'd11398: dataIn1 = 32'd376
; 
32'd11399: dataIn1 = 32'd431
; 
32'd11400: dataIn1 = 32'd466
; 
32'd11401: dataIn1 = 32'd473
; 
32'd11402: dataIn1 = 32'd475
; 
32'd11403: dataIn1 = 32'd492
; 
32'd11404: dataIn1 = 32'd502
; 
32'd11405: dataIn1 = 32'd541
; 
32'd11406: dataIn1 = 32'd542
; 
32'd11407: dataIn1 = 32'd546
; 
32'd11408: dataIn1 = 32'd567
; 
32'd11409: dataIn1 = 32'd577
; 
32'd11410: dataIn1 = 32'd580
; 
32'd11411: dataIn1 = 32'd605
; 
32'd11412: dataIn1 = 32'd613
; 
32'd11413: dataIn1 = 32'd615
; 
32'd11414: dataIn1 = 32'd666
; 
32'd11415: dataIn1 = 32'd678
; 
32'd11416: dataIn1 = 32'd686
; 
32'd11417: dataIn1 = 32'd690
; 
32'd11418: dataIn1 = 32'd693
; 
32'd11419: dataIn1 = 32'd719
; 
32'd11420: dataIn1 = 32'd741
; 
32'd11421: dataIn1 = 32'd744
; 
32'd11422: dataIn1 = 32'd751
; 
32'd11423: dataIn1 = 32'd755
; 
32'd11424: dataIn1 = 32'd762
; 
32'd11425: dataIn1 = 32'd794
; 
32'd11426: dataIn1 = 32'd98
; 
32'd11427: dataIn1 = 32'd100
; 
32'd11428: dataIn1 = 32'd125
; 
32'd11429: dataIn1 = 32'd130
; 
32'd11430: dataIn1 = 32'd135
; 
32'd11431: dataIn1 = 32'd144
; 
32'd11432: dataIn1 = 32'd147
; 
32'd11433: dataIn1 = 32'd154
; 
32'd11434: dataIn1 = 32'd197
; 
32'd11435: dataIn1 = 32'd230
; 
32'd11436: dataIn1 = 32'd232
; 
32'd11437: dataIn1 = 32'd233
; 
32'd11438: dataIn1 = 32'd240
; 
32'd11439: dataIn1 = 32'd263
; 
32'd11440: dataIn1 = 32'd279
; 
32'd11441: dataIn1 = 32'd307
; 
32'd11442: dataIn1 = 32'd320
; 
32'd11443: dataIn1 = 32'd397
; 
32'd11444: dataIn1 = 32'd403
; 
32'd11445: dataIn1 = 32'd404
; 
32'd11446: dataIn1 = 32'd405
; 
32'd11447: dataIn1 = 32'd406
; 
32'd11448: dataIn1 = 32'd425
; 
32'd11449: dataIn1 = 32'd433
; 
32'd11450: dataIn1 = 32'd465
; 
32'd11451: dataIn1 = 32'd477
; 
32'd11452: dataIn1 = 32'd478
; 
32'd11453: dataIn1 = 32'd482
; 
32'd11454: dataIn1 = 32'd485
; 
32'd11455: dataIn1 = 32'd522
; 
32'd11456: dataIn1 = 32'd561
; 
32'd11457: dataIn1 = 32'd564
; 
32'd11458: dataIn1 = 32'd583
; 
32'd11459: dataIn1 = 32'd585
; 
32'd11460: dataIn1 = 32'd587
; 
32'd11461: dataIn1 = 32'd591
; 
32'd11462: dataIn1 = 32'd595
; 
32'd11463: dataIn1 = 32'd599
; 
32'd11464: dataIn1 = 32'd626
; 
32'd11465: dataIn1 = 32'd646
; 
32'd11466: dataIn1 = 32'd664
; 
32'd11467: dataIn1 = 32'd672
; 
32'd11468: dataIn1 = 32'd682
; 
32'd11469: dataIn1 = 32'd785
; 
32'd11470: dataIn1 = 32'd80
; 
32'd11471: dataIn1 = 32'd119
; 
32'd11472: dataIn1 = 32'd135
; 
32'd11473: dataIn1 = 32'd146
; 
32'd11474: dataIn1 = 32'd170
; 
32'd11475: dataIn1 = 32'd174
; 
32'd11476: dataIn1 = 32'd177
; 
32'd11477: dataIn1 = 32'd208
; 
32'd11478: dataIn1 = 32'd210
; 
32'd11479: dataIn1 = 32'd211
; 
32'd11480: dataIn1 = 32'd217
; 
32'd11481: dataIn1 = 32'd232
; 
32'd11482: dataIn1 = 32'd281
; 
32'd11483: dataIn1 = 32'd282
; 
32'd11484: dataIn1 = 32'd294
; 
32'd11485: dataIn1 = 32'd295
; 
32'd11486: dataIn1 = 32'd334
; 
32'd11487: dataIn1 = 32'd354
; 
32'd11488: dataIn1 = 32'd368
; 
32'd11489: dataIn1 = 32'd376
; 
32'd11490: dataIn1 = 32'd381
; 
32'd11491: dataIn1 = 32'd389
; 
32'd11492: dataIn1 = 32'd390
; 
32'd11493: dataIn1 = 32'd394
; 
32'd11494: dataIn1 = 32'd395
; 
32'd11495: dataIn1 = 32'd410
; 
32'd11496: dataIn1 = 32'd411
; 
32'd11497: dataIn1 = 32'd493
; 
32'd11498: dataIn1 = 32'd506
; 
32'd11499: dataIn1 = 32'd529
; 
32'd11500: dataIn1 = 32'd546
; 
32'd11501: dataIn1 = 32'd556
; 
32'd11502: dataIn1 = 32'd590
; 
32'd11503: dataIn1 = 32'd606
; 
32'd11504: dataIn1 = 32'd621
; 
32'd11505: dataIn1 = 32'd632
; 
32'd11506: dataIn1 = 32'd646
; 
32'd11507: dataIn1 = 32'd671
; 
32'd11508: dataIn1 = 32'd681
; 
32'd11509: dataIn1 = 32'd696
; 
32'd11510: dataIn1 = 32'd703
; 
32'd11511: dataIn1 = 32'd734
; 
32'd11512: dataIn1 = 32'd766
; 
32'd11513: dataIn1 = 32'd85
; 
32'd11514: dataIn1 = 32'd98
; 
32'd11515: dataIn1 = 32'd125
; 
32'd11516: dataIn1 = 32'd126
; 
32'd11517: dataIn1 = 32'd145
; 
32'd11518: dataIn1 = 32'd166
; 
32'd11519: dataIn1 = 32'd178
; 
32'd11520: dataIn1 = 32'd238
; 
32'd11521: dataIn1 = 32'd259
; 
32'd11522: dataIn1 = 32'd260
; 
32'd11523: dataIn1 = 32'd284
; 
32'd11524: dataIn1 = 32'd311
; 
32'd11525: dataIn1 = 32'd343
; 
32'd11526: dataIn1 = 32'd362
; 
32'd11527: dataIn1 = 32'd365
; 
32'd11528: dataIn1 = 32'd421
; 
32'd11529: dataIn1 = 32'd433
; 
32'd11530: dataIn1 = 32'd449
; 
32'd11531: dataIn1 = 32'd569
; 
32'd11532: dataIn1 = 32'd576
; 
32'd11533: dataIn1 = 32'd588
; 
32'd11534: dataIn1 = 32'd598
; 
32'd11535: dataIn1 = 32'd629
; 
32'd11536: dataIn1 = 32'd667
; 
32'd11537: dataIn1 = 32'd670
; 
32'd11538: dataIn1 = 32'd673
; 
32'd11539: dataIn1 = 32'd694
; 
32'd11540: dataIn1 = 32'd700
; 
32'd11541: dataIn1 = 32'd707
; 
32'd11542: dataIn1 = 32'd734
; 
32'd11543: dataIn1 = 32'd747
; 
32'd11544: dataIn1 = 32'd759
; 
32'd11545: dataIn1 = 32'd770
; 
32'd11546: dataIn1 = 32'd778
; 
32'd11547: dataIn1 = 32'd783
; 
32'd11548: dataIn1 = 32'd82
; 
32'd11549: dataIn1 = 32'd100
; 
32'd11550: dataIn1 = 32'd108
; 
32'd11551: dataIn1 = 32'd115
; 
32'd11552: dataIn1 = 32'd121
; 
32'd11553: dataIn1 = 32'd122
; 
32'd11554: dataIn1 = 32'd126
; 
32'd11555: dataIn1 = 32'd148
; 
32'd11556: dataIn1 = 32'd159
; 
32'd11557: dataIn1 = 32'd190
; 
32'd11558: dataIn1 = 32'd193
; 
32'd11559: dataIn1 = 32'd198
; 
32'd11560: dataIn1 = 32'd202
; 
32'd11561: dataIn1 = 32'd210
; 
32'd11562: dataIn1 = 32'd212
; 
32'd11563: dataIn1 = 32'd232
; 
32'd11564: dataIn1 = 32'd239
; 
32'd11565: dataIn1 = 32'd248
; 
32'd11566: dataIn1 = 32'd262
; 
32'd11567: dataIn1 = 32'd273
; 
32'd11568: dataIn1 = 32'd278
; 
32'd11569: dataIn1 = 32'd285
; 
32'd11570: dataIn1 = 32'd293
; 
32'd11571: dataIn1 = 32'd301
; 
32'd11572: dataIn1 = 32'd306
; 
32'd11573: dataIn1 = 32'd322
; 
32'd11574: dataIn1 = 32'd344
; 
32'd11575: dataIn1 = 32'd346
; 
32'd11576: dataIn1 = 32'd365
; 
32'd11577: dataIn1 = 32'd369
; 
32'd11578: dataIn1 = 32'd377
; 
32'd11579: dataIn1 = 32'd378
; 
32'd11580: dataIn1 = 32'd385
; 
32'd11581: dataIn1 = 32'd394
; 
32'd11582: dataIn1 = 32'd396
; 
32'd11583: dataIn1 = 32'd401
; 
32'd11584: dataIn1 = 32'd434
; 
32'd11585: dataIn1 = 32'd452
; 
32'd11586: dataIn1 = 32'd481
; 
32'd11587: dataIn1 = 32'd483
; 
32'd11588: dataIn1 = 32'd528
; 
32'd11589: dataIn1 = 32'd531
; 
32'd11590: dataIn1 = 32'd543
; 
32'd11591: dataIn1 = 32'd569
; 
32'd11592: dataIn1 = 32'd588
; 
32'd11593: dataIn1 = 32'd604
; 
32'd11594: dataIn1 = 32'd627
; 
32'd11595: dataIn1 = 32'd632
; 
32'd11596: dataIn1 = 32'd646
; 
32'd11597: dataIn1 = 32'd660
; 
32'd11598: dataIn1 = 32'd679
; 
32'd11599: dataIn1 = 32'd691
; 
32'd11600: dataIn1 = 32'd692
; 
32'd11601: dataIn1 = 32'd709
; 
32'd11602: dataIn1 = 32'd711
; 
32'd11603: dataIn1 = 32'd740
; 
32'd11604: dataIn1 = 32'd753
; 
32'd11605: dataIn1 = 32'd770
; 
32'd11606: dataIn1 = 32'd776
; 
32'd11607: dataIn1 = 32'd796
; 
32'd11608: dataIn1 = 32'd100
; 
32'd11609: dataIn1 = 32'd118
; 
32'd11610: dataIn1 = 32'd119
; 
32'd11611: dataIn1 = 32'd132
; 
32'd11612: dataIn1 = 32'd154
; 
32'd11613: dataIn1 = 32'd163
; 
32'd11614: dataIn1 = 32'd171
; 
32'd11615: dataIn1 = 32'd204
; 
32'd11616: dataIn1 = 32'd215
; 
32'd11617: dataIn1 = 32'd231
; 
32'd11618: dataIn1 = 32'd233
; 
32'd11619: dataIn1 = 32'd242
; 
32'd11620: dataIn1 = 32'd250
; 
32'd11621: dataIn1 = 32'd287
; 
32'd11622: dataIn1 = 32'd298
; 
32'd11623: dataIn1 = 32'd301
; 
32'd11624: dataIn1 = 32'd317
; 
32'd11625: dataIn1 = 32'd319
; 
32'd11626: dataIn1 = 32'd333
; 
32'd11627: dataIn1 = 32'd359
; 
32'd11628: dataIn1 = 32'd379
; 
32'd11629: dataIn1 = 32'd390
; 
32'd11630: dataIn1 = 32'd393
; 
32'd11631: dataIn1 = 32'd414
; 
32'd11632: dataIn1 = 32'd444
; 
32'd11633: dataIn1 = 32'd472
; 
32'd11634: dataIn1 = 32'd480
; 
32'd11635: dataIn1 = 32'd486
; 
32'd11636: dataIn1 = 32'd499
; 
32'd11637: dataIn1 = 32'd506
; 
32'd11638: dataIn1 = 32'd563
; 
32'd11639: dataIn1 = 32'd567
; 
32'd11640: dataIn1 = 32'd573
; 
32'd11641: dataIn1 = 32'd610
; 
32'd11642: dataIn1 = 32'd619
; 
32'd11643: dataIn1 = 32'd636
; 
32'd11644: dataIn1 = 32'd646
; 
32'd11645: dataIn1 = 32'd649
; 
32'd11646: dataIn1 = 32'd659
; 
32'd11647: dataIn1 = 32'd675
; 
32'd11648: dataIn1 = 32'd682
; 
32'd11649: dataIn1 = 32'd708
; 
32'd11650: dataIn1 = 32'd728
; 
32'd11651: dataIn1 = 32'd730
; 
32'd11652: dataIn1 = 32'd755
; 
32'd11653: dataIn1 = 32'd758
; 
32'd11654: dataIn1 = 32'd764
; 
32'd11655: dataIn1 = 32'd776
; 
32'd11656: dataIn1 = 32'd99
; 
32'd11657: dataIn1 = 32'd105
; 
32'd11658: dataIn1 = 32'd119
; 
32'd11659: dataIn1 = 32'd120
; 
32'd11660: dataIn1 = 32'd124
; 
32'd11661: dataIn1 = 32'd131
; 
32'd11662: dataIn1 = 32'd177
; 
32'd11663: dataIn1 = 32'd193
; 
32'd11664: dataIn1 = 32'd211
; 
32'd11665: dataIn1 = 32'd246
; 
32'd11666: dataIn1 = 32'd286
; 
32'd11667: dataIn1 = 32'd300
; 
32'd11668: dataIn1 = 32'd343
; 
32'd11669: dataIn1 = 32'd391
; 
32'd11670: dataIn1 = 32'd396
; 
32'd11671: dataIn1 = 32'd422
; 
32'd11672: dataIn1 = 32'd425
; 
32'd11673: dataIn1 = 32'd487
; 
32'd11674: dataIn1 = 32'd493
; 
32'd11675: dataIn1 = 32'd498
; 
32'd11676: dataIn1 = 32'd514
; 
32'd11677: dataIn1 = 32'd521
; 
32'd11678: dataIn1 = 32'd530
; 
32'd11679: dataIn1 = 32'd532
; 
32'd11680: dataIn1 = 32'd541
; 
32'd11681: dataIn1 = 32'd586
; 
32'd11682: dataIn1 = 32'd610
; 
32'd11683: dataIn1 = 32'd660
; 
32'd11684: dataIn1 = 32'd668
; 
32'd11685: dataIn1 = 32'd669
; 
32'd11686: dataIn1 = 32'd686
; 
32'd11687: dataIn1 = 32'd700
; 
32'd11688: dataIn1 = 32'd713
; 
32'd11689: dataIn1 = 32'd730
; 
32'd11690: dataIn1 = 32'd739
; 
32'd11691: dataIn1 = 32'd747
; 
32'd11692: dataIn1 = 32'd752
; 
32'd11693: dataIn1 = 32'd784
; 
32'd11694: dataIn1 = 32'd785
; 
32'd11695: dataIn1 = 32'd88
; 
32'd11696: dataIn1 = 32'd115
; 
32'd11697: dataIn1 = 32'd155
; 
32'd11698: dataIn1 = 32'd168
; 
32'd11699: dataIn1 = 32'd169
; 
32'd11700: dataIn1 = 32'd171
; 
32'd11701: dataIn1 = 32'd198
; 
32'd11702: dataIn1 = 32'd213
; 
32'd11703: dataIn1 = 32'd214
; 
32'd11704: dataIn1 = 32'd233
; 
32'd11705: dataIn1 = 32'd262
; 
32'd11706: dataIn1 = 32'd264
; 
32'd11707: dataIn1 = 32'd273
; 
32'd11708: dataIn1 = 32'd277
; 
32'd11709: dataIn1 = 32'd297
; 
32'd11710: dataIn1 = 32'd355
; 
32'd11711: dataIn1 = 32'd358
; 
32'd11712: dataIn1 = 32'd359
; 
32'd11713: dataIn1 = 32'd363
; 
32'd11714: dataIn1 = 32'd381
; 
32'd11715: dataIn1 = 32'd405
; 
32'd11716: dataIn1 = 32'd415
; 
32'd11717: dataIn1 = 32'd420
; 
32'd11718: dataIn1 = 32'd454
; 
32'd11719: dataIn1 = 32'd455
; 
32'd11720: dataIn1 = 32'd471
; 
32'd11721: dataIn1 = 32'd472
; 
32'd11722: dataIn1 = 32'd487
; 
32'd11723: dataIn1 = 32'd489
; 
32'd11724: dataIn1 = 32'd503
; 
32'd11725: dataIn1 = 32'd519
; 
32'd11726: dataIn1 = 32'd565
; 
32'd11727: dataIn1 = 32'd569
; 
32'd11728: dataIn1 = 32'd570
; 
32'd11729: dataIn1 = 32'd580
; 
32'd11730: dataIn1 = 32'd627
; 
32'd11731: dataIn1 = 32'd678
; 
32'd11732: dataIn1 = 32'd680
; 
32'd11733: dataIn1 = 32'd703
; 
32'd11734: dataIn1 = 32'd708
; 
32'd11735: dataIn1 = 32'd713
; 
32'd11736: dataIn1 = 32'd716
; 
32'd11737: dataIn1 = 32'd745
; 
32'd11738: dataIn1 = 32'd764
; 
32'd11739: dataIn1 = 32'd778
; 
32'd11740: dataIn1 = 32'd789
; 
32'd11741: dataIn1 = 32'd158
; 
32'd11742: dataIn1 = 32'd179
; 
32'd11743: dataIn1 = 32'd191
; 
32'd11744: dataIn1 = 32'd235
; 
32'd11745: dataIn1 = 32'd247
; 
32'd11746: dataIn1 = 32'd264
; 
32'd11747: dataIn1 = 32'd279
; 
32'd11748: dataIn1 = 32'd293
; 
32'd11749: dataIn1 = 32'd323
; 
32'd11750: dataIn1 = 32'd364
; 
32'd11751: dataIn1 = 32'd367
; 
32'd11752: dataIn1 = 32'd380
; 
32'd11753: dataIn1 = 32'd389
; 
32'd11754: dataIn1 = 32'd408
; 
32'd11755: dataIn1 = 32'd427
; 
32'd11756: dataIn1 = 32'd436
; 
32'd11757: dataIn1 = 32'd456
; 
32'd11758: dataIn1 = 32'd458
; 
32'd11759: dataIn1 = 32'd461
; 
32'd11760: dataIn1 = 32'd480
; 
32'd11761: dataIn1 = 32'd503
; 
32'd11762: dataIn1 = 32'd507
; 
32'd11763: dataIn1 = 32'd509
; 
32'd11764: dataIn1 = 32'd551
; 
32'd11765: dataIn1 = 32'd574
; 
32'd11766: dataIn1 = 32'd624
; 
32'd11767: dataIn1 = 32'd635
; 
32'd11768: dataIn1 = 32'd642
; 
32'd11769: dataIn1 = 32'd673
; 
32'd11770: dataIn1 = 32'd696
; 
32'd11771: dataIn1 = 32'd718
; 
32'd11772: dataIn1 = 32'd730
; 
32'd11773: dataIn1 = 32'd731
; 
32'd11774: dataIn1 = 32'd745
; 
32'd11775: dataIn1 = 32'd749
; 
32'd11776: dataIn1 = 32'd752
; 
32'd11777: dataIn1 = 32'd755
; 
32'd11778: dataIn1 = 32'd100
; 
32'd11779: dataIn1 = 32'd101
; 
32'd11780: dataIn1 = 32'd117
; 
32'd11781: dataIn1 = 32'd145
; 
32'd11782: dataIn1 = 32'd153
; 
32'd11783: dataIn1 = 32'd160
; 
32'd11784: dataIn1 = 32'd170
; 
32'd11785: dataIn1 = 32'd183
; 
32'd11786: dataIn1 = 32'd226
; 
32'd11787: dataIn1 = 32'd254
; 
32'd11788: dataIn1 = 32'd276
; 
32'd11789: dataIn1 = 32'd300
; 
32'd11790: dataIn1 = 32'd308
; 
32'd11791: dataIn1 = 32'd321
; 
32'd11792: dataIn1 = 32'd324
; 
32'd11793: dataIn1 = 32'd333
; 
32'd11794: dataIn1 = 32'd341
; 
32'd11795: dataIn1 = 32'd347
; 
32'd11796: dataIn1 = 32'd349
; 
32'd11797: dataIn1 = 32'd384
; 
32'd11798: dataIn1 = 32'd411
; 
32'd11799: dataIn1 = 32'd424
; 
32'd11800: dataIn1 = 32'd444
; 
32'd11801: dataIn1 = 32'd455
; 
32'd11802: dataIn1 = 32'd496
; 
32'd11803: dataIn1 = 32'd510
; 
32'd11804: dataIn1 = 32'd532
; 
32'd11805: dataIn1 = 32'd593
; 
32'd11806: dataIn1 = 32'd612
; 
32'd11807: dataIn1 = 32'd636
; 
32'd11808: dataIn1 = 32'd640
; 
32'd11809: dataIn1 = 32'd651
; 
32'd11810: dataIn1 = 32'd670
; 
32'd11811: dataIn1 = 32'd712
; 
32'd11812: dataIn1 = 32'd719
; 
32'd11813: dataIn1 = 32'd744
; 
32'd11814: dataIn1 = 32'd793
; 
32'd11815: dataIn1 = 32'd100
; 
32'd11816: dataIn1 = 32'd114
; 
32'd11817: dataIn1 = 32'd167
; 
32'd11818: dataIn1 = 32'd182
; 
32'd11819: dataIn1 = 32'd200
; 
32'd11820: dataIn1 = 32'd245
; 
32'd11821: dataIn1 = 32'd310
; 
32'd11822: dataIn1 = 32'd320
; 
32'd11823: dataIn1 = 32'd356
; 
32'd11824: dataIn1 = 32'd379
; 
32'd11825: dataIn1 = 32'd425
; 
32'd11826: dataIn1 = 32'd451
; 
32'd11827: dataIn1 = 32'd465
; 
32'd11828: dataIn1 = 32'd470
; 
32'd11829: dataIn1 = 32'd487
; 
32'd11830: dataIn1 = 32'd496
; 
32'd11831: dataIn1 = 32'd507
; 
32'd11832: dataIn1 = 32'd557
; 
32'd11833: dataIn1 = 32'd561
; 
32'd11834: dataIn1 = 32'd566
; 
32'd11835: dataIn1 = 32'd620
; 
32'd11836: dataIn1 = 32'd629
; 
32'd11837: dataIn1 = 32'd633
; 
32'd11838: dataIn1 = 32'd636
; 
32'd11839: dataIn1 = 32'd695
; 
32'd11840: dataIn1 = 32'd705
; 
32'd11841: dataIn1 = 32'd735
; 
32'd11842: dataIn1 = 32'd738
; 
32'd11843: dataIn1 = 32'd795
; 
32'd11844: dataIn1 = 32'd799
; 
32'd11845: dataIn1 = 32'd102
; 
32'd11846: dataIn1 = 32'd172
; 
32'd11847: dataIn1 = 32'd179
; 
32'd11848: dataIn1 = 32'd182
; 
32'd11849: dataIn1 = 32'd203
; 
32'd11850: dataIn1 = 32'd205
; 
32'd11851: dataIn1 = 32'd212
; 
32'd11852: dataIn1 = 32'd218
; 
32'd11853: dataIn1 = 32'd229
; 
32'd11854: dataIn1 = 32'd274
; 
32'd11855: dataIn1 = 32'd288
; 
32'd11856: dataIn1 = 32'd301
; 
32'd11857: dataIn1 = 32'd310
; 
32'd11858: dataIn1 = 32'd314
; 
32'd11859: dataIn1 = 32'd316
; 
32'd11860: dataIn1 = 32'd319
; 
32'd11861: dataIn1 = 32'd361
; 
32'd11862: dataIn1 = 32'd377
; 
32'd11863: dataIn1 = 32'd389
; 
32'd11864: dataIn1 = 32'd392
; 
32'd11865: dataIn1 = 32'd402
; 
32'd11866: dataIn1 = 32'd464
; 
32'd11867: dataIn1 = 32'd475
; 
32'd11868: dataIn1 = 32'd529
; 
32'd11869: dataIn1 = 32'd530
; 
32'd11870: dataIn1 = 32'd545
; 
32'd11871: dataIn1 = 32'd562
; 
32'd11872: dataIn1 = 32'd566
; 
32'd11873: dataIn1 = 32'd568
; 
32'd11874: dataIn1 = 32'd571
; 
32'd11875: dataIn1 = 32'd579
; 
32'd11876: dataIn1 = 32'd581
; 
32'd11877: dataIn1 = 32'd604
; 
32'd11878: dataIn1 = 32'd632
; 
32'd11879: dataIn1 = 32'd634
; 
32'd11880: dataIn1 = 32'd636
; 
32'd11881: dataIn1 = 32'd654
; 
32'd11882: dataIn1 = 32'd662
; 
32'd11883: dataIn1 = 32'd669
; 
32'd11884: dataIn1 = 32'd699
; 
32'd11885: dataIn1 = 32'd702
; 
32'd11886: dataIn1 = 32'd707
; 
32'd11887: dataIn1 = 32'd739
; 
32'd11888: dataIn1 = 32'd800
; 
32'd11889: dataIn1 = 32'd103
; 
32'd11890: dataIn1 = 32'd113
; 
32'd11891: dataIn1 = 32'd114
; 
32'd11892: dataIn1 = 32'd124
; 
32'd11893: dataIn1 = 32'd134
; 
32'd11894: dataIn1 = 32'd146
; 
32'd11895: dataIn1 = 32'd148
; 
32'd11896: dataIn1 = 32'd176
; 
32'd11897: dataIn1 = 32'd187
; 
32'd11898: dataIn1 = 32'd204
; 
32'd11899: dataIn1 = 32'd210
; 
32'd11900: dataIn1 = 32'd213
; 
32'd11901: dataIn1 = 32'd231
; 
32'd11902: dataIn1 = 32'd232
; 
32'd11903: dataIn1 = 32'd235
; 
32'd11904: dataIn1 = 32'd236
; 
32'd11905: dataIn1 = 32'd251
; 
32'd11906: dataIn1 = 32'd260
; 
32'd11907: dataIn1 = 32'd268
; 
32'd11908: dataIn1 = 32'd305
; 
32'd11909: dataIn1 = 32'd332
; 
32'd11910: dataIn1 = 32'd339
; 
32'd11911: dataIn1 = 32'd340
; 
32'd11912: dataIn1 = 32'd352
; 
32'd11913: dataIn1 = 32'd354
; 
32'd11914: dataIn1 = 32'd364
; 
32'd11915: dataIn1 = 32'd375
; 
32'd11916: dataIn1 = 32'd392
; 
32'd11917: dataIn1 = 32'd411
; 
32'd11918: dataIn1 = 32'd417
; 
32'd11919: dataIn1 = 32'd438
; 
32'd11920: dataIn1 = 32'd458
; 
32'd11921: dataIn1 = 32'd467
; 
32'd11922: dataIn1 = 32'd496
; 
32'd11923: dataIn1 = 32'd503
; 
32'd11924: dataIn1 = 32'd510
; 
32'd11925: dataIn1 = 32'd552
; 
32'd11926: dataIn1 = 32'd603
; 
32'd11927: dataIn1 = 32'd630
; 
32'd11928: dataIn1 = 32'd634
; 
32'd11929: dataIn1 = 32'd658
; 
32'd11930: dataIn1 = 32'd665
; 
32'd11931: dataIn1 = 32'd679
; 
32'd11932: dataIn1 = 32'd689
; 
32'd11933: dataIn1 = 32'd710
; 
32'd11934: dataIn1 = 32'd734
; 
32'd11935: dataIn1 = 32'd742
; 
32'd11936: dataIn1 = 32'd757
; 
32'd11937: dataIn1 = 32'd771
; 
32'd11938: dataIn1 = 32'd779
; 
32'd11939: dataIn1 = 32'd782
; 
32'd11940: dataIn1 = 32'd785
; 
32'd11941: dataIn1 = 32'd800
; 
32'd11942: dataIn1 = 32'd117
; 
32'd11943: dataIn1 = 32'd127
; 
32'd11944: dataIn1 = 32'd135
; 
32'd11945: dataIn1 = 32'd177
; 
32'd11946: dataIn1 = 32'd195
; 
32'd11947: dataIn1 = 32'd230
; 
32'd11948: dataIn1 = 32'd263
; 
32'd11949: dataIn1 = 32'd276
; 
32'd11950: dataIn1 = 32'd282
; 
32'd11951: dataIn1 = 32'd300
; 
32'd11952: dataIn1 = 32'd318
; 
32'd11953: dataIn1 = 32'd323
; 
32'd11954: dataIn1 = 32'd347
; 
32'd11955: dataIn1 = 32'd356
; 
32'd11956: dataIn1 = 32'd364
; 
32'd11957: dataIn1 = 32'd374
; 
32'd11958: dataIn1 = 32'd397
; 
32'd11959: dataIn1 = 32'd399
; 
32'd11960: dataIn1 = 32'd402
; 
32'd11961: dataIn1 = 32'd431
; 
32'd11962: dataIn1 = 32'd513
; 
32'd11963: dataIn1 = 32'd515
; 
32'd11964: dataIn1 = 32'd531
; 
32'd11965: dataIn1 = 32'd593
; 
32'd11966: dataIn1 = 32'd620
; 
32'd11967: dataIn1 = 32'd624
; 
32'd11968: dataIn1 = 32'd626
; 
32'd11969: dataIn1 = 32'd629
; 
32'd11970: dataIn1 = 32'd645
; 
32'd11971: dataIn1 = 32'd664
; 
32'd11972: dataIn1 = 32'd666
; 
32'd11973: dataIn1 = 32'd675
; 
32'd11974: dataIn1 = 32'd699
; 
32'd11975: dataIn1 = 32'd708
; 
32'd11976: dataIn1 = 32'd711
; 
32'd11977: dataIn1 = 32'd712
; 
32'd11978: dataIn1 = 32'd713
; 
32'd11979: dataIn1 = 32'd715
; 
32'd11980: dataIn1 = 32'd747
; 
32'd11981: dataIn1 = 32'd758
; 
32'd11982: dataIn1 = 32'd132
; 
32'd11983: dataIn1 = 32'd146
; 
32'd11984: dataIn1 = 32'd171
; 
32'd11985: dataIn1 = 32'd174
; 
32'd11986: dataIn1 = 32'd183
; 
32'd11987: dataIn1 = 32'd206
; 
32'd11988: dataIn1 = 32'd207
; 
32'd11989: dataIn1 = 32'd208
; 
32'd11990: dataIn1 = 32'd225
; 
32'd11991: dataIn1 = 32'd232
; 
32'd11992: dataIn1 = 32'd233
; 
32'd11993: dataIn1 = 32'd245
; 
32'd11994: dataIn1 = 32'd246
; 
32'd11995: dataIn1 = 32'd285
; 
32'd11996: dataIn1 = 32'd290
; 
32'd11997: dataIn1 = 32'd293
; 
32'd11998: dataIn1 = 32'd359
; 
32'd11999: dataIn1 = 32'd370
; 
32'd12000: dataIn1 = 32'd412
; 
32'd12001: dataIn1 = 32'd440
; 
32'd12002: dataIn1 = 32'd441
; 
32'd12003: dataIn1 = 32'd454
; 
32'd12004: dataIn1 = 32'd461
; 
32'd12005: dataIn1 = 32'd466
; 
32'd12006: dataIn1 = 32'd479
; 
32'd12007: dataIn1 = 32'd485
; 
32'd12008: dataIn1 = 32'd488
; 
32'd12009: dataIn1 = 32'd494
; 
32'd12010: dataIn1 = 32'd496
; 
32'd12011: dataIn1 = 32'd530
; 
32'd12012: dataIn1 = 32'd550
; 
32'd12013: dataIn1 = 32'd574
; 
32'd12014: dataIn1 = 32'd592
; 
32'd12015: dataIn1 = 32'd628
; 
32'd12016: dataIn1 = 32'd683
; 
32'd12017: dataIn1 = 32'd690
; 
32'd12018: dataIn1 = 32'd723
; 
32'd12019: dataIn1 = 32'd754
; 
32'd12020: dataIn1 = 32'd769
; 
32'd12021: dataIn1 = 32'd775
; 
32'd12022: dataIn1 = 32'd776
; 
32'd12023: dataIn1 = 32'd788
; 
32'd12024: dataIn1 = 32'd790
; 
32'd12025: dataIn1 = 32'd799
; 
32'd12026: dataIn1 = 32'd103
; 
32'd12027: dataIn1 = 32'd120
; 
32'd12028: dataIn1 = 32'd130
; 
32'd12029: dataIn1 = 32'd181
; 
32'd12030: dataIn1 = 32'd203
; 
32'd12031: dataIn1 = 32'd218
; 
32'd12032: dataIn1 = 32'd233
; 
32'd12033: dataIn1 = 32'd245
; 
32'd12034: dataIn1 = 32'd267
; 
32'd12035: dataIn1 = 32'd276
; 
32'd12036: dataIn1 = 32'd283
; 
32'd12037: dataIn1 = 32'd298
; 
32'd12038: dataIn1 = 32'd305
; 
32'd12039: dataIn1 = 32'd310
; 
32'd12040: dataIn1 = 32'd317
; 
32'd12041: dataIn1 = 32'd329
; 
32'd12042: dataIn1 = 32'd339
; 
32'd12043: dataIn1 = 32'd367
; 
32'd12044: dataIn1 = 32'd396
; 
32'd12045: dataIn1 = 32'd399
; 
32'd12046: dataIn1 = 32'd407
; 
32'd12047: dataIn1 = 32'd411
; 
32'd12048: dataIn1 = 32'd438
; 
32'd12049: dataIn1 = 32'd439
; 
32'd12050: dataIn1 = 32'd463
; 
32'd12051: dataIn1 = 32'd469
; 
32'd12052: dataIn1 = 32'd475
; 
32'd12053: dataIn1 = 32'd476
; 
32'd12054: dataIn1 = 32'd485
; 
32'd12055: dataIn1 = 32'd505
; 
32'd12056: dataIn1 = 32'd537
; 
32'd12057: dataIn1 = 32'd539
; 
32'd12058: dataIn1 = 32'd553
; 
32'd12059: dataIn1 = 32'd560
; 
32'd12060: dataIn1 = 32'd576
; 
32'd12061: dataIn1 = 32'd606
; 
32'd12062: dataIn1 = 32'd619
; 
32'd12063: dataIn1 = 32'd635
; 
32'd12064: dataIn1 = 32'd664
; 
32'd12065: dataIn1 = 32'd665
; 
32'd12066: dataIn1 = 32'd686
; 
32'd12067: dataIn1 = 32'd695
; 
32'd12068: dataIn1 = 32'd696
; 
32'd12069: dataIn1 = 32'd705
; 
32'd12070: dataIn1 = 32'd707
; 
32'd12071: dataIn1 = 32'd753
; 
32'd12072: dataIn1 = 32'd775
; 
32'd12073: dataIn1 = 32'd796
; 
32'd12074: dataIn1 = 32'd116
; 
32'd12075: dataIn1 = 32'd168
; 
32'd12076: dataIn1 = 32'd210
; 
32'd12077: dataIn1 = 32'd226
; 
32'd12078: dataIn1 = 32'd249
; 
32'd12079: dataIn1 = 32'd260
; 
32'd12080: dataIn1 = 32'd272
; 
32'd12081: dataIn1 = 32'd279
; 
32'd12082: dataIn1 = 32'd288
; 
32'd12083: dataIn1 = 32'd296
; 
32'd12084: dataIn1 = 32'd302
; 
32'd12085: dataIn1 = 32'd305
; 
32'd12086: dataIn1 = 32'd319
; 
32'd12087: dataIn1 = 32'd336
; 
32'd12088: dataIn1 = 32'd344
; 
32'd12089: dataIn1 = 32'd358
; 
32'd12090: dataIn1 = 32'd382
; 
32'd12091: dataIn1 = 32'd397
; 
32'd12092: dataIn1 = 32'd419
; 
32'd12093: dataIn1 = 32'd420
; 
32'd12094: dataIn1 = 32'd422
; 
32'd12095: dataIn1 = 32'd427
; 
32'd12096: dataIn1 = 32'd487
; 
32'd12097: dataIn1 = 32'd549
; 
32'd12098: dataIn1 = 32'd552
; 
32'd12099: dataIn1 = 32'd554
; 
32'd12100: dataIn1 = 32'd558
; 
32'd12101: dataIn1 = 32'd562
; 
32'd12102: dataIn1 = 32'd583
; 
32'd12103: dataIn1 = 32'd594
; 
32'd12104: dataIn1 = 32'd600
; 
32'd12105: dataIn1 = 32'd616
; 
32'd12106: dataIn1 = 32'd622
; 
32'd12107: dataIn1 = 32'd637
; 
32'd12108: dataIn1 = 32'd647
; 
32'd12109: dataIn1 = 32'd649
; 
32'd12110: dataIn1 = 32'd652
; 
32'd12111: dataIn1 = 32'd667
; 
32'd12112: dataIn1 = 32'd678
; 
32'd12113: dataIn1 = 32'd683
; 
32'd12114: dataIn1 = 32'd692
; 
32'd12115: dataIn1 = 32'd696
; 
32'd12116: dataIn1 = 32'd697
; 
32'd12117: dataIn1 = 32'd708
; 
32'd12118: dataIn1 = 32'd727
; 
32'd12119: dataIn1 = 32'd744
; 
32'd12120: dataIn1 = 32'd748
; 
32'd12121: dataIn1 = 32'd750
; 
32'd12122: dataIn1 = 32'd775
; 
32'd12123: dataIn1 = 32'd110
; 
32'd12124: dataIn1 = 32'd117
; 
32'd12125: dataIn1 = 32'd118
; 
32'd12126: dataIn1 = 32'd140
; 
32'd12127: dataIn1 = 32'd152
; 
32'd12128: dataIn1 = 32'd153
; 
32'd12129: dataIn1 = 32'd155
; 
32'd12130: dataIn1 = 32'd160
; 
32'd12131: dataIn1 = 32'd203
; 
32'd12132: dataIn1 = 32'd221
; 
32'd12133: dataIn1 = 32'd246
; 
32'd12134: dataIn1 = 32'd267
; 
32'd12135: dataIn1 = 32'd269
; 
32'd12136: dataIn1 = 32'd271
; 
32'd12137: dataIn1 = 32'd279
; 
32'd12138: dataIn1 = 32'd310
; 
32'd12139: dataIn1 = 32'd313
; 
32'd12140: dataIn1 = 32'd315
; 
32'd12141: dataIn1 = 32'd363
; 
32'd12142: dataIn1 = 32'd380
; 
32'd12143: dataIn1 = 32'd398
; 
32'd12144: dataIn1 = 32'd428
; 
32'd12145: dataIn1 = 32'd449
; 
32'd12146: dataIn1 = 32'd472
; 
32'd12147: dataIn1 = 32'd475
; 
32'd12148: dataIn1 = 32'd494
; 
32'd12149: dataIn1 = 32'd499
; 
32'd12150: dataIn1 = 32'd512
; 
32'd12151: dataIn1 = 32'd539
; 
32'd12152: dataIn1 = 32'd547
; 
32'd12153: dataIn1 = 32'd552
; 
32'd12154: dataIn1 = 32'd563
; 
32'd12155: dataIn1 = 32'd571
; 
32'd12156: dataIn1 = 32'd572
; 
32'd12157: dataIn1 = 32'd584
; 
32'd12158: dataIn1 = 32'd603
; 
32'd12159: dataIn1 = 32'd636
; 
32'd12160: dataIn1 = 32'd649
; 
32'd12161: dataIn1 = 32'd677
; 
32'd12162: dataIn1 = 32'd681
; 
32'd12163: dataIn1 = 32'd702
; 
32'd12164: dataIn1 = 32'd722
; 
32'd12165: dataIn1 = 32'd764
; 
32'd12166: dataIn1 = 32'd768
; 
32'd12167: dataIn1 = 32'd100
; 
32'd12168: dataIn1 = 32'd129
; 
32'd12169: dataIn1 = 32'd135
; 
32'd12170: dataIn1 = 32'd150
; 
32'd12171: dataIn1 = 32'd164
; 
32'd12172: dataIn1 = 32'd173
; 
32'd12173: dataIn1 = 32'd181
; 
32'd12174: dataIn1 = 32'd189
; 
32'd12175: dataIn1 = 32'd191
; 
32'd12176: dataIn1 = 32'd198
; 
32'd12177: dataIn1 = 32'd218
; 
32'd12178: dataIn1 = 32'd235
; 
32'd12179: dataIn1 = 32'd253
; 
32'd12180: dataIn1 = 32'd268
; 
32'd12181: dataIn1 = 32'd276
; 
32'd12182: dataIn1 = 32'd314
; 
32'd12183: dataIn1 = 32'd320
; 
32'd12184: dataIn1 = 32'd321
; 
32'd12185: dataIn1 = 32'd329
; 
32'd12186: dataIn1 = 32'd364
; 
32'd12187: dataIn1 = 32'd370
; 
32'd12188: dataIn1 = 32'd376
; 
32'd12189: dataIn1 = 32'd379
; 
32'd12190: dataIn1 = 32'd380
; 
32'd12191: dataIn1 = 32'd387
; 
32'd12192: dataIn1 = 32'd398
; 
32'd12193: dataIn1 = 32'd404
; 
32'd12194: dataIn1 = 32'd411
; 
32'd12195: dataIn1 = 32'd421
; 
32'd12196: dataIn1 = 32'd447
; 
32'd12197: dataIn1 = 32'd473
; 
32'd12198: dataIn1 = 32'd474
; 
32'd12199: dataIn1 = 32'd477
; 
32'd12200: dataIn1 = 32'd502
; 
32'd12201: dataIn1 = 32'd522
; 
32'd12202: dataIn1 = 32'd553
; 
32'd12203: dataIn1 = 32'd563
; 
32'd12204: dataIn1 = 32'd568
; 
32'd12205: dataIn1 = 32'd572
; 
32'd12206: dataIn1 = 32'd574
; 
32'd12207: dataIn1 = 32'd589
; 
32'd12208: dataIn1 = 32'd593
; 
32'd12209: dataIn1 = 32'd631
; 
32'd12210: dataIn1 = 32'd633
; 
32'd12211: dataIn1 = 32'd683
; 
32'd12212: dataIn1 = 32'd696
; 
32'd12213: dataIn1 = 32'd700
; 
32'd12214: dataIn1 = 32'd726
; 
32'd12215: dataIn1 = 32'd764
; 
32'd12216: dataIn1 = 32'd779
; 
32'd12217: dataIn1 = 32'd97
; 
32'd12218: dataIn1 = 32'd109
; 
32'd12219: dataIn1 = 32'd126
; 
32'd12220: dataIn1 = 32'd131
; 
32'd12221: dataIn1 = 32'd143
; 
32'd12222: dataIn1 = 32'd166
; 
32'd12223: dataIn1 = 32'd205
; 
32'd12224: dataIn1 = 32'd222
; 
32'd12225: dataIn1 = 32'd234
; 
32'd12226: dataIn1 = 32'd236
; 
32'd12227: dataIn1 = 32'd239
; 
32'd12228: dataIn1 = 32'd241
; 
32'd12229: dataIn1 = 32'd251
; 
32'd12230: dataIn1 = 32'd253
; 
32'd12231: dataIn1 = 32'd260
; 
32'd12232: dataIn1 = 32'd263
; 
32'd12233: dataIn1 = 32'd311
; 
32'd12234: dataIn1 = 32'd339
; 
32'd12235: dataIn1 = 32'd343
; 
32'd12236: dataIn1 = 32'd344
; 
32'd12237: dataIn1 = 32'd348
; 
32'd12238: dataIn1 = 32'd391
; 
32'd12239: dataIn1 = 32'd393
; 
32'd12240: dataIn1 = 32'd398
; 
32'd12241: dataIn1 = 32'd416
; 
32'd12242: dataIn1 = 32'd423
; 
32'd12243: dataIn1 = 32'd446
; 
32'd12244: dataIn1 = 32'd538
; 
32'd12245: dataIn1 = 32'd566
; 
32'd12246: dataIn1 = 32'd582
; 
32'd12247: dataIn1 = 32'd602
; 
32'd12248: dataIn1 = 32'd619
; 
32'd12249: dataIn1 = 32'd628
; 
32'd12250: dataIn1 = 32'd655
; 
32'd12251: dataIn1 = 32'd686
; 
32'd12252: dataIn1 = 32'd762
; 
32'd12253: dataIn1 = 32'd105
; 
32'd12254: dataIn1 = 32'd107
; 
32'd12255: dataIn1 = 32'd109
; 
32'd12256: dataIn1 = 32'd121
; 
32'd12257: dataIn1 = 32'd130
; 
32'd12258: dataIn1 = 32'd136
; 
32'd12259: dataIn1 = 32'd144
; 
32'd12260: dataIn1 = 32'd170
; 
32'd12261: dataIn1 = 32'd175
; 
32'd12262: dataIn1 = 32'd190
; 
32'd12263: dataIn1 = 32'd198
; 
32'd12264: dataIn1 = 32'd200
; 
32'd12265: dataIn1 = 32'd232
; 
32'd12266: dataIn1 = 32'd236
; 
32'd12267: dataIn1 = 32'd289
; 
32'd12268: dataIn1 = 32'd306
; 
32'd12269: dataIn1 = 32'd313
; 
32'd12270: dataIn1 = 32'd316
; 
32'd12271: dataIn1 = 32'd352
; 
32'd12272: dataIn1 = 32'd357
; 
32'd12273: dataIn1 = 32'd359
; 
32'd12274: dataIn1 = 32'd360
; 
32'd12275: dataIn1 = 32'd369
; 
32'd12276: dataIn1 = 32'd389
; 
32'd12277: dataIn1 = 32'd391
; 
32'd12278: dataIn1 = 32'd395
; 
32'd12279: dataIn1 = 32'd444
; 
32'd12280: dataIn1 = 32'd450
; 
32'd12281: dataIn1 = 32'd461
; 
32'd12282: dataIn1 = 32'd500
; 
32'd12283: dataIn1 = 32'd510
; 
32'd12284: dataIn1 = 32'd520
; 
32'd12285: dataIn1 = 32'd529
; 
32'd12286: dataIn1 = 32'd540
; 
32'd12287: dataIn1 = 32'd547
; 
32'd12288: dataIn1 = 32'd582
; 
32'd12289: dataIn1 = 32'd585
; 
32'd12290: dataIn1 = 32'd586
; 
32'd12291: dataIn1 = 32'd587
; 
32'd12292: dataIn1 = 32'd595
; 
32'd12293: dataIn1 = 32'd631
; 
32'd12294: dataIn1 = 32'd634
; 
32'd12295: dataIn1 = 32'd644
; 
32'd12296: dataIn1 = 32'd646
; 
32'd12297: dataIn1 = 32'd651
; 
32'd12298: dataIn1 = 32'd664
; 
32'd12299: dataIn1 = 32'd683
; 
32'd12300: dataIn1 = 32'd699
; 
32'd12301: dataIn1 = 32'd705
; 
32'd12302: dataIn1 = 32'd713
; 
32'd12303: dataIn1 = 32'd716
; 
32'd12304: dataIn1 = 32'd749
; 
32'd12305: dataIn1 = 32'd752
; 
32'd12306: dataIn1 = 32'd753
; 
32'd12307: dataIn1 = 32'd754
; 
32'd12308: dataIn1 = 32'd765
; 
32'd12309: dataIn1 = 32'd767
; 
32'd12310: dataIn1 = 32'd770
; 
32'd12311: dataIn1 = 32'd771
; 
32'd12312: dataIn1 = 32'd782
; 
32'd12313: dataIn1 = 32'd783
; 
32'd12314: dataIn1 = 32'd793
; 
32'd12315: dataIn1 = 32'd106
; 
32'd12316: dataIn1 = 32'd115
; 
32'd12317: dataIn1 = 32'd122
; 
32'd12318: dataIn1 = 32'd201
; 
32'd12319: dataIn1 = 32'd203
; 
32'd12320: dataIn1 = 32'd211
; 
32'd12321: dataIn1 = 32'd236
; 
32'd12322: dataIn1 = 32'd249
; 
32'd12323: dataIn1 = 32'd256
; 
32'd12324: dataIn1 = 32'd310
; 
32'd12325: dataIn1 = 32'd311
; 
32'd12326: dataIn1 = 32'd326
; 
32'd12327: dataIn1 = 32'd329
; 
32'd12328: dataIn1 = 32'd343
; 
32'd12329: dataIn1 = 32'd355
; 
32'd12330: dataIn1 = 32'd362
; 
32'd12331: dataIn1 = 32'd380
; 
32'd12332: dataIn1 = 32'd416
; 
32'd12333: dataIn1 = 32'd479
; 
32'd12334: dataIn1 = 32'd483
; 
32'd12335: dataIn1 = 32'd486
; 
32'd12336: dataIn1 = 32'd496
; 
32'd12337: dataIn1 = 32'd497
; 
32'd12338: dataIn1 = 32'd498
; 
32'd12339: dataIn1 = 32'd525
; 
32'd12340: dataIn1 = 32'd534
; 
32'd12341: dataIn1 = 32'd550
; 
32'd12342: dataIn1 = 32'd556
; 
32'd12343: dataIn1 = 32'd575
; 
32'd12344: dataIn1 = 32'd576
; 
32'd12345: dataIn1 = 32'd614
; 
32'd12346: dataIn1 = 32'd632
; 
32'd12347: dataIn1 = 32'd633
; 
32'd12348: dataIn1 = 32'd647
; 
32'd12349: dataIn1 = 32'd648
; 
32'd12350: dataIn1 = 32'd663
; 
32'd12351: dataIn1 = 32'd666
; 
32'd12352: dataIn1 = 32'd672
; 
32'd12353: dataIn1 = 32'd693
; 
32'd12354: dataIn1 = 32'd726
; 
32'd12355: dataIn1 = 32'd740
; 
32'd12356: dataIn1 = 32'd743
; 
32'd12357: dataIn1 = 32'd759
; 
32'd12358: dataIn1 = 32'd774
; 
32'd12359: dataIn1 = 32'd781
; 
32'd12360: dataIn1 = 32'd115
; 
32'd12361: dataIn1 = 32'd124
; 
32'd12362: dataIn1 = 32'd126
; 
32'd12363: dataIn1 = 32'd145
; 
32'd12364: dataIn1 = 32'd148
; 
32'd12365: dataIn1 = 32'd168
; 
32'd12366: dataIn1 = 32'd173
; 
32'd12367: dataIn1 = 32'd183
; 
32'd12368: dataIn1 = 32'd184
; 
32'd12369: dataIn1 = 32'd221
; 
32'd12370: dataIn1 = 32'd236
; 
32'd12371: dataIn1 = 32'd263
; 
32'd12372: dataIn1 = 32'd274
; 
32'd12373: dataIn1 = 32'd304
; 
32'd12374: dataIn1 = 32'd325
; 
32'd12375: dataIn1 = 32'd348
; 
32'd12376: dataIn1 = 32'd366
; 
32'd12377: dataIn1 = 32'd367
; 
32'd12378: dataIn1 = 32'd412
; 
32'd12379: dataIn1 = 32'd433
; 
32'd12380: dataIn1 = 32'd446
; 
32'd12381: dataIn1 = 32'd468
; 
32'd12382: dataIn1 = 32'd525
; 
32'd12383: dataIn1 = 32'd546
; 
32'd12384: dataIn1 = 32'd548
; 
32'd12385: dataIn1 = 32'd559
; 
32'd12386: dataIn1 = 32'd561
; 
32'd12387: dataIn1 = 32'd564
; 
32'd12388: dataIn1 = 32'd566
; 
32'd12389: dataIn1 = 32'd571
; 
32'd12390: dataIn1 = 32'd583
; 
32'd12391: dataIn1 = 32'd585
; 
32'd12392: dataIn1 = 32'd590
; 
32'd12393: dataIn1 = 32'd604
; 
32'd12394: dataIn1 = 32'd608
; 
32'd12395: dataIn1 = 32'd612
; 
32'd12396: dataIn1 = 32'd616
; 
32'd12397: dataIn1 = 32'd650
; 
32'd12398: dataIn1 = 32'd658
; 
32'd12399: dataIn1 = 32'd670
; 
32'd12400: dataIn1 = 32'd683
; 
32'd12401: dataIn1 = 32'd688
; 
32'd12402: dataIn1 = 32'd718
; 
32'd12403: dataIn1 = 32'd737
; 
32'd12404: dataIn1 = 32'd760
; 
32'd12405: dataIn1 = 32'd797
; 
32'd12406: dataIn1 = 32'd798
; 
32'd12407: dataIn1 = 32'd116
; 
32'd12408: dataIn1 = 32'd151
; 
32'd12409: dataIn1 = 32'd157
; 
32'd12410: dataIn1 = 32'd167
; 
32'd12411: dataIn1 = 32'd219
; 
32'd12412: dataIn1 = 32'd256
; 
32'd12413: dataIn1 = 32'd259
; 
32'd12414: dataIn1 = 32'd262
; 
32'd12415: dataIn1 = 32'd288
; 
32'd12416: dataIn1 = 32'd289
; 
32'd12417: dataIn1 = 32'd309
; 
32'd12418: dataIn1 = 32'd314
; 
32'd12419: dataIn1 = 32'd333
; 
32'd12420: dataIn1 = 32'd337
; 
32'd12421: dataIn1 = 32'd344
; 
32'd12422: dataIn1 = 32'd363
; 
32'd12423: dataIn1 = 32'd383
; 
32'd12424: dataIn1 = 32'd397
; 
32'd12425: dataIn1 = 32'd405
; 
32'd12426: dataIn1 = 32'd433
; 
32'd12427: dataIn1 = 32'd434
; 
32'd12428: dataIn1 = 32'd449
; 
32'd12429: dataIn1 = 32'd469
; 
32'd12430: dataIn1 = 32'd472
; 
32'd12431: dataIn1 = 32'd479
; 
32'd12432: dataIn1 = 32'd485
; 
32'd12433: dataIn1 = 32'd487
; 
32'd12434: dataIn1 = 32'd504
; 
32'd12435: dataIn1 = 32'd520
; 
32'd12436: dataIn1 = 32'd521
; 
32'd12437: dataIn1 = 32'd522
; 
32'd12438: dataIn1 = 32'd548
; 
32'd12439: dataIn1 = 32'd558
; 
32'd12440: dataIn1 = 32'd586
; 
32'd12441: dataIn1 = 32'd605
; 
32'd12442: dataIn1 = 32'd622
; 
32'd12443: dataIn1 = 32'd666
; 
32'd12444: dataIn1 = 32'd691
; 
32'd12445: dataIn1 = 32'd696
; 
32'd12446: dataIn1 = 32'd715
; 
32'd12447: dataIn1 = 32'd719
; 
32'd12448: dataIn1 = 32'd764
; 
32'd12449: dataIn1 = 32'd766
; 
32'd12450: dataIn1 = 32'd770
; 
32'd12451: dataIn1 = 32'd774
; 
32'd12452: dataIn1 = 32'd791
; 
32'd12453: dataIn1 = 32'd123
; 
32'd12454: dataIn1 = 32'd142
; 
32'd12455: dataIn1 = 32'd147
; 
32'd12456: dataIn1 = 32'd171
; 
32'd12457: dataIn1 = 32'd173
; 
32'd12458: dataIn1 = 32'd186
; 
32'd12459: dataIn1 = 32'd192
; 
32'd12460: dataIn1 = 32'd203
; 
32'd12461: dataIn1 = 32'd204
; 
32'd12462: dataIn1 = 32'd208
; 
32'd12463: dataIn1 = 32'd217
; 
32'd12464: dataIn1 = 32'd232
; 
32'd12465: dataIn1 = 32'd248
; 
32'd12466: dataIn1 = 32'd258
; 
32'd12467: dataIn1 = 32'd273
; 
32'd12468: dataIn1 = 32'd298
; 
32'd12469: dataIn1 = 32'd304
; 
32'd12470: dataIn1 = 32'd305
; 
32'd12471: dataIn1 = 32'd331
; 
32'd12472: dataIn1 = 32'd363
; 
32'd12473: dataIn1 = 32'd414
; 
32'd12474: dataIn1 = 32'd434
; 
32'd12475: dataIn1 = 32'd449
; 
32'd12476: dataIn1 = 32'd471
; 
32'd12477: dataIn1 = 32'd479
; 
32'd12478: dataIn1 = 32'd505
; 
32'd12479: dataIn1 = 32'd526
; 
32'd12480: dataIn1 = 32'd531
; 
32'd12481: dataIn1 = 32'd538
; 
32'd12482: dataIn1 = 32'd547
; 
32'd12483: dataIn1 = 32'd558
; 
32'd12484: dataIn1 = 32'd588
; 
32'd12485: dataIn1 = 32'd609
; 
32'd12486: dataIn1 = 32'd624
; 
32'd12487: dataIn1 = 32'd632
; 
32'd12488: dataIn1 = 32'd647
; 
32'd12489: dataIn1 = 32'd706
; 
32'd12490: dataIn1 = 32'd711
; 
32'd12491: dataIn1 = 32'd769
; 
32'd12492: dataIn1 = 32'd777
; 
32'd12493: dataIn1 = 32'd114
; 
32'd12494: dataIn1 = 32'd120
; 
32'd12495: dataIn1 = 32'd127
; 
32'd12496: dataIn1 = 32'd143
; 
32'd12497: dataIn1 = 32'd180
; 
32'd12498: dataIn1 = 32'd202
; 
32'd12499: dataIn1 = 32'd203
; 
32'd12500: dataIn1 = 32'd205
; 
32'd12501: dataIn1 = 32'd207
; 
32'd12502: dataIn1 = 32'd218
; 
32'd12503: dataIn1 = 32'd219
; 
32'd12504: dataIn1 = 32'd228
; 
32'd12505: dataIn1 = 32'd244
; 
32'd12506: dataIn1 = 32'd265
; 
32'd12507: dataIn1 = 32'd285
; 
32'd12508: dataIn1 = 32'd293
; 
32'd12509: dataIn1 = 32'd315
; 
32'd12510: dataIn1 = 32'd333
; 
32'd12511: dataIn1 = 32'd336
; 
32'd12512: dataIn1 = 32'd345
; 
32'd12513: dataIn1 = 32'd346
; 
32'd12514: dataIn1 = 32'd354
; 
32'd12515: dataIn1 = 32'd363
; 
32'd12516: dataIn1 = 32'd380
; 
32'd12517: dataIn1 = 32'd384
; 
32'd12518: dataIn1 = 32'd386
; 
32'd12519: dataIn1 = 32'd399
; 
32'd12520: dataIn1 = 32'd414
; 
32'd12521: dataIn1 = 32'd450
; 
32'd12522: dataIn1 = 32'd473
; 
32'd12523: dataIn1 = 32'd509
; 
32'd12524: dataIn1 = 32'd511
; 
32'd12525: dataIn1 = 32'd513
; 
32'd12526: dataIn1 = 32'd524
; 
32'd12527: dataIn1 = 32'd526
; 
32'd12528: dataIn1 = 32'd533
; 
32'd12529: dataIn1 = 32'd576
; 
32'd12530: dataIn1 = 32'd591
; 
32'd12531: dataIn1 = 32'd611
; 
32'd12532: dataIn1 = 32'd624
; 
32'd12533: dataIn1 = 32'd636
; 
32'd12534: dataIn1 = 32'd659
; 
32'd12535: dataIn1 = 32'd684
; 
32'd12536: dataIn1 = 32'd696
; 
32'd12537: dataIn1 = 32'd700
; 
32'd12538: dataIn1 = 32'd701
; 
32'd12539: dataIn1 = 32'd705
; 
32'd12540: dataIn1 = 32'd731
; 
32'd12541: dataIn1 = 32'd738
; 
32'd12542: dataIn1 = 32'd771
; 
32'd12543: dataIn1 = 32'd781
; 
32'd12544: dataIn1 = 32'd167
; 
32'd12545: dataIn1 = 32'd218
; 
32'd12546: dataIn1 = 32'd258
; 
32'd12547: dataIn1 = 32'd263
; 
32'd12548: dataIn1 = 32'd264
; 
32'd12549: dataIn1 = 32'd278
; 
32'd12550: dataIn1 = 32'd304
; 
32'd12551: dataIn1 = 32'd314
; 
32'd12552: dataIn1 = 32'd338
; 
32'd12553: dataIn1 = 32'd356
; 
32'd12554: dataIn1 = 32'd377
; 
32'd12555: dataIn1 = 32'd398
; 
32'd12556: dataIn1 = 32'd413
; 
32'd12557: dataIn1 = 32'd422
; 
32'd12558: dataIn1 = 32'd426
; 
32'd12559: dataIn1 = 32'd441
; 
32'd12560: dataIn1 = 32'd452
; 
32'd12561: dataIn1 = 32'd465
; 
32'd12562: dataIn1 = 32'd477
; 
32'd12563: dataIn1 = 32'd504
; 
32'd12564: dataIn1 = 32'd505
; 
32'd12565: dataIn1 = 32'd508
; 
32'd12566: dataIn1 = 32'd515
; 
32'd12567: dataIn1 = 32'd590
; 
32'd12568: dataIn1 = 32'd611
; 
32'd12569: dataIn1 = 32'd618
; 
32'd12570: dataIn1 = 32'd711
; 
32'd12571: dataIn1 = 32'd743
; 
32'd12572: dataIn1 = 32'd748
; 
32'd12573: dataIn1 = 32'd761
; 
32'd12574: dataIn1 = 32'd770
; 
32'd12575: dataIn1 = 32'd776
; 
32'd12576: dataIn1 = 32'd777
; 
32'd12577: dataIn1 = 32'd784
; 
32'd12578: dataIn1 = 32'd789
; 
32'd12579: dataIn1 = 32'd165
; 
32'd12580: dataIn1 = 32'd181
; 
32'd12581: dataIn1 = 32'd189
; 
32'd12582: dataIn1 = 32'd190
; 
32'd12583: dataIn1 = 32'd196
; 
32'd12584: dataIn1 = 32'd214
; 
32'd12585: dataIn1 = 32'd280
; 
32'd12586: dataIn1 = 32'd283
; 
32'd12587: dataIn1 = 32'd299
; 
32'd12588: dataIn1 = 32'd301
; 
32'd12589: dataIn1 = 32'd308
; 
32'd12590: dataIn1 = 32'd334
; 
32'd12591: dataIn1 = 32'd346
; 
32'd12592: dataIn1 = 32'd351
; 
32'd12593: dataIn1 = 32'd357
; 
32'd12594: dataIn1 = 32'd362
; 
32'd12595: dataIn1 = 32'd368
; 
32'd12596: dataIn1 = 32'd399
; 
32'd12597: dataIn1 = 32'd430
; 
32'd12598: dataIn1 = 32'd433
; 
32'd12599: dataIn1 = 32'd442
; 
32'd12600: dataIn1 = 32'd446
; 
32'd12601: dataIn1 = 32'd449
; 
32'd12602: dataIn1 = 32'd476
; 
32'd12603: dataIn1 = 32'd568
; 
32'd12604: dataIn1 = 32'd604
; 
32'd12605: dataIn1 = 32'd640
; 
32'd12606: dataIn1 = 32'd649
; 
32'd12607: dataIn1 = 32'd670
; 
32'd12608: dataIn1 = 32'd680
; 
32'd12609: dataIn1 = 32'd702
; 
32'd12610: dataIn1 = 32'd722
; 
32'd12611: dataIn1 = 32'd752
; 
32'd12612: dataIn1 = 32'd788
; 
32'd12613: dataIn1 = 32'd107
; 
32'd12614: dataIn1 = 32'd120
; 
32'd12615: dataIn1 = 32'd144
; 
32'd12616: dataIn1 = 32'd153
; 
32'd12617: dataIn1 = 32'd157
; 
32'd12618: dataIn1 = 32'd190
; 
32'd12619: dataIn1 = 32'd211
; 
32'd12620: dataIn1 = 32'd253
; 
32'd12621: dataIn1 = 32'd300
; 
32'd12622: dataIn1 = 32'd309
; 
32'd12623: dataIn1 = 32'd334
; 
32'd12624: dataIn1 = 32'd340
; 
32'd12625: dataIn1 = 32'd346
; 
32'd12626: dataIn1 = 32'd368
; 
32'd12627: dataIn1 = 32'd388
; 
32'd12628: dataIn1 = 32'd390
; 
32'd12629: dataIn1 = 32'd410
; 
32'd12630: dataIn1 = 32'd426
; 
32'd12631: dataIn1 = 32'd454
; 
32'd12632: dataIn1 = 32'd490
; 
32'd12633: dataIn1 = 32'd514
; 
32'd12634: dataIn1 = 32'd525
; 
32'd12635: dataIn1 = 32'd536
; 
32'd12636: dataIn1 = 32'd559
; 
32'd12637: dataIn1 = 32'd588
; 
32'd12638: dataIn1 = 32'd605
; 
32'd12639: dataIn1 = 32'd621
; 
32'd12640: dataIn1 = 32'd622
; 
32'd12641: dataIn1 = 32'd627
; 
32'd12642: dataIn1 = 32'd675
; 
32'd12643: dataIn1 = 32'd680
; 
32'd12644: dataIn1 = 32'd684
; 
32'd12645: dataIn1 = 32'd689
; 
32'd12646: dataIn1 = 32'd703
; 
32'd12647: dataIn1 = 32'd732
; 
32'd12648: dataIn1 = 32'd747
; 
32'd12649: dataIn1 = 32'd752
; 
32'd12650: dataIn1 = 32'd783
; 
32'd12651: dataIn1 = 32'd792
; 
32'd12652: dataIn1 = 32'd112
; 
32'd12653: dataIn1 = 32'd133
; 
32'd12654: dataIn1 = 32'd139
; 
32'd12655: dataIn1 = 32'd144
; 
32'd12656: dataIn1 = 32'd152
; 
32'd12657: dataIn1 = 32'd189
; 
32'd12658: dataIn1 = 32'd190
; 
32'd12659: dataIn1 = 32'd208
; 
32'd12660: dataIn1 = 32'd261
; 
32'd12661: dataIn1 = 32'd269
; 
32'd12662: dataIn1 = 32'd271
; 
32'd12663: dataIn1 = 32'd280
; 
32'd12664: dataIn1 = 32'd294
; 
32'd12665: dataIn1 = 32'd300
; 
32'd12666: dataIn1 = 32'd339
; 
32'd12667: dataIn1 = 32'd345
; 
32'd12668: dataIn1 = 32'd353
; 
32'd12669: dataIn1 = 32'd370
; 
32'd12670: dataIn1 = 32'd381
; 
32'd12671: dataIn1 = 32'd383
; 
32'd12672: dataIn1 = 32'd389
; 
32'd12673: dataIn1 = 32'd395
; 
32'd12674: dataIn1 = 32'd398
; 
32'd12675: dataIn1 = 32'd455
; 
32'd12676: dataIn1 = 32'd473
; 
32'd12677: dataIn1 = 32'd487
; 
32'd12678: dataIn1 = 32'd508
; 
32'd12679: dataIn1 = 32'd509
; 
32'd12680: dataIn1 = 32'd549
; 
32'd12681: dataIn1 = 32'd562
; 
32'd12682: dataIn1 = 32'd598
; 
32'd12683: dataIn1 = 32'd614
; 
32'd12684: dataIn1 = 32'd637
; 
32'd12685: dataIn1 = 32'd658
; 
32'd12686: dataIn1 = 32'd678
; 
32'd12687: dataIn1 = 32'd693
; 
32'd12688: dataIn1 = 32'd702
; 
32'd12689: dataIn1 = 32'd721
; 
32'd12690: dataIn1 = 32'd737
; 
32'd12691: dataIn1 = 32'd753
; 
32'd12692: dataIn1 = 32'd755
; 
32'd12693: dataIn1 = 32'd769
; 
32'd12694: dataIn1 = 32'd776
; 
32'd12695: dataIn1 = 32'd799
; 
32'd12696: dataIn1 = 32'd144
; 
32'd12697: dataIn1 = 32'd161
; 
32'd12698: dataIn1 = 32'd162
; 
32'd12699: dataIn1 = 32'd176
; 
32'd12700: dataIn1 = 32'd187
; 
32'd12701: dataIn1 = 32'd220
; 
32'd12702: dataIn1 = 32'd233
; 
32'd12703: dataIn1 = 32'd240
; 
32'd12704: dataIn1 = 32'd256
; 
32'd12705: dataIn1 = 32'd264
; 
32'd12706: dataIn1 = 32'd280
; 
32'd12707: dataIn1 = 32'd316
; 
32'd12708: dataIn1 = 32'd332
; 
32'd12709: dataIn1 = 32'd336
; 
32'd12710: dataIn1 = 32'd343
; 
32'd12711: dataIn1 = 32'd353
; 
32'd12712: dataIn1 = 32'd363
; 
32'd12713: dataIn1 = 32'd378
; 
32'd12714: dataIn1 = 32'd392
; 
32'd12715: dataIn1 = 32'd412
; 
32'd12716: dataIn1 = 32'd483
; 
32'd12717: dataIn1 = 32'd489
; 
32'd12718: dataIn1 = 32'd493
; 
32'd12719: dataIn1 = 32'd508
; 
32'd12720: dataIn1 = 32'd516
; 
32'd12721: dataIn1 = 32'd541
; 
32'd12722: dataIn1 = 32'd549
; 
32'd12723: dataIn1 = 32'd557
; 
32'd12724: dataIn1 = 32'd582
; 
32'd12725: dataIn1 = 32'd592
; 
32'd12726: dataIn1 = 32'd608
; 
32'd12727: dataIn1 = 32'd638
; 
32'd12728: dataIn1 = 32'd666
; 
32'd12729: dataIn1 = 32'd668
; 
32'd12730: dataIn1 = 32'd681
; 
32'd12731: dataIn1 = 32'd692
; 
32'd12732: dataIn1 = 32'd709
; 
32'd12733: dataIn1 = 32'd710
; 
32'd12734: dataIn1 = 32'd717
; 
32'd12735: dataIn1 = 32'd765
; 
32'd12736: dataIn1 = 32'd788
; 
32'd12737: dataIn1 = 32'd133
; 
32'd12738: dataIn1 = 32'd144
; 
32'd12739: dataIn1 = 32'd158
; 
32'd12740: dataIn1 = 32'd161
; 
32'd12741: dataIn1 = 32'd178
; 
32'd12742: dataIn1 = 32'd198
; 
32'd12743: dataIn1 = 32'd200
; 
32'd12744: dataIn1 = 32'd222
; 
32'd12745: dataIn1 = 32'd258
; 
32'd12746: dataIn1 = 32'd275
; 
32'd12747: dataIn1 = 32'd277
; 
32'd12748: dataIn1 = 32'd278
; 
32'd12749: dataIn1 = 32'd286
; 
32'd12750: dataIn1 = 32'd303
; 
32'd12751: dataIn1 = 32'd338
; 
32'd12752: dataIn1 = 32'd353
; 
32'd12753: dataIn1 = 32'd374
; 
32'd12754: dataIn1 = 32'd405
; 
32'd12755: dataIn1 = 32'd414
; 
32'd12756: dataIn1 = 32'd423
; 
32'd12757: dataIn1 = 32'd427
; 
32'd12758: dataIn1 = 32'd460
; 
32'd12759: dataIn1 = 32'd472
; 
32'd12760: dataIn1 = 32'd525
; 
32'd12761: dataIn1 = 32'd535
; 
32'd12762: dataIn1 = 32'd583
; 
32'd12763: dataIn1 = 32'd599
; 
32'd12764: dataIn1 = 32'd619
; 
32'd12765: dataIn1 = 32'd657
; 
32'd12766: dataIn1 = 32'd679
; 
32'd12767: dataIn1 = 32'd694
; 
32'd12768: dataIn1 = 32'd702
; 
32'd12769: dataIn1 = 32'd703
; 
32'd12770: dataIn1 = 32'd717
; 
32'd12771: dataIn1 = 32'd739
; 
32'd12772: dataIn1 = 32'd743
; 
32'd12773: dataIn1 = 32'd764
; 
32'd12774: dataIn1 = 32'd789
; 
32'd12775: dataIn1 = 32'd794
; 
32'd12776: dataIn1 = 32'd796
; 
32'd12777: dataIn1 = 32'd115
; 
32'd12778: dataIn1 = 32'd146
; 
32'd12779: dataIn1 = 32'd150
; 
32'd12780: dataIn1 = 32'd199
; 
32'd12781: dataIn1 = 32'd217
; 
32'd12782: dataIn1 = 32'd238
; 
32'd12783: dataIn1 = 32'd311
; 
32'd12784: dataIn1 = 32'd319
; 
32'd12785: dataIn1 = 32'd346
; 
32'd12786: dataIn1 = 32'd366
; 
32'd12787: dataIn1 = 32'd397
; 
32'd12788: dataIn1 = 32'd409
; 
32'd12789: dataIn1 = 32'd416
; 
32'd12790: dataIn1 = 32'd481
; 
32'd12791: dataIn1 = 32'd487
; 
32'd12792: dataIn1 = 32'd493
; 
32'd12793: dataIn1 = 32'd511
; 
32'd12794: dataIn1 = 32'd525
; 
32'd12795: dataIn1 = 32'd531
; 
32'd12796: dataIn1 = 32'd543
; 
32'd12797: dataIn1 = 32'd589
; 
32'd12798: dataIn1 = 32'd592
; 
32'd12799: dataIn1 = 32'd607
; 
32'd12800: dataIn1 = 32'd615
; 
32'd12801: dataIn1 = 32'd655
; 
32'd12802: dataIn1 = 32'd673
; 
32'd12803: dataIn1 = 32'd676
; 
32'd12804: dataIn1 = 32'd710
; 
32'd12805: dataIn1 = 32'd781
; 
32'd12806: dataIn1 = 32'd124
; 
32'd12807: dataIn1 = 32'd131
; 
32'd12808: dataIn1 = 32'd151
; 
32'd12809: dataIn1 = 32'd152
; 
32'd12810: dataIn1 = 32'd156
; 
32'd12811: dataIn1 = 32'd200
; 
32'd12812: dataIn1 = 32'd210
; 
32'd12813: dataIn1 = 32'd215
; 
32'd12814: dataIn1 = 32'd275
; 
32'd12815: dataIn1 = 32'd283
; 
32'd12816: dataIn1 = 32'd289
; 
32'd12817: dataIn1 = 32'd309
; 
32'd12818: dataIn1 = 32'd326
; 
32'd12819: dataIn1 = 32'd329
; 
32'd12820: dataIn1 = 32'd356
; 
32'd12821: dataIn1 = 32'd371
; 
32'd12822: dataIn1 = 32'd377
; 
32'd12823: dataIn1 = 32'd400
; 
32'd12824: dataIn1 = 32'd421
; 
32'd12825: dataIn1 = 32'd437
; 
32'd12826: dataIn1 = 32'd441
; 
32'd12827: dataIn1 = 32'd451
; 
32'd12828: dataIn1 = 32'd458
; 
32'd12829: dataIn1 = 32'd466
; 
32'd12830: dataIn1 = 32'd467
; 
32'd12831: dataIn1 = 32'd470
; 
32'd12832: dataIn1 = 32'd471
; 
32'd12833: dataIn1 = 32'd480
; 
32'd12834: dataIn1 = 32'd493
; 
32'd12835: dataIn1 = 32'd576
; 
32'd12836: dataIn1 = 32'd585
; 
32'd12837: dataIn1 = 32'd589
; 
32'd12838: dataIn1 = 32'd635
; 
32'd12839: dataIn1 = 32'd643
; 
32'd12840: dataIn1 = 32'd712
; 
32'd12841: dataIn1 = 32'd716
; 
32'd12842: dataIn1 = 32'd790
; 
32'd12843: dataIn1 = 32'd791
; 
32'd12844: dataIn1 = 32'd113
; 
32'd12845: dataIn1 = 32'd117
; 
32'd12846: dataIn1 = 32'd137
; 
32'd12847: dataIn1 = 32'd145
; 
32'd12848: dataIn1 = 32'd150
; 
32'd12849: dataIn1 = 32'd204
; 
32'd12850: dataIn1 = 32'd212
; 
32'd12851: dataIn1 = 32'd215
; 
32'd12852: dataIn1 = 32'd234
; 
32'd12853: dataIn1 = 32'd270
; 
32'd12854: dataIn1 = 32'd286
; 
32'd12855: dataIn1 = 32'd287
; 
32'd12856: dataIn1 = 32'd292
; 
32'd12857: dataIn1 = 32'd299
; 
32'd12858: dataIn1 = 32'd343
; 
32'd12859: dataIn1 = 32'd377
; 
32'd12860: dataIn1 = 32'd378
; 
32'd12861: dataIn1 = 32'd388
; 
32'd12862: dataIn1 = 32'd389
; 
32'd12863: dataIn1 = 32'd460
; 
32'd12864: dataIn1 = 32'd475
; 
32'd12865: dataIn1 = 32'd482
; 
32'd12866: dataIn1 = 32'd574
; 
32'd12867: dataIn1 = 32'd602
; 
32'd12868: dataIn1 = 32'd612
; 
32'd12869: dataIn1 = 32'd613
; 
32'd12870: dataIn1 = 32'd630
; 
32'd12871: dataIn1 = 32'd643
; 
32'd12872: dataIn1 = 32'd646
; 
32'd12873: dataIn1 = 32'd666
; 
32'd12874: dataIn1 = 32'd677
; 
32'd12875: dataIn1 = 32'd678
; 
32'd12876: dataIn1 = 32'd684
; 
32'd12877: dataIn1 = 32'd687
; 
32'd12878: dataIn1 = 32'd688
; 
32'd12879: dataIn1 = 32'd721
; 
32'd12880: dataIn1 = 32'd759
; 
32'd12881: dataIn1 = 32'd769
; 
32'd12882: dataIn1 = 32'd770
; 
32'd12883: dataIn1 = 32'd772
; 
32'd12884: dataIn1 = 32'd787
; 
32'd12885: dataIn1 = 32'd795
; 
32'd12886: dataIn1 = 32'd129
; 
32'd12887: dataIn1 = 32'd138
; 
32'd12888: dataIn1 = 32'd165
; 
32'd12889: dataIn1 = 32'd196
; 
32'd12890: dataIn1 = 32'd221
; 
32'd12891: dataIn1 = 32'd225
; 
32'd12892: dataIn1 = 32'd243
; 
32'd12893: dataIn1 = 32'd263
; 
32'd12894: dataIn1 = 32'd281
; 
32'd12895: dataIn1 = 32'd310
; 
32'd12896: dataIn1 = 32'd359
; 
32'd12897: dataIn1 = 32'd369
; 
32'd12898: dataIn1 = 32'd389
; 
32'd12899: dataIn1 = 32'd416
; 
32'd12900: dataIn1 = 32'd427
; 
32'd12901: dataIn1 = 32'd453
; 
32'd12902: dataIn1 = 32'd487
; 
32'd12903: dataIn1 = 32'd502
; 
32'd12904: dataIn1 = 32'd506
; 
32'd12905: dataIn1 = 32'd522
; 
32'd12906: dataIn1 = 32'd562
; 
32'd12907: dataIn1 = 32'd574
; 
32'd12908: dataIn1 = 32'd578
; 
32'd12909: dataIn1 = 32'd592
; 
32'd12910: dataIn1 = 32'd600
; 
32'd12911: dataIn1 = 32'd605
; 
32'd12912: dataIn1 = 32'd611
; 
32'd12913: dataIn1 = 32'd623
; 
32'd12914: dataIn1 = 32'd633
; 
32'd12915: dataIn1 = 32'd634
; 
32'd12916: dataIn1 = 32'd667
; 
32'd12917: dataIn1 = 32'd668
; 
32'd12918: dataIn1 = 32'd678
; 
32'd12919: dataIn1 = 32'd706
; 
32'd12920: dataIn1 = 32'd719
; 
32'd12921: dataIn1 = 32'd722
; 
32'd12922: dataIn1 = 32'd726
; 
32'd12923: dataIn1 = 32'd727
; 
32'd12924: dataIn1 = 32'd773
; 
32'd12925: dataIn1 = 32'd785
; 
32'd12926: dataIn1 = 32'd125
; 
32'd12927: dataIn1 = 32'd141
; 
32'd12928: dataIn1 = 32'd157
; 
32'd12929: dataIn1 = 32'd204
; 
32'd12930: dataIn1 = 32'd228
; 
32'd12931: dataIn1 = 32'd240
; 
32'd12932: dataIn1 = 32'd254
; 
32'd12933: dataIn1 = 32'd275
; 
32'd12934: dataIn1 = 32'd277
; 
32'd12935: dataIn1 = 32'd284
; 
32'd12936: dataIn1 = 32'd287
; 
32'd12937: dataIn1 = 32'd294
; 
32'd12938: dataIn1 = 32'd339
; 
32'd12939: dataIn1 = 32'd341
; 
32'd12940: dataIn1 = 32'd360
; 
32'd12941: dataIn1 = 32'd384
; 
32'd12942: dataIn1 = 32'd412
; 
32'd12943: dataIn1 = 32'd426
; 
32'd12944: dataIn1 = 32'd444
; 
32'd12945: dataIn1 = 32'd449
; 
32'd12946: dataIn1 = 32'd479
; 
32'd12947: dataIn1 = 32'd491
; 
32'd12948: dataIn1 = 32'd498
; 
32'd12949: dataIn1 = 32'd516
; 
32'd12950: dataIn1 = 32'd537
; 
32'd12951: dataIn1 = 32'd542
; 
32'd12952: dataIn1 = 32'd552
; 
32'd12953: dataIn1 = 32'd560
; 
32'd12954: dataIn1 = 32'd561
; 
32'd12955: dataIn1 = 32'd620
; 
32'd12956: dataIn1 = 32'd645
; 
32'd12957: dataIn1 = 32'd672
; 
32'd12958: dataIn1 = 32'd686
; 
32'd12959: dataIn1 = 32'd691
; 
32'd12960: dataIn1 = 32'd719
; 
32'd12961: dataIn1 = 32'd720
; 
32'd12962: dataIn1 = 32'd731
; 
32'd12963: dataIn1 = 32'd744
; 
32'd12964: dataIn1 = 32'd764
; 
32'd12965: dataIn1 = 32'd765
; 
32'd12966: dataIn1 = 32'd767
; 
32'd12967: dataIn1 = 32'd783
; 
32'd12968: dataIn1 = 32'd796
; 
32'd12969: dataIn1 = 32'd122
; 
32'd12970: dataIn1 = 32'd136
; 
32'd12971: dataIn1 = 32'd154
; 
32'd12972: dataIn1 = 32'd172
; 
32'd12973: dataIn1 = 32'd198
; 
32'd12974: dataIn1 = 32'd219
; 
32'd12975: dataIn1 = 32'd294
; 
32'd12976: dataIn1 = 32'd335
; 
32'd12977: dataIn1 = 32'd340
; 
32'd12978: dataIn1 = 32'd355
; 
32'd12979: dataIn1 = 32'd359
; 
32'd12980: dataIn1 = 32'd364
; 
32'd12981: dataIn1 = 32'd373
; 
32'd12982: dataIn1 = 32'd437
; 
32'd12983: dataIn1 = 32'd447
; 
32'd12984: dataIn1 = 32'd509
; 
32'd12985: dataIn1 = 32'd533
; 
32'd12986: dataIn1 = 32'd569
; 
32'd12987: dataIn1 = 32'd602
; 
32'd12988: dataIn1 = 32'd613
; 
32'd12989: dataIn1 = 32'd617
; 
32'd12990: dataIn1 = 32'd660
; 
32'd12991: dataIn1 = 32'd674
; 
32'd12992: dataIn1 = 32'd685
; 
32'd12993: dataIn1 = 32'd689
; 
32'd12994: dataIn1 = 32'd692
; 
32'd12995: dataIn1 = 32'd700
; 
32'd12996: dataIn1 = 32'd713
; 
32'd12997: dataIn1 = 32'd741
; 
32'd12998: dataIn1 = 32'd763
; 
32'd12999: dataIn1 = 32'd125
; 
32'd13000: dataIn1 = 32'd138
; 
32'd13001: dataIn1 = 32'd145
; 
32'd13002: dataIn1 = 32'd157
; 
32'd13003: dataIn1 = 32'd158
; 
32'd13004: dataIn1 = 32'd160
; 
32'd13005: dataIn1 = 32'd163
; 
32'd13006: dataIn1 = 32'd174
; 
32'd13007: dataIn1 = 32'd193
; 
32'd13008: dataIn1 = 32'd198
; 
32'd13009: dataIn1 = 32'd201
; 
32'd13010: dataIn1 = 32'd205
; 
32'd13011: dataIn1 = 32'd229
; 
32'd13012: dataIn1 = 32'd239
; 
32'd13013: dataIn1 = 32'd241
; 
32'd13014: dataIn1 = 32'd243
; 
32'd13015: dataIn1 = 32'd253
; 
32'd13016: dataIn1 = 32'd264
; 
32'd13017: dataIn1 = 32'd266
; 
32'd13018: dataIn1 = 32'd290
; 
32'd13019: dataIn1 = 32'd335
; 
32'd13020: dataIn1 = 32'd350
; 
32'd13021: dataIn1 = 32'd351
; 
32'd13022: dataIn1 = 32'd360
; 
32'd13023: dataIn1 = 32'd388
; 
32'd13024: dataIn1 = 32'd391
; 
32'd13025: dataIn1 = 32'd403
; 
32'd13026: dataIn1 = 32'd462
; 
32'd13027: dataIn1 = 32'd466
; 
32'd13028: dataIn1 = 32'd533
; 
32'd13029: dataIn1 = 32'd540
; 
32'd13030: dataIn1 = 32'd559
; 
32'd13031: dataIn1 = 32'd577
; 
32'd13032: dataIn1 = 32'd578
; 
32'd13033: dataIn1 = 32'd588
; 
32'd13034: dataIn1 = 32'd602
; 
32'd13035: dataIn1 = 32'd607
; 
32'd13036: dataIn1 = 32'd611
; 
32'd13037: dataIn1 = 32'd623
; 
32'd13038: dataIn1 = 32'd651
; 
32'd13039: dataIn1 = 32'd662
; 
32'd13040: dataIn1 = 32'd670
; 
32'd13041: dataIn1 = 32'd677
; 
32'd13042: dataIn1 = 32'd685
; 
32'd13043: dataIn1 = 32'd696
; 
32'd13044: dataIn1 = 32'd718
; 
32'd13045: dataIn1 = 32'd733
; 
32'd13046: dataIn1 = 32'd763
; 
32'd13047: dataIn1 = 32'd769
; 
32'd13048: dataIn1 = 32'd772
; 
32'd13049: dataIn1 = 32'd781
; 
32'd13050: dataIn1 = 32'd117
; 
32'd13051: dataIn1 = 32'd119
; 
32'd13052: dataIn1 = 32'd157
; 
32'd13053: dataIn1 = 32'd167
; 
32'd13054: dataIn1 = 32'd254
; 
32'd13055: dataIn1 = 32'd257
; 
32'd13056: dataIn1 = 32'd274
; 
32'd13057: dataIn1 = 32'd288
; 
32'd13058: dataIn1 = 32'd315
; 
32'd13059: dataIn1 = 32'd339
; 
32'd13060: dataIn1 = 32'd365
; 
32'd13061: dataIn1 = 32'd398
; 
32'd13062: dataIn1 = 32'd422
; 
32'd13063: dataIn1 = 32'd435
; 
32'd13064: dataIn1 = 32'd442
; 
32'd13065: dataIn1 = 32'd456
; 
32'd13066: dataIn1 = 32'd467
; 
32'd13067: dataIn1 = 32'd477
; 
32'd13068: dataIn1 = 32'd485
; 
32'd13069: dataIn1 = 32'd486
; 
32'd13070: dataIn1 = 32'd491
; 
32'd13071: dataIn1 = 32'd499
; 
32'd13072: dataIn1 = 32'd558
; 
32'd13073: dataIn1 = 32'd562
; 
32'd13074: dataIn1 = 32'd574
; 
32'd13075: dataIn1 = 32'd638
; 
32'd13076: dataIn1 = 32'd639
; 
32'd13077: dataIn1 = 32'd642
; 
32'd13078: dataIn1 = 32'd648
; 
32'd13079: dataIn1 = 32'd674
; 
32'd13080: dataIn1 = 32'd740
; 
32'd13081: dataIn1 = 32'd751
; 
32'd13082: dataIn1 = 32'd773
; 
32'd13083: dataIn1 = 32'd774
; 
32'd13084: dataIn1 = 32'd788
; 
32'd13085: dataIn1 = 32'd796
; 
32'd13086: dataIn1 = 32'd125
; 
32'd13087: dataIn1 = 32'd140
; 
32'd13088: dataIn1 = 32'd197
; 
32'd13089: dataIn1 = 32'd199
; 
32'd13090: dataIn1 = 32'd205
; 
32'd13091: dataIn1 = 32'd283
; 
32'd13092: dataIn1 = 32'd285
; 
32'd13093: dataIn1 = 32'd291
; 
32'd13094: dataIn1 = 32'd293
; 
32'd13095: dataIn1 = 32'd330
; 
32'd13096: dataIn1 = 32'd370
; 
32'd13097: dataIn1 = 32'd375
; 
32'd13098: dataIn1 = 32'd414
; 
32'd13099: dataIn1 = 32'd446
; 
32'd13100: dataIn1 = 32'd472
; 
32'd13101: dataIn1 = 32'd475
; 
32'd13102: dataIn1 = 32'd504
; 
32'd13103: dataIn1 = 32'd556
; 
32'd13104: dataIn1 = 32'd589
; 
32'd13105: dataIn1 = 32'd612
; 
32'd13106: dataIn1 = 32'd617
; 
32'd13107: dataIn1 = 32'd629
; 
32'd13108: dataIn1 = 32'd640
; 
32'd13109: dataIn1 = 32'd689
; 
32'd13110: dataIn1 = 32'd690
; 
32'd13111: dataIn1 = 32'd694
; 
32'd13112: dataIn1 = 32'd716
; 
32'd13113: dataIn1 = 32'd719
; 
32'd13114: dataIn1 = 32'd741
; 
32'd13115: dataIn1 = 32'd756
; 
32'd13116: dataIn1 = 32'd757
; 
32'd13117: dataIn1 = 32'd774
; 
32'd13118: dataIn1 = 32'd779
; 
32'd13119: dataIn1 = 32'd781
; 
32'd13120: dataIn1 = 32'd783
; 
32'd13121: dataIn1 = 32'd127
; 
32'd13122: dataIn1 = 32'd128
; 
32'd13123: dataIn1 = 32'd139
; 
32'd13124: dataIn1 = 32'd151
; 
32'd13125: dataIn1 = 32'd233
; 
32'd13126: dataIn1 = 32'd235
; 
32'd13127: dataIn1 = 32'd237
; 
32'd13128: dataIn1 = 32'd246
; 
32'd13129: dataIn1 = 32'd252
; 
32'd13130: dataIn1 = 32'd265
; 
32'd13131: dataIn1 = 32'd275
; 
32'd13132: dataIn1 = 32'd292
; 
32'd13133: dataIn1 = 32'd293
; 
32'd13134: dataIn1 = 32'd302
; 
32'd13135: dataIn1 = 32'd322
; 
32'd13136: dataIn1 = 32'd326
; 
32'd13137: dataIn1 = 32'd330
; 
32'd13138: dataIn1 = 32'd338
; 
32'd13139: dataIn1 = 32'd354
; 
32'd13140: dataIn1 = 32'd385
; 
32'd13141: dataIn1 = 32'd438
; 
32'd13142: dataIn1 = 32'd453
; 
32'd13143: dataIn1 = 32'd473
; 
32'd13144: dataIn1 = 32'd496
; 
32'd13145: dataIn1 = 32'd530
; 
32'd13146: dataIn1 = 32'd536
; 
32'd13147: dataIn1 = 32'd551
; 
32'd13148: dataIn1 = 32'd595
; 
32'd13149: dataIn1 = 32'd685
; 
32'd13150: dataIn1 = 32'd689
; 
32'd13151: dataIn1 = 32'd707
; 
32'd13152: dataIn1 = 32'd717
; 
32'd13153: dataIn1 = 32'd718
; 
32'd13154: dataIn1 = 32'd734
; 
32'd13155: dataIn1 = 32'd735
; 
32'd13156: dataIn1 = 32'd749
; 
32'd13157: dataIn1 = 32'd764
; 
32'd13158: dataIn1 = 32'd784
; 
32'd13159: dataIn1 = 32'd126
; 
32'd13160: dataIn1 = 32'd130
; 
32'd13161: dataIn1 = 32'd146
; 
32'd13162: dataIn1 = 32'd174
; 
32'd13163: dataIn1 = 32'd185
; 
32'd13164: dataIn1 = 32'd186
; 
32'd13165: dataIn1 = 32'd199
; 
32'd13166: dataIn1 = 32'd222
; 
32'd13167: dataIn1 = 32'd234
; 
32'd13168: dataIn1 = 32'd246
; 
32'd13169: dataIn1 = 32'd252
; 
32'd13170: dataIn1 = 32'd264
; 
32'd13171: dataIn1 = 32'd268
; 
32'd13172: dataIn1 = 32'd287
; 
32'd13173: dataIn1 = 32'd297
; 
32'd13174: dataIn1 = 32'd311
; 
32'd13175: dataIn1 = 32'd312
; 
32'd13176: dataIn1 = 32'd313
; 
32'd13177: dataIn1 = 32'd316
; 
32'd13178: dataIn1 = 32'd318
; 
32'd13179: dataIn1 = 32'd326
; 
32'd13180: dataIn1 = 32'd331
; 
32'd13181: dataIn1 = 32'd341
; 
32'd13182: dataIn1 = 32'd344
; 
32'd13183: dataIn1 = 32'd348
; 
32'd13184: dataIn1 = 32'd353
; 
32'd13185: dataIn1 = 32'd362
; 
32'd13186: dataIn1 = 32'd369
; 
32'd13187: dataIn1 = 32'd402
; 
32'd13188: dataIn1 = 32'd415
; 
32'd13189: dataIn1 = 32'd428
; 
32'd13190: dataIn1 = 32'd454
; 
32'd13191: dataIn1 = 32'd460
; 
32'd13192: dataIn1 = 32'd473
; 
32'd13193: dataIn1 = 32'd491
; 
32'd13194: dataIn1 = 32'd531
; 
32'd13195: dataIn1 = 32'd534
; 
32'd13196: dataIn1 = 32'd536
; 
32'd13197: dataIn1 = 32'd537
; 
32'd13198: dataIn1 = 32'd573
; 
32'd13199: dataIn1 = 32'd575
; 
32'd13200: dataIn1 = 32'd620
; 
32'd13201: dataIn1 = 32'd644
; 
32'd13202: dataIn1 = 32'd648
; 
32'd13203: dataIn1 = 32'd659
; 
32'd13204: dataIn1 = 32'd663
; 
32'd13205: dataIn1 = 32'd777
; 
32'd13206: dataIn1 = 32'd799
; 
32'd13207: dataIn1 = 32'd128
; 
32'd13208: dataIn1 = 32'd160
; 
32'd13209: dataIn1 = 32'd209
; 
32'd13210: dataIn1 = 32'd240
; 
32'd13211: dataIn1 = 32'd249
; 
32'd13212: dataIn1 = 32'd252
; 
32'd13213: dataIn1 = 32'd259
; 
32'd13214: dataIn1 = 32'd267
; 
32'd13215: dataIn1 = 32'd281
; 
32'd13216: dataIn1 = 32'd287
; 
32'd13217: dataIn1 = 32'd288
; 
32'd13218: dataIn1 = 32'd292
; 
32'd13219: dataIn1 = 32'd305
; 
32'd13220: dataIn1 = 32'd326
; 
32'd13221: dataIn1 = 32'd337
; 
32'd13222: dataIn1 = 32'd338
; 
32'd13223: dataIn1 = 32'd359
; 
32'd13224: dataIn1 = 32'd370
; 
32'd13225: dataIn1 = 32'd376
; 
32'd13226: dataIn1 = 32'd380
; 
32'd13227: dataIn1 = 32'd450
; 
32'd13228: dataIn1 = 32'd466
; 
32'd13229: dataIn1 = 32'd501
; 
32'd13230: dataIn1 = 32'd525
; 
32'd13231: dataIn1 = 32'd538
; 
32'd13232: dataIn1 = 32'd542
; 
32'd13233: dataIn1 = 32'd552
; 
32'd13234: dataIn1 = 32'd606
; 
32'd13235: dataIn1 = 32'd614
; 
32'd13236: dataIn1 = 32'd626
; 
32'd13237: dataIn1 = 32'd642
; 
32'd13238: dataIn1 = 32'd679
; 
32'd13239: dataIn1 = 32'd684
; 
32'd13240: dataIn1 = 32'd687
; 
32'd13241: dataIn1 = 32'd730
; 
32'd13242: dataIn1 = 32'd756
; 
32'd13243: dataIn1 = 32'd770
; 
32'd13244: dataIn1 = 32'd797
; 
32'd13245: dataIn1 = 32'd133
; 
32'd13246: dataIn1 = 32'd145
; 
32'd13247: dataIn1 = 32'd147
; 
32'd13248: dataIn1 = 32'd153
; 
32'd13249: dataIn1 = 32'd164
; 
32'd13250: dataIn1 = 32'd178
; 
32'd13251: dataIn1 = 32'd191
; 
32'd13252: dataIn1 = 32'd202
; 
32'd13253: dataIn1 = 32'd228
; 
32'd13254: dataIn1 = 32'd238
; 
32'd13255: dataIn1 = 32'd263
; 
32'd13256: dataIn1 = 32'd301
; 
32'd13257: dataIn1 = 32'd322
; 
32'd13258: dataIn1 = 32'd378
; 
32'd13259: dataIn1 = 32'd380
; 
32'd13260: dataIn1 = 32'd407
; 
32'd13261: dataIn1 = 32'd426
; 
32'd13262: dataIn1 = 32'd439
; 
32'd13263: dataIn1 = 32'd446
; 
32'd13264: dataIn1 = 32'd452
; 
32'd13265: dataIn1 = 32'd460
; 
32'd13266: dataIn1 = 32'd461
; 
32'd13267: dataIn1 = 32'd487
; 
32'd13268: dataIn1 = 32'd488
; 
32'd13269: dataIn1 = 32'd491
; 
32'd13270: dataIn1 = 32'd495
; 
32'd13271: dataIn1 = 32'd505
; 
32'd13272: dataIn1 = 32'd542
; 
32'd13273: dataIn1 = 32'd558
; 
32'd13274: dataIn1 = 32'd575
; 
32'd13275: dataIn1 = 32'd580
; 
32'd13276: dataIn1 = 32'd607
; 
32'd13277: dataIn1 = 32'd610
; 
32'd13278: dataIn1 = 32'd637
; 
32'd13279: dataIn1 = 32'd655
; 
32'd13280: dataIn1 = 32'd690
; 
32'd13281: dataIn1 = 32'd691
; 
32'd13282: dataIn1 = 32'd714
; 
32'd13283: dataIn1 = 32'd725
; 
32'd13284: dataIn1 = 32'd735
; 
32'd13285: dataIn1 = 32'd189
; 
32'd13286: dataIn1 = 32'd196
; 
32'd13287: dataIn1 = 32'd217
; 
32'd13288: dataIn1 = 32'd239
; 
32'd13289: dataIn1 = 32'd247
; 
32'd13290: dataIn1 = 32'd270
; 
32'd13291: dataIn1 = 32'd286
; 
32'd13292: dataIn1 = 32'd288
; 
32'd13293: dataIn1 = 32'd317
; 
32'd13294: dataIn1 = 32'd318
; 
32'd13295: dataIn1 = 32'd321
; 
32'd13296: dataIn1 = 32'd337
; 
32'd13297: dataIn1 = 32'd343
; 
32'd13298: dataIn1 = 32'd385
; 
32'd13299: dataIn1 = 32'd392
; 
32'd13300: dataIn1 = 32'd409
; 
32'd13301: dataIn1 = 32'd425
; 
32'd13302: dataIn1 = 32'd444
; 
32'd13303: dataIn1 = 32'd449
; 
32'd13304: dataIn1 = 32'd457
; 
32'd13305: dataIn1 = 32'd470
; 
32'd13306: dataIn1 = 32'd478
; 
32'd13307: dataIn1 = 32'd493
; 
32'd13308: dataIn1 = 32'd531
; 
32'd13309: dataIn1 = 32'd553
; 
32'd13310: dataIn1 = 32'd599
; 
32'd13311: dataIn1 = 32'd613
; 
32'd13312: dataIn1 = 32'd626
; 
32'd13313: dataIn1 = 32'd685
; 
32'd13314: dataIn1 = 32'd741
; 
32'd13315: dataIn1 = 32'd754
; 
32'd13316: dataIn1 = 32'd766
; 
32'd13317: dataIn1 = 32'd135
; 
32'd13318: dataIn1 = 32'd158
; 
32'd13319: dataIn1 = 32'd168
; 
32'd13320: dataIn1 = 32'd170
; 
32'd13321: dataIn1 = 32'd190
; 
32'd13322: dataIn1 = 32'd204
; 
32'd13323: dataIn1 = 32'd219
; 
32'd13324: dataIn1 = 32'd225
; 
32'd13325: dataIn1 = 32'd239
; 
32'd13326: dataIn1 = 32'd251
; 
32'd13327: dataIn1 = 32'd254
; 
32'd13328: dataIn1 = 32'd267
; 
32'd13329: dataIn1 = 32'd270
; 
32'd13330: dataIn1 = 32'd278
; 
32'd13331: dataIn1 = 32'd286
; 
32'd13332: dataIn1 = 32'd309
; 
32'd13333: dataIn1 = 32'd314
; 
32'd13334: dataIn1 = 32'd328
; 
32'd13335: dataIn1 = 32'd336
; 
32'd13336: dataIn1 = 32'd338
; 
32'd13337: dataIn1 = 32'd344
; 
32'd13338: dataIn1 = 32'd367
; 
32'd13339: dataIn1 = 32'd382
; 
32'd13340: dataIn1 = 32'd386
; 
32'd13341: dataIn1 = 32'd388
; 
32'd13342: dataIn1 = 32'd396
; 
32'd13343: dataIn1 = 32'd397
; 
32'd13344: dataIn1 = 32'd411
; 
32'd13345: dataIn1 = 32'd419
; 
32'd13346: dataIn1 = 32'd424
; 
32'd13347: dataIn1 = 32'd514
; 
32'd13348: dataIn1 = 32'd529
; 
32'd13349: dataIn1 = 32'd540
; 
32'd13350: dataIn1 = 32'd544
; 
32'd13351: dataIn1 = 32'd568
; 
32'd13352: dataIn1 = 32'd569
; 
32'd13353: dataIn1 = 32'd570
; 
32'd13354: dataIn1 = 32'd572
; 
32'd13355: dataIn1 = 32'd638
; 
32'd13356: dataIn1 = 32'd641
; 
32'd13357: dataIn1 = 32'd661
; 
32'd13358: dataIn1 = 32'd670
; 
32'd13359: dataIn1 = 32'd693
; 
32'd13360: dataIn1 = 32'd732
; 
32'd13361: dataIn1 = 32'd737
; 
32'd13362: dataIn1 = 32'd754
; 
32'd13363: dataIn1 = 32'd758
; 
32'd13364: dataIn1 = 32'd762
; 
32'd13365: dataIn1 = 32'd768
; 
32'd13366: dataIn1 = 32'd774
; 
32'd13367: dataIn1 = 32'd786
; 
32'd13368: dataIn1 = 32'd789
; 
32'd13369: dataIn1 = 32'd128
; 
32'd13370: dataIn1 = 32'd138
; 
32'd13371: dataIn1 = 32'd168
; 
32'd13372: dataIn1 = 32'd169
; 
32'd13373: dataIn1 = 32'd240
; 
32'd13374: dataIn1 = 32'd249
; 
32'd13375: dataIn1 = 32'd274
; 
32'd13376: dataIn1 = 32'd326
; 
32'd13377: dataIn1 = 32'd331
; 
32'd13378: dataIn1 = 32'd350
; 
32'd13379: dataIn1 = 32'd396
; 
32'd13380: dataIn1 = 32'd402
; 
32'd13381: dataIn1 = 32'd409
; 
32'd13382: dataIn1 = 32'd422
; 
32'd13383: dataIn1 = 32'd426
; 
32'd13384: dataIn1 = 32'd431
; 
32'd13385: dataIn1 = 32'd450
; 
32'd13386: dataIn1 = 32'd469
; 
32'd13387: dataIn1 = 32'd486
; 
32'd13388: dataIn1 = 32'd541
; 
32'd13389: dataIn1 = 32'd542
; 
32'd13390: dataIn1 = 32'd548
; 
32'd13391: dataIn1 = 32'd565
; 
32'd13392: dataIn1 = 32'd567
; 
32'd13393: dataIn1 = 32'd574
; 
32'd13394: dataIn1 = 32'd582
; 
32'd13395: dataIn1 = 32'd592
; 
32'd13396: dataIn1 = 32'd597
; 
32'd13397: dataIn1 = 32'd617
; 
32'd13398: dataIn1 = 32'd632
; 
32'd13399: dataIn1 = 32'd678
; 
32'd13400: dataIn1 = 32'd686
; 
32'd13401: dataIn1 = 32'd691
; 
32'd13402: dataIn1 = 32'd694
; 
32'd13403: dataIn1 = 32'd743
; 
32'd13404: dataIn1 = 32'd755
; 
32'd13405: dataIn1 = 32'd758
; 
32'd13406: dataIn1 = 32'd762
; 
32'd13407: dataIn1 = 32'd767
; 
32'd13408: dataIn1 = 32'd785
; 
32'd13409: dataIn1 = 32'd133
; 
32'd13410: dataIn1 = 32'd142
; 
32'd13411: dataIn1 = 32'd153
; 
32'd13412: dataIn1 = 32'd157
; 
32'd13413: dataIn1 = 32'd181
; 
32'd13414: dataIn1 = 32'd186
; 
32'd13415: dataIn1 = 32'd204
; 
32'd13416: dataIn1 = 32'd221
; 
32'd13417: dataIn1 = 32'd242
; 
32'd13418: dataIn1 = 32'd269
; 
32'd13419: dataIn1 = 32'd271
; 
32'd13420: dataIn1 = 32'd277
; 
32'd13421: dataIn1 = 32'd279
; 
32'd13422: dataIn1 = 32'd281
; 
32'd13423: dataIn1 = 32'd292
; 
32'd13424: dataIn1 = 32'd294
; 
32'd13425: dataIn1 = 32'd307
; 
32'd13426: dataIn1 = 32'd316
; 
32'd13427: dataIn1 = 32'd330
; 
32'd13428: dataIn1 = 32'd357
; 
32'd13429: dataIn1 = 32'd363
; 
32'd13430: dataIn1 = 32'd367
; 
32'd13431: dataIn1 = 32'd389
; 
32'd13432: dataIn1 = 32'd404
; 
32'd13433: dataIn1 = 32'd410
; 
32'd13434: dataIn1 = 32'd416
; 
32'd13435: dataIn1 = 32'd434
; 
32'd13436: dataIn1 = 32'd443
; 
32'd13437: dataIn1 = 32'd457
; 
32'd13438: dataIn1 = 32'd484
; 
32'd13439: dataIn1 = 32'd506
; 
32'd13440: dataIn1 = 32'd517
; 
32'd13441: dataIn1 = 32'd524
; 
32'd13442: dataIn1 = 32'd530
; 
32'd13443: dataIn1 = 32'd536
; 
32'd13444: dataIn1 = 32'd540
; 
32'd13445: dataIn1 = 32'd570
; 
32'd13446: dataIn1 = 32'd571
; 
32'd13447: dataIn1 = 32'd596
; 
32'd13448: dataIn1 = 32'd600
; 
32'd13449: dataIn1 = 32'd664
; 
32'd13450: dataIn1 = 32'd671
; 
32'd13451: dataIn1 = 32'd674
; 
32'd13452: dataIn1 = 32'd682
; 
32'd13453: dataIn1 = 32'd692
; 
32'd13454: dataIn1 = 32'd702
; 
32'd13455: dataIn1 = 32'd733
; 
32'd13456: dataIn1 = 32'd748
; 
32'd13457: dataIn1 = 32'd774
; 
32'd13458: dataIn1 = 32'd783
; 
32'd13459: dataIn1 = 32'd800
; 
32'd13460: dataIn1 = 32'd127
; 
32'd13461: dataIn1 = 32'd146
; 
32'd13462: dataIn1 = 32'd151
; 
32'd13463: dataIn1 = 32'd157
; 
32'd13464: dataIn1 = 32'd201
; 
32'd13465: dataIn1 = 32'd207
; 
32'd13466: dataIn1 = 32'd214
; 
32'd13467: dataIn1 = 32'd224
; 
32'd13468: dataIn1 = 32'd256
; 
32'd13469: dataIn1 = 32'd265
; 
32'd13470: dataIn1 = 32'd282
; 
32'd13471: dataIn1 = 32'd308
; 
32'd13472: dataIn1 = 32'd309
; 
32'd13473: dataIn1 = 32'd317
; 
32'd13474: dataIn1 = 32'd318
; 
32'd13475: dataIn1 = 32'd319
; 
32'd13476: dataIn1 = 32'd321
; 
32'd13477: dataIn1 = 32'd376
; 
32'd13478: dataIn1 = 32'd384
; 
32'd13479: dataIn1 = 32'd385
; 
32'd13480: dataIn1 = 32'd418
; 
32'd13481: dataIn1 = 32'd445
; 
32'd13482: dataIn1 = 32'd464
; 
32'd13483: dataIn1 = 32'd515
; 
32'd13484: dataIn1 = 32'd520
; 
32'd13485: dataIn1 = 32'd539
; 
32'd13486: dataIn1 = 32'd561
; 
32'd13487: dataIn1 = 32'd584
; 
32'd13488: dataIn1 = 32'd643
; 
32'd13489: dataIn1 = 32'd654
; 
32'd13490: dataIn1 = 32'd662
; 
32'd13491: dataIn1 = 32'd664
; 
32'd13492: dataIn1 = 32'd675
; 
32'd13493: dataIn1 = 32'd710
; 
32'd13494: dataIn1 = 32'd719
; 
32'd13495: dataIn1 = 32'd761
; 
32'd13496: dataIn1 = 32'd780
; 
32'd13497: dataIn1 = 32'd797
; 
32'd13498: dataIn1 = 32'd132
; 
32'd13499: dataIn1 = 32'd136
; 
32'd13500: dataIn1 = 32'd154
; 
32'd13501: dataIn1 = 32'd169
; 
32'd13502: dataIn1 = 32'd211
; 
32'd13503: dataIn1 = 32'd302
; 
32'd13504: dataIn1 = 32'd317
; 
32'd13505: dataIn1 = 32'd326
; 
32'd13506: dataIn1 = 32'd328
; 
32'd13507: dataIn1 = 32'd340
; 
32'd13508: dataIn1 = 32'd349
; 
32'd13509: dataIn1 = 32'd351
; 
32'd13510: dataIn1 = 32'd381
; 
32'd13511: dataIn1 = 32'd412
; 
32'd13512: dataIn1 = 32'd470
; 
32'd13513: dataIn1 = 32'd484
; 
32'd13514: dataIn1 = 32'd546
; 
32'd13515: dataIn1 = 32'd554
; 
32'd13516: dataIn1 = 32'd561
; 
32'd13517: dataIn1 = 32'd599
; 
32'd13518: dataIn1 = 32'd632
; 
32'd13519: dataIn1 = 32'd666
; 
32'd13520: dataIn1 = 32'd688
; 
32'd13521: dataIn1 = 32'd703
; 
32'd13522: dataIn1 = 32'd718
; 
32'd13523: dataIn1 = 32'd734
; 
32'd13524: dataIn1 = 32'd790
; 
32'd13525: dataIn1 = 32'd161
; 
32'd13526: dataIn1 = 32'd184
; 
32'd13527: dataIn1 = 32'd185
; 
32'd13528: dataIn1 = 32'd193
; 
32'd13529: dataIn1 = 32'd201
; 
32'd13530: dataIn1 = 32'd229
; 
32'd13531: dataIn1 = 32'd232
; 
32'd13532: dataIn1 = 32'd236
; 
32'd13533: dataIn1 = 32'd256
; 
32'd13534: dataIn1 = 32'd259
; 
32'd13535: dataIn1 = 32'd289
; 
32'd13536: dataIn1 = 32'd304
; 
32'd13537: dataIn1 = 32'd314
; 
32'd13538: dataIn1 = 32'd374
; 
32'd13539: dataIn1 = 32'd413
; 
32'd13540: dataIn1 = 32'd483
; 
32'd13541: dataIn1 = 32'd544
; 
32'd13542: dataIn1 = 32'd545
; 
32'd13543: dataIn1 = 32'd552
; 
32'd13544: dataIn1 = 32'd568
; 
32'd13545: dataIn1 = 32'd589
; 
32'd13546: dataIn1 = 32'd617
; 
32'd13547: dataIn1 = 32'd639
; 
32'd13548: dataIn1 = 32'd681
; 
32'd13549: dataIn1 = 32'd692
; 
32'd13550: dataIn1 = 32'd701
; 
32'd13551: dataIn1 = 32'd710
; 
32'd13552: dataIn1 = 32'd752
; 
32'd13553: dataIn1 = 32'd769
; 
32'd13554: dataIn1 = 32'd772
; 
32'd13555: dataIn1 = 32'd777
; 
32'd13556: dataIn1 = 32'd136
; 
32'd13557: dataIn1 = 32'd147
; 
32'd13558: dataIn1 = 32'd150
; 
32'd13559: dataIn1 = 32'd152
; 
32'd13560: dataIn1 = 32'd166
; 
32'd13561: dataIn1 = 32'd169
; 
32'd13562: dataIn1 = 32'd203
; 
32'd13563: dataIn1 = 32'd250
; 
32'd13564: dataIn1 = 32'd264
; 
32'd13565: dataIn1 = 32'd277
; 
32'd13566: dataIn1 = 32'd299
; 
32'd13567: dataIn1 = 32'd317
; 
32'd13568: dataIn1 = 32'd324
; 
32'd13569: dataIn1 = 32'd329
; 
32'd13570: dataIn1 = 32'd353
; 
32'd13571: dataIn1 = 32'd402
; 
32'd13572: dataIn1 = 32'd414
; 
32'd13573: dataIn1 = 32'd421
; 
32'd13574: dataIn1 = 32'd452
; 
32'd13575: dataIn1 = 32'd500
; 
32'd13576: dataIn1 = 32'd518
; 
32'd13577: dataIn1 = 32'd561
; 
32'd13578: dataIn1 = 32'd641
; 
32'd13579: dataIn1 = 32'd655
; 
32'd13580: dataIn1 = 32'd687
; 
32'd13581: dataIn1 = 32'd689
; 
32'd13582: dataIn1 = 32'd692
; 
32'd13583: dataIn1 = 32'd715
; 
32'd13584: dataIn1 = 32'd724
; 
32'd13585: dataIn1 = 32'd736
; 
32'd13586: dataIn1 = 32'd749
; 
32'd13587: dataIn1 = 32'd763
; 
32'd13588: dataIn1 = 32'd767
; 
32'd13589: dataIn1 = 32'd787
; 
32'd13590: dataIn1 = 32'd789
; 
32'd13591: dataIn1 = 32'd798
; 
32'd13592: dataIn1 = 32'd800
; 
32'd13593: dataIn1 = 32'd135
; 
32'd13594: dataIn1 = 32'd136
; 
32'd13595: dataIn1 = 32'd150
; 
32'd13596: dataIn1 = 32'd179
; 
32'd13597: dataIn1 = 32'd181
; 
32'd13598: dataIn1 = 32'd183
; 
32'd13599: dataIn1 = 32'd205
; 
32'd13600: dataIn1 = 32'd207
; 
32'd13601: dataIn1 = 32'd218
; 
32'd13602: dataIn1 = 32'd309
; 
32'd13603: dataIn1 = 32'd353
; 
32'd13604: dataIn1 = 32'd360
; 
32'd13605: dataIn1 = 32'd418
; 
32'd13606: dataIn1 = 32'd421
; 
32'd13607: dataIn1 = 32'd434
; 
32'd13608: dataIn1 = 32'd454
; 
32'd13609: dataIn1 = 32'd474
; 
32'd13610: dataIn1 = 32'd485
; 
32'd13611: dataIn1 = 32'd492
; 
32'd13612: dataIn1 = 32'd497
; 
32'd13613: dataIn1 = 32'd521
; 
32'd13614: dataIn1 = 32'd536
; 
32'd13615: dataIn1 = 32'd539
; 
32'd13616: dataIn1 = 32'd558
; 
32'd13617: dataIn1 = 32'd565
; 
32'd13618: dataIn1 = 32'd567
; 
32'd13619: dataIn1 = 32'd571
; 
32'd13620: dataIn1 = 32'd575
; 
32'd13621: dataIn1 = 32'd585
; 
32'd13622: dataIn1 = 32'd588
; 
32'd13623: dataIn1 = 32'd618
; 
32'd13624: dataIn1 = 32'd620
; 
32'd13625: dataIn1 = 32'd628
; 
32'd13626: dataIn1 = 32'd655
; 
32'd13627: dataIn1 = 32'd670
; 
32'd13628: dataIn1 = 32'd680
; 
32'd13629: dataIn1 = 32'd682
; 
32'd13630: dataIn1 = 32'd703
; 
32'd13631: dataIn1 = 32'd717
; 
32'd13632: dataIn1 = 32'd751
; 
32'd13633: dataIn1 = 32'd758
; 
32'd13634: dataIn1 = 32'd765
; 
32'd13635: dataIn1 = 32'd774
; 
32'd13636: dataIn1 = 32'd787
; 
32'd13637: dataIn1 = 32'd138
; 
32'd13638: dataIn1 = 32'd145
; 
32'd13639: dataIn1 = 32'd171
; 
32'd13640: dataIn1 = 32'd192
; 
32'd13641: dataIn1 = 32'd218
; 
32'd13642: dataIn1 = 32'd224
; 
32'd13643: dataIn1 = 32'd293
; 
32'd13644: dataIn1 = 32'd340
; 
32'd13645: dataIn1 = 32'd365
; 
32'd13646: dataIn1 = 32'd367
; 
32'd13647: dataIn1 = 32'd368
; 
32'd13648: dataIn1 = 32'd372
; 
32'd13649: dataIn1 = 32'd383
; 
32'd13650: dataIn1 = 32'd384
; 
32'd13651: dataIn1 = 32'd389
; 
32'd13652: dataIn1 = 32'd402
; 
32'd13653: dataIn1 = 32'd412
; 
32'd13654: dataIn1 = 32'd420
; 
32'd13655: dataIn1 = 32'd433
; 
32'd13656: dataIn1 = 32'd439
; 
32'd13657: dataIn1 = 32'd452
; 
32'd13658: dataIn1 = 32'd476
; 
32'd13659: dataIn1 = 32'd489
; 
32'd13660: dataIn1 = 32'd512
; 
32'd13661: dataIn1 = 32'd521
; 
32'd13662: dataIn1 = 32'd544
; 
32'd13663: dataIn1 = 32'd551
; 
32'd13664: dataIn1 = 32'd554
; 
32'd13665: dataIn1 = 32'd557
; 
32'd13666: dataIn1 = 32'd611
; 
32'd13667: dataIn1 = 32'd614
; 
32'd13668: dataIn1 = 32'd638
; 
32'd13669: dataIn1 = 32'd659
; 
32'd13670: dataIn1 = 32'd660
; 
32'd13671: dataIn1 = 32'd661
; 
32'd13672: dataIn1 = 32'd691
; 
32'd13673: dataIn1 = 32'd725
; 
32'd13674: dataIn1 = 32'd731
; 
32'd13675: dataIn1 = 32'd754
; 
32'd13676: dataIn1 = 32'd799
; 
32'd13677: dataIn1 = 32'd142
; 
32'd13678: dataIn1 = 32'd144
; 
32'd13679: dataIn1 = 32'd169
; 
32'd13680: dataIn1 = 32'd175
; 
32'd13681: dataIn1 = 32'd177
; 
32'd13682: dataIn1 = 32'd218
; 
32'd13683: dataIn1 = 32'd225
; 
32'd13684: dataIn1 = 32'd246
; 
32'd13685: dataIn1 = 32'd265
; 
32'd13686: dataIn1 = 32'd285
; 
32'd13687: dataIn1 = 32'd298
; 
32'd13688: dataIn1 = 32'd329
; 
32'd13689: dataIn1 = 32'd347
; 
32'd13690: dataIn1 = 32'd374
; 
32'd13691: dataIn1 = 32'd380
; 
32'd13692: dataIn1 = 32'd387
; 
32'd13693: dataIn1 = 32'd390
; 
32'd13694: dataIn1 = 32'd399
; 
32'd13695: dataIn1 = 32'd403
; 
32'd13696: dataIn1 = 32'd425
; 
32'd13697: dataIn1 = 32'd433
; 
32'd13698: dataIn1 = 32'd438
; 
32'd13699: dataIn1 = 32'd463
; 
32'd13700: dataIn1 = 32'd503
; 
32'd13701: dataIn1 = 32'd504
; 
32'd13702: dataIn1 = 32'd509
; 
32'd13703: dataIn1 = 32'd552
; 
32'd13704: dataIn1 = 32'd556
; 
32'd13705: dataIn1 = 32'd560
; 
32'd13706: dataIn1 = 32'd595
; 
32'd13707: dataIn1 = 32'd605
; 
32'd13708: dataIn1 = 32'd615
; 
32'd13709: dataIn1 = 32'd630
; 
32'd13710: dataIn1 = 32'd635
; 
32'd13711: dataIn1 = 32'd648
; 
32'd13712: dataIn1 = 32'd668
; 
32'd13713: dataIn1 = 32'd713
; 
32'd13714: dataIn1 = 32'd729
; 
32'd13715: dataIn1 = 32'd740
; 
32'd13716: dataIn1 = 32'd762
; 
32'd13717: dataIn1 = 32'd768
; 
32'd13718: dataIn1 = 32'd782
; 
32'd13719: dataIn1 = 32'd144
; 
32'd13720: dataIn1 = 32'd171
; 
32'd13721: dataIn1 = 32'd204
; 
32'd13722: dataIn1 = 32'd216
; 
32'd13723: dataIn1 = 32'd223
; 
32'd13724: dataIn1 = 32'd227
; 
32'd13725: dataIn1 = 32'd237
; 
32'd13726: dataIn1 = 32'd246
; 
32'd13727: dataIn1 = 32'd281
; 
32'd13728: dataIn1 = 32'd289
; 
32'd13729: dataIn1 = 32'd294
; 
32'd13730: dataIn1 = 32'd306
; 
32'd13731: dataIn1 = 32'd337
; 
32'd13732: dataIn1 = 32'd351
; 
32'd13733: dataIn1 = 32'd359
; 
32'd13734: dataIn1 = 32'd397
; 
32'd13735: dataIn1 = 32'd403
; 
32'd13736: dataIn1 = 32'd441
; 
32'd13737: dataIn1 = 32'd445
; 
32'd13738: dataIn1 = 32'd476
; 
32'd13739: dataIn1 = 32'd484
; 
32'd13740: dataIn1 = 32'd499
; 
32'd13741: dataIn1 = 32'd515
; 
32'd13742: dataIn1 = 32'd521
; 
32'd13743: dataIn1 = 32'd587
; 
32'd13744: dataIn1 = 32'd591
; 
32'd13745: dataIn1 = 32'd628
; 
32'd13746: dataIn1 = 32'd637
; 
32'd13747: dataIn1 = 32'd647
; 
32'd13748: dataIn1 = 32'd704
; 
32'd13749: dataIn1 = 32'd709
; 
32'd13750: dataIn1 = 32'd711
; 
32'd13751: dataIn1 = 32'd738
; 
32'd13752: dataIn1 = 32'd800
; 
32'd13753: dataIn1 = 32'd158
; 
32'd13754: dataIn1 = 32'd188
; 
32'd13755: dataIn1 = 32'd250
; 
32'd13756: dataIn1 = 32'd293
; 
32'd13757: dataIn1 = 32'd323
; 
32'd13758: dataIn1 = 32'd335
; 
32'd13759: dataIn1 = 32'd338
; 
32'd13760: dataIn1 = 32'd346
; 
32'd13761: dataIn1 = 32'd349
; 
32'd13762: dataIn1 = 32'd356
; 
32'd13763: dataIn1 = 32'd361
; 
32'd13764: dataIn1 = 32'd423
; 
32'd13765: dataIn1 = 32'd431
; 
32'd13766: dataIn1 = 32'd451
; 
32'd13767: dataIn1 = 32'd454
; 
32'd13768: dataIn1 = 32'd459
; 
32'd13769: dataIn1 = 32'd466
; 
32'd13770: dataIn1 = 32'd472
; 
32'd13771: dataIn1 = 32'd473
; 
32'd13772: dataIn1 = 32'd480
; 
32'd13773: dataIn1 = 32'd483
; 
32'd13774: dataIn1 = 32'd489
; 
32'd13775: dataIn1 = 32'd490
; 
32'd13776: dataIn1 = 32'd520
; 
32'd13777: dataIn1 = 32'd527
; 
32'd13778: dataIn1 = 32'd529
; 
32'd13779: dataIn1 = 32'd540
; 
32'd13780: dataIn1 = 32'd548
; 
32'd13781: dataIn1 = 32'd556
; 
32'd13782: dataIn1 = 32'd561
; 
32'd13783: dataIn1 = 32'd575
; 
32'd13784: dataIn1 = 32'd586
; 
32'd13785: dataIn1 = 32'd589
; 
32'd13786: dataIn1 = 32'd617
; 
32'd13787: dataIn1 = 32'd623
; 
32'd13788: dataIn1 = 32'd647
; 
32'd13789: dataIn1 = 32'd686
; 
32'd13790: dataIn1 = 32'd703
; 
32'd13791: dataIn1 = 32'd722
; 
32'd13792: dataIn1 = 32'd793
; 
32'd13793: dataIn1 = 32'd158
; 
32'd13794: dataIn1 = 32'd178
; 
32'd13795: dataIn1 = 32'd182
; 
32'd13796: dataIn1 = 32'd190
; 
32'd13797: dataIn1 = 32'd220
; 
32'd13798: dataIn1 = 32'd241
; 
32'd13799: dataIn1 = 32'd244
; 
32'd13800: dataIn1 = 32'd245
; 
32'd13801: dataIn1 = 32'd290
; 
32'd13802: dataIn1 = 32'd305
; 
32'd13803: dataIn1 = 32'd324
; 
32'd13804: dataIn1 = 32'd335
; 
32'd13805: dataIn1 = 32'd344
; 
32'd13806: dataIn1 = 32'd363
; 
32'd13807: dataIn1 = 32'd444
; 
32'd13808: dataIn1 = 32'd454
; 
32'd13809: dataIn1 = 32'd465
; 
32'd13810: dataIn1 = 32'd498
; 
32'd13811: dataIn1 = 32'd539
; 
32'd13812: dataIn1 = 32'd542
; 
32'd13813: dataIn1 = 32'd548
; 
32'd13814: dataIn1 = 32'd589
; 
32'd13815: dataIn1 = 32'd632
; 
32'd13816: dataIn1 = 32'd634
; 
32'd13817: dataIn1 = 32'd650
; 
32'd13818: dataIn1 = 32'd663
; 
32'd13819: dataIn1 = 32'd670
; 
32'd13820: dataIn1 = 32'd695
; 
32'd13821: dataIn1 = 32'd708
; 
32'd13822: dataIn1 = 32'd752
; 
32'd13823: dataIn1 = 32'd150
; 
32'd13824: dataIn1 = 32'd164
; 
32'd13825: dataIn1 = 32'd171
; 
32'd13826: dataIn1 = 32'd205
; 
32'd13827: dataIn1 = 32'd220
; 
32'd13828: dataIn1 = 32'd227
; 
32'd13829: dataIn1 = 32'd229
; 
32'd13830: dataIn1 = 32'd243
; 
32'd13831: dataIn1 = 32'd250
; 
32'd13832: dataIn1 = 32'd255
; 
32'd13833: dataIn1 = 32'd270
; 
32'd13834: dataIn1 = 32'd272
; 
32'd13835: dataIn1 = 32'd277
; 
32'd13836: dataIn1 = 32'd295
; 
32'd13837: dataIn1 = 32'd396
; 
32'd13838: dataIn1 = 32'd401
; 
32'd13839: dataIn1 = 32'd460
; 
32'd13840: dataIn1 = 32'd468
; 
32'd13841: dataIn1 = 32'd496
; 
32'd13842: dataIn1 = 32'd510
; 
32'd13843: dataIn1 = 32'd519
; 
32'd13844: dataIn1 = 32'd528
; 
32'd13845: dataIn1 = 32'd554
; 
32'd13846: dataIn1 = 32'd566
; 
32'd13847: dataIn1 = 32'd567
; 
32'd13848: dataIn1 = 32'd581
; 
32'd13849: dataIn1 = 32'd624
; 
32'd13850: dataIn1 = 32'd628
; 
32'd13851: dataIn1 = 32'd644
; 
32'd13852: dataIn1 = 32'd650
; 
32'd13853: dataIn1 = 32'd690
; 
32'd13854: dataIn1 = 32'd691
; 
32'd13855: dataIn1 = 32'd693
; 
32'd13856: dataIn1 = 32'd700
; 
32'd13857: dataIn1 = 32'd711
; 
32'd13858: dataIn1 = 32'd792
; 
32'd13859: dataIn1 = 32'd142
; 
32'd13860: dataIn1 = 32'd150
; 
32'd13861: dataIn1 = 32'd170
; 
32'd13862: dataIn1 = 32'd185
; 
32'd13863: dataIn1 = 32'd209
; 
32'd13864: dataIn1 = 32'd211
; 
32'd13865: dataIn1 = 32'd232
; 
32'd13866: dataIn1 = 32'd241
; 
32'd13867: dataIn1 = 32'd253
; 
32'd13868: dataIn1 = 32'd281
; 
32'd13869: dataIn1 = 32'd290
; 
32'd13870: dataIn1 = 32'd300
; 
32'd13871: dataIn1 = 32'd320
; 
32'd13872: dataIn1 = 32'd328
; 
32'd13873: dataIn1 = 32'd364
; 
32'd13874: dataIn1 = 32'd372
; 
32'd13875: dataIn1 = 32'd376
; 
32'd13876: dataIn1 = 32'd380
; 
32'd13877: dataIn1 = 32'd382
; 
32'd13878: dataIn1 = 32'd396
; 
32'd13879: dataIn1 = 32'd407
; 
32'd13880: dataIn1 = 32'd420
; 
32'd13881: dataIn1 = 32'd437
; 
32'd13882: dataIn1 = 32'd480
; 
32'd13883: dataIn1 = 32'd484
; 
32'd13884: dataIn1 = 32'd499
; 
32'd13885: dataIn1 = 32'd505
; 
32'd13886: dataIn1 = 32'd512
; 
32'd13887: dataIn1 = 32'd605
; 
32'd13888: dataIn1 = 32'd617
; 
32'd13889: dataIn1 = 32'd643
; 
32'd13890: dataIn1 = 32'd645
; 
32'd13891: dataIn1 = 32'd656
; 
32'd13892: dataIn1 = 32'd683
; 
32'd13893: dataIn1 = 32'd684
; 
32'd13894: dataIn1 = 32'd686
; 
32'd13895: dataIn1 = 32'd705
; 
32'd13896: dataIn1 = 32'd740
; 
32'd13897: dataIn1 = 32'd772
; 
32'd13898: dataIn1 = 32'd800
; 
32'd13899: dataIn1 = 32'd149
; 
32'd13900: dataIn1 = 32'd205
; 
32'd13901: dataIn1 = 32'd213
; 
32'd13902: dataIn1 = 32'd243
; 
32'd13903: dataIn1 = 32'd251
; 
32'd13904: dataIn1 = 32'd257
; 
32'd13905: dataIn1 = 32'd265
; 
32'd13906: dataIn1 = 32'd272
; 
32'd13907: dataIn1 = 32'd273
; 
32'd13908: dataIn1 = 32'd280
; 
32'd13909: dataIn1 = 32'd289
; 
32'd13910: dataIn1 = 32'd312
; 
32'd13911: dataIn1 = 32'd323
; 
32'd13912: dataIn1 = 32'd338
; 
32'd13913: dataIn1 = 32'd353
; 
32'd13914: dataIn1 = 32'd366
; 
32'd13915: dataIn1 = 32'd369
; 
32'd13916: dataIn1 = 32'd422
; 
32'd13917: dataIn1 = 32'd431
; 
32'd13918: dataIn1 = 32'd440
; 
32'd13919: dataIn1 = 32'd441
; 
32'd13920: dataIn1 = 32'd463
; 
32'd13921: dataIn1 = 32'd466
; 
32'd13922: dataIn1 = 32'd467
; 
32'd13923: dataIn1 = 32'd470
; 
32'd13924: dataIn1 = 32'd498
; 
32'd13925: dataIn1 = 32'd532
; 
32'd13926: dataIn1 = 32'd535
; 
32'd13927: dataIn1 = 32'd545
; 
32'd13928: dataIn1 = 32'd562
; 
32'd13929: dataIn1 = 32'd648
; 
32'd13930: dataIn1 = 32'd677
; 
32'd13931: dataIn1 = 32'd687
; 
32'd13932: dataIn1 = 32'd692
; 
32'd13933: dataIn1 = 32'd700
; 
32'd13934: dataIn1 = 32'd716
; 
32'd13935: dataIn1 = 32'd729
; 
32'd13936: dataIn1 = 32'd751
; 
32'd13937: dataIn1 = 32'd774
; 
32'd13938: dataIn1 = 32'd775
; 
32'd13939: dataIn1 = 32'd787
; 
32'd13940: dataIn1 = 32'd157
; 
32'd13941: dataIn1 = 32'd172
; 
32'd13942: dataIn1 = 32'd195
; 
32'd13943: dataIn1 = 32'd220
; 
32'd13944: dataIn1 = 32'd228
; 
32'd13945: dataIn1 = 32'd234
; 
32'd13946: dataIn1 = 32'd262
; 
32'd13947: dataIn1 = 32'd267
; 
32'd13948: dataIn1 = 32'd321
; 
32'd13949: dataIn1 = 32'd338
; 
32'd13950: dataIn1 = 32'd382
; 
32'd13951: dataIn1 = 32'd388
; 
32'd13952: dataIn1 = 32'd405
; 
32'd13953: dataIn1 = 32'd408
; 
32'd13954: dataIn1 = 32'd410
; 
32'd13955: dataIn1 = 32'd415
; 
32'd13956: dataIn1 = 32'd427
; 
32'd13957: dataIn1 = 32'd428
; 
32'd13958: dataIn1 = 32'd430
; 
32'd13959: dataIn1 = 32'd456
; 
32'd13960: dataIn1 = 32'd459
; 
32'd13961: dataIn1 = 32'd484
; 
32'd13962: dataIn1 = 32'd490
; 
32'd13963: dataIn1 = 32'd491
; 
32'd13964: dataIn1 = 32'd500
; 
32'd13965: dataIn1 = 32'd522
; 
32'd13966: dataIn1 = 32'd524
; 
32'd13967: dataIn1 = 32'd531
; 
32'd13968: dataIn1 = 32'd536
; 
32'd13969: dataIn1 = 32'd541
; 
32'd13970: dataIn1 = 32'd543
; 
32'd13971: dataIn1 = 32'd554
; 
32'd13972: dataIn1 = 32'd556
; 
32'd13973: dataIn1 = 32'd610
; 
32'd13974: dataIn1 = 32'd646
; 
32'd13975: dataIn1 = 32'd658
; 
32'd13976: dataIn1 = 32'd682
; 
32'd13977: dataIn1 = 32'd702
; 
32'd13978: dataIn1 = 32'd764
; 
32'd13979: dataIn1 = 32'd767
; 
32'd13980: dataIn1 = 32'd775
; 
32'd13981: dataIn1 = 32'd147
; 
32'd13982: dataIn1 = 32'd170
; 
32'd13983: dataIn1 = 32'd181
; 
32'd13984: dataIn1 = 32'd184
; 
32'd13985: dataIn1 = 32'd207
; 
32'd13986: dataIn1 = 32'd227
; 
32'd13987: dataIn1 = 32'd231
; 
32'd13988: dataIn1 = 32'd239
; 
32'd13989: dataIn1 = 32'd244
; 
32'd13990: dataIn1 = 32'd249
; 
32'd13991: dataIn1 = 32'd261
; 
32'd13992: dataIn1 = 32'd283
; 
32'd13993: dataIn1 = 32'd306
; 
32'd13994: dataIn1 = 32'd309
; 
32'd13995: dataIn1 = 32'd374
; 
32'd13996: dataIn1 = 32'd454
; 
32'd13997: dataIn1 = 32'd477
; 
32'd13998: dataIn1 = 32'd483
; 
32'd13999: dataIn1 = 32'd488
; 
32'd14000: dataIn1 = 32'd522
; 
32'd14001: dataIn1 = 32'd538
; 
32'd14002: dataIn1 = 32'd551
; 
32'd14003: dataIn1 = 32'd561
; 
32'd14004: dataIn1 = 32'd583
; 
32'd14005: dataIn1 = 32'd627
; 
32'd14006: dataIn1 = 32'd630
; 
32'd14007: dataIn1 = 32'd631
; 
32'd14008: dataIn1 = 32'd649
; 
32'd14009: dataIn1 = 32'd652
; 
32'd14010: dataIn1 = 32'd675
; 
32'd14011: dataIn1 = 32'd682
; 
32'd14012: dataIn1 = 32'd684
; 
32'd14013: dataIn1 = 32'd771
; 
32'd14014: dataIn1 = 32'd797
; 
32'd14015: dataIn1 = 32'd799
; 
32'd14016: dataIn1 = 32'd154
; 
32'd14017: dataIn1 = 32'd178
; 
32'd14018: dataIn1 = 32'd192
; 
32'd14019: dataIn1 = 32'd199
; 
32'd14020: dataIn1 = 32'd243
; 
32'd14021: dataIn1 = 32'd274
; 
32'd14022: dataIn1 = 32'd282
; 
32'd14023: dataIn1 = 32'd288
; 
32'd14024: dataIn1 = 32'd294
; 
32'd14025: dataIn1 = 32'd321
; 
32'd14026: dataIn1 = 32'd349
; 
32'd14027: dataIn1 = 32'd363
; 
32'd14028: dataIn1 = 32'd371
; 
32'd14029: dataIn1 = 32'd400
; 
32'd14030: dataIn1 = 32'd405
; 
32'd14031: dataIn1 = 32'd419
; 
32'd14032: dataIn1 = 32'd422
; 
32'd14033: dataIn1 = 32'd439
; 
32'd14034: dataIn1 = 32'd440
; 
32'd14035: dataIn1 = 32'd450
; 
32'd14036: dataIn1 = 32'd455
; 
32'd14037: dataIn1 = 32'd467
; 
32'd14038: dataIn1 = 32'd476
; 
32'd14039: dataIn1 = 32'd542
; 
32'd14040: dataIn1 = 32'd547
; 
32'd14041: dataIn1 = 32'd555
; 
32'd14042: dataIn1 = 32'd606
; 
32'd14043: dataIn1 = 32'd644
; 
32'd14044: dataIn1 = 32'd649
; 
32'd14045: dataIn1 = 32'd656
; 
32'd14046: dataIn1 = 32'd659
; 
32'd14047: dataIn1 = 32'd661
; 
32'd14048: dataIn1 = 32'd674
; 
32'd14049: dataIn1 = 32'd698
; 
32'd14050: dataIn1 = 32'd700
; 
32'd14051: dataIn1 = 32'd730
; 
32'd14052: dataIn1 = 32'd733
; 
32'd14053: dataIn1 = 32'd737
; 
32'd14054: dataIn1 = 32'd753
; 
32'd14055: dataIn1 = 32'd773
; 
32'd14056: dataIn1 = 32'd788
; 
32'd14057: dataIn1 = 32'd798
; 
32'd14058: dataIn1 = 32'd148
; 
32'd14059: dataIn1 = 32'd151
; 
32'd14060: dataIn1 = 32'd152
; 
32'd14061: dataIn1 = 32'd165
; 
32'd14062: dataIn1 = 32'd196
; 
32'd14063: dataIn1 = 32'd200
; 
32'd14064: dataIn1 = 32'd202
; 
32'd14065: dataIn1 = 32'd208
; 
32'd14066: dataIn1 = 32'd211
; 
32'd14067: dataIn1 = 32'd227
; 
32'd14068: dataIn1 = 32'd237
; 
32'd14069: dataIn1 = 32'd247
; 
32'd14070: dataIn1 = 32'd252
; 
32'd14071: dataIn1 = 32'd262
; 
32'd14072: dataIn1 = 32'd273
; 
32'd14073: dataIn1 = 32'd299
; 
32'd14074: dataIn1 = 32'd311
; 
32'd14075: dataIn1 = 32'd324
; 
32'd14076: dataIn1 = 32'd330
; 
32'd14077: dataIn1 = 32'd338
; 
32'd14078: dataIn1 = 32'd339
; 
32'd14079: dataIn1 = 32'd344
; 
32'd14080: dataIn1 = 32'd360
; 
32'd14081: dataIn1 = 32'd372
; 
32'd14082: dataIn1 = 32'd400
; 
32'd14083: dataIn1 = 32'd414
; 
32'd14084: dataIn1 = 32'd415
; 
32'd14085: dataIn1 = 32'd433
; 
32'd14086: dataIn1 = 32'd443
; 
32'd14087: dataIn1 = 32'd448
; 
32'd14088: dataIn1 = 32'd465
; 
32'd14089: dataIn1 = 32'd511
; 
32'd14090: dataIn1 = 32'd533
; 
32'd14091: dataIn1 = 32'd560
; 
32'd14092: dataIn1 = 32'd573
; 
32'd14093: dataIn1 = 32'd587
; 
32'd14094: dataIn1 = 32'd606
; 
32'd14095: dataIn1 = 32'd633
; 
32'd14096: dataIn1 = 32'd657
; 
32'd14097: dataIn1 = 32'd702
; 
32'd14098: dataIn1 = 32'd704
; 
32'd14099: dataIn1 = 32'd721
; 
32'd14100: dataIn1 = 32'd757
; 
32'd14101: dataIn1 = 32'd765
; 
32'd14102: dataIn1 = 32'd776
; 
32'd14103: dataIn1 = 32'd791
; 
32'd14104: dataIn1 = 32'd797
; 
32'd14105: dataIn1 = 32'd155
; 
32'd14106: dataIn1 = 32'd162
; 
32'd14107: dataIn1 = 32'd179
; 
32'd14108: dataIn1 = 32'd182
; 
32'd14109: dataIn1 = 32'd183
; 
32'd14110: dataIn1 = 32'd185
; 
32'd14111: dataIn1 = 32'd189
; 
32'd14112: dataIn1 = 32'd194
; 
32'd14113: dataIn1 = 32'd228
; 
32'd14114: dataIn1 = 32'd236
; 
32'd14115: dataIn1 = 32'd239
; 
32'd14116: dataIn1 = 32'd252
; 
32'd14117: dataIn1 = 32'd261
; 
32'd14118: dataIn1 = 32'd264
; 
32'd14119: dataIn1 = 32'd281
; 
32'd14120: dataIn1 = 32'd291
; 
32'd14121: dataIn1 = 32'd310
; 
32'd14122: dataIn1 = 32'd334
; 
32'd14123: dataIn1 = 32'd340
; 
32'd14124: dataIn1 = 32'd354
; 
32'd14125: dataIn1 = 32'd370
; 
32'd14126: dataIn1 = 32'd377
; 
32'd14127: dataIn1 = 32'd387
; 
32'd14128: dataIn1 = 32'd400
; 
32'd14129: dataIn1 = 32'd416
; 
32'd14130: dataIn1 = 32'd428
; 
32'd14131: dataIn1 = 32'd431
; 
32'd14132: dataIn1 = 32'd452
; 
32'd14133: dataIn1 = 32'd465
; 
32'd14134: dataIn1 = 32'd480
; 
32'd14135: dataIn1 = 32'd517
; 
32'd14136: dataIn1 = 32'd557
; 
32'd14137: dataIn1 = 32'd597
; 
32'd14138: dataIn1 = 32'd599
; 
32'd14139: dataIn1 = 32'd626
; 
32'd14140: dataIn1 = 32'd682
; 
32'd14141: dataIn1 = 32'd728
; 
32'd14142: dataIn1 = 32'd759
; 
32'd14143: dataIn1 = 32'd766
; 
32'd14144: dataIn1 = 32'd776
; 
32'd14145: dataIn1 = 32'd792
; 
32'd14146: dataIn1 = 32'd797
; 
32'd14147: dataIn1 = 32'd190
; 
32'd14148: dataIn1 = 32'd218
; 
32'd14149: dataIn1 = 32'd220
; 
32'd14150: dataIn1 = 32'd243
; 
32'd14151: dataIn1 = 32'd255
; 
32'd14152: dataIn1 = 32'd272
; 
32'd14153: dataIn1 = 32'd281
; 
32'd14154: dataIn1 = 32'd322
; 
32'd14155: dataIn1 = 32'd347
; 
32'd14156: dataIn1 = 32'd350
; 
32'd14157: dataIn1 = 32'd373
; 
32'd14158: dataIn1 = 32'd379
; 
32'd14159: dataIn1 = 32'd388
; 
32'd14160: dataIn1 = 32'd390
; 
32'd14161: dataIn1 = 32'd397
; 
32'd14162: dataIn1 = 32'd402
; 
32'd14163: dataIn1 = 32'd427
; 
32'd14164: dataIn1 = 32'd430
; 
32'd14165: dataIn1 = 32'd498
; 
32'd14166: dataIn1 = 32'd524
; 
32'd14167: dataIn1 = 32'd535
; 
32'd14168: dataIn1 = 32'd549
; 
32'd14169: dataIn1 = 32'd563
; 
32'd14170: dataIn1 = 32'd593
; 
32'd14171: dataIn1 = 32'd614
; 
32'd14172: dataIn1 = 32'd628
; 
32'd14173: dataIn1 = 32'd646
; 
32'd14174: dataIn1 = 32'd655
; 
32'd14175: dataIn1 = 32'd682
; 
32'd14176: dataIn1 = 32'd699
; 
32'd14177: dataIn1 = 32'd700
; 
32'd14178: dataIn1 = 32'd708
; 
32'd14179: dataIn1 = 32'd716
; 
32'd14180: dataIn1 = 32'd720
; 
32'd14181: dataIn1 = 32'd730
; 
32'd14182: dataIn1 = 32'd745
; 
32'd14183: dataIn1 = 32'd756
; 
32'd14184: dataIn1 = 32'd764
; 
32'd14185: dataIn1 = 32'd771
; 
32'd14186: dataIn1 = 32'd780
; 
32'd14187: dataIn1 = 32'd782
; 
32'd14188: dataIn1 = 32'd797
; 
32'd14189: dataIn1 = 32'd800
; 
32'd14190: dataIn1 = 32'd176
; 
32'd14191: dataIn1 = 32'd178
; 
32'd14192: dataIn1 = 32'd181
; 
32'd14193: dataIn1 = 32'd185
; 
32'd14194: dataIn1 = 32'd201
; 
32'd14195: dataIn1 = 32'd206
; 
32'd14196: dataIn1 = 32'd212
; 
32'd14197: dataIn1 = 32'd218
; 
32'd14198: dataIn1 = 32'd225
; 
32'd14199: dataIn1 = 32'd227
; 
32'd14200: dataIn1 = 32'd230
; 
32'd14201: dataIn1 = 32'd246
; 
32'd14202: dataIn1 = 32'd248
; 
32'd14203: dataIn1 = 32'd267
; 
32'd14204: dataIn1 = 32'd272
; 
32'd14205: dataIn1 = 32'd282
; 
32'd14206: dataIn1 = 32'd328
; 
32'd14207: dataIn1 = 32'd342
; 
32'd14208: dataIn1 = 32'd351
; 
32'd14209: dataIn1 = 32'd361
; 
32'd14210: dataIn1 = 32'd373
; 
32'd14211: dataIn1 = 32'd420
; 
32'd14212: dataIn1 = 32'd430
; 
32'd14213: dataIn1 = 32'd438
; 
32'd14214: dataIn1 = 32'd468
; 
32'd14215: dataIn1 = 32'd481
; 
32'd14216: dataIn1 = 32'd482
; 
32'd14217: dataIn1 = 32'd490
; 
32'd14218: dataIn1 = 32'd491
; 
32'd14219: dataIn1 = 32'd494
; 
32'd14220: dataIn1 = 32'd503
; 
32'd14221: dataIn1 = 32'd533
; 
32'd14222: dataIn1 = 32'd536
; 
32'd14223: dataIn1 = 32'd562
; 
32'd14224: dataIn1 = 32'd583
; 
32'd14225: dataIn1 = 32'd588
; 
32'd14226: dataIn1 = 32'd624
; 
32'd14227: dataIn1 = 32'd631
; 
32'd14228: dataIn1 = 32'd638
; 
32'd14229: dataIn1 = 32'd640
; 
32'd14230: dataIn1 = 32'd645
; 
32'd14231: dataIn1 = 32'd649
; 
32'd14232: dataIn1 = 32'd668
; 
32'd14233: dataIn1 = 32'd669
; 
32'd14234: dataIn1 = 32'd675
; 
32'd14235: dataIn1 = 32'd684
; 
32'd14236: dataIn1 = 32'd703
; 
32'd14237: dataIn1 = 32'd708
; 
32'd14238: dataIn1 = 32'd753
; 
32'd14239: dataIn1 = 32'd767
; 
32'd14240: dataIn1 = 32'd790
; 
32'd14241: dataIn1 = 32'd157
; 
32'd14242: dataIn1 = 32'd178
; 
32'd14243: dataIn1 = 32'd188
; 
32'd14244: dataIn1 = 32'd189
; 
32'd14245: dataIn1 = 32'd216
; 
32'd14246: dataIn1 = 32'd222
; 
32'd14247: dataIn1 = 32'd226
; 
32'd14248: dataIn1 = 32'd246
; 
32'd14249: dataIn1 = 32'd252
; 
32'd14250: dataIn1 = 32'd256
; 
32'd14251: dataIn1 = 32'd269
; 
32'd14252: dataIn1 = 32'd293
; 
32'd14253: dataIn1 = 32'd316
; 
32'd14254: dataIn1 = 32'd321
; 
32'd14255: dataIn1 = 32'd326
; 
32'd14256: dataIn1 = 32'd328
; 
32'd14257: dataIn1 = 32'd332
; 
32'd14258: dataIn1 = 32'd353
; 
32'd14259: dataIn1 = 32'd357
; 
32'd14260: dataIn1 = 32'd372
; 
32'd14261: dataIn1 = 32'd374
; 
32'd14262: dataIn1 = 32'd379
; 
32'd14263: dataIn1 = 32'd391
; 
32'd14264: dataIn1 = 32'd425
; 
32'd14265: dataIn1 = 32'd441
; 
32'd14266: dataIn1 = 32'd454
; 
32'd14267: dataIn1 = 32'd461
; 
32'd14268: dataIn1 = 32'd469
; 
32'd14269: dataIn1 = 32'd502
; 
32'd14270: dataIn1 = 32'd503
; 
32'd14271: dataIn1 = 32'd520
; 
32'd14272: dataIn1 = 32'd534
; 
32'd14273: dataIn1 = 32'd563
; 
32'd14274: dataIn1 = 32'd569
; 
32'd14275: dataIn1 = 32'd585
; 
32'd14276: dataIn1 = 32'd587
; 
32'd14277: dataIn1 = 32'd615
; 
32'd14278: dataIn1 = 32'd619
; 
32'd14279: dataIn1 = 32'd625
; 
32'd14280: dataIn1 = 32'd630
; 
32'd14281: dataIn1 = 32'd634
; 
32'd14282: dataIn1 = 32'd645
; 
32'd14283: dataIn1 = 32'd696
; 
32'd14284: dataIn1 = 32'd738
; 
32'd14285: dataIn1 = 32'd744
; 
32'd14286: dataIn1 = 32'd755
; 
32'd14287: dataIn1 = 32'd762
; 
32'd14288: dataIn1 = 32'd778
; 
32'd14289: dataIn1 = 32'd787
; 
32'd14290: dataIn1 = 32'd794
; 
32'd14291: dataIn1 = 32'd795
; 
32'd14292: dataIn1 = 32'd796
; 
32'd14293: dataIn1 = 32'd148
; 
32'd14294: dataIn1 = 32'd156
; 
32'd14295: dataIn1 = 32'd164
; 
32'd14296: dataIn1 = 32'd165
; 
32'd14297: dataIn1 = 32'd176
; 
32'd14298: dataIn1 = 32'd178
; 
32'd14299: dataIn1 = 32'd181
; 
32'd14300: dataIn1 = 32'd186
; 
32'd14301: dataIn1 = 32'd194
; 
32'd14302: dataIn1 = 32'd214
; 
32'd14303: dataIn1 = 32'd223
; 
32'd14304: dataIn1 = 32'd235
; 
32'd14305: dataIn1 = 32'd259
; 
32'd14306: dataIn1 = 32'd267
; 
32'd14307: dataIn1 = 32'd335
; 
32'd14308: dataIn1 = 32'd352
; 
32'd14309: dataIn1 = 32'd353
; 
32'd14310: dataIn1 = 32'd388
; 
32'd14311: dataIn1 = 32'd398
; 
32'd14312: dataIn1 = 32'd418
; 
32'd14313: dataIn1 = 32'd429
; 
32'd14314: dataIn1 = 32'd442
; 
32'd14315: dataIn1 = 32'd455
; 
32'd14316: dataIn1 = 32'd462
; 
32'd14317: dataIn1 = 32'd480
; 
32'd14318: dataIn1 = 32'd489
; 
32'd14319: dataIn1 = 32'd503
; 
32'd14320: dataIn1 = 32'd515
; 
32'd14321: dataIn1 = 32'd529
; 
32'd14322: dataIn1 = 32'd539
; 
32'd14323: dataIn1 = 32'd542
; 
32'd14324: dataIn1 = 32'd546
; 
32'd14325: dataIn1 = 32'd587
; 
32'd14326: dataIn1 = 32'd589
; 
32'd14327: dataIn1 = 32'd593
; 
32'd14328: dataIn1 = 32'd600
; 
32'd14329: dataIn1 = 32'd646
; 
32'd14330: dataIn1 = 32'd655
; 
32'd14331: dataIn1 = 32'd671
; 
32'd14332: dataIn1 = 32'd713
; 
32'd14333: dataIn1 = 32'd726
; 
32'd14334: dataIn1 = 32'd728
; 
32'd14335: dataIn1 = 32'd784
; 
32'd14336: dataIn1 = 32'd790
; 
32'd14337: dataIn1 = 32'd176
; 
32'd14338: dataIn1 = 32'd200
; 
32'd14339: dataIn1 = 32'd203
; 
32'd14340: dataIn1 = 32'd204
; 
32'd14341: dataIn1 = 32'd215
; 
32'd14342: dataIn1 = 32'd223
; 
32'd14343: dataIn1 = 32'd257
; 
32'd14344: dataIn1 = 32'd258
; 
32'd14345: dataIn1 = 32'd279
; 
32'd14346: dataIn1 = 32'd285
; 
32'd14347: dataIn1 = 32'd300
; 
32'd14348: dataIn1 = 32'd339
; 
32'd14349: dataIn1 = 32'd371
; 
32'd14350: dataIn1 = 32'd393
; 
32'd14351: dataIn1 = 32'd396
; 
32'd14352: dataIn1 = 32'd448
; 
32'd14353: dataIn1 = 32'd450
; 
32'd14354: dataIn1 = 32'd483
; 
32'd14355: dataIn1 = 32'd510
; 
32'd14356: dataIn1 = 32'd515
; 
32'd14357: dataIn1 = 32'd531
; 
32'd14358: dataIn1 = 32'd537
; 
32'd14359: dataIn1 = 32'd575
; 
32'd14360: dataIn1 = 32'd578
; 
32'd14361: dataIn1 = 32'd579
; 
32'd14362: dataIn1 = 32'd580
; 
32'd14363: dataIn1 = 32'd589
; 
32'd14364: dataIn1 = 32'd611
; 
32'd14365: dataIn1 = 32'd634
; 
32'd14366: dataIn1 = 32'd654
; 
32'd14367: dataIn1 = 32'd664
; 
32'd14368: dataIn1 = 32'd666
; 
32'd14369: dataIn1 = 32'd674
; 
32'd14370: dataIn1 = 32'd717
; 
32'd14371: dataIn1 = 32'd718
; 
32'd14372: dataIn1 = 32'd752
; 
32'd14373: dataIn1 = 32'd765
; 
32'd14374: dataIn1 = 32'd158
; 
32'd14375: dataIn1 = 32'd174
; 
32'd14376: dataIn1 = 32'd196
; 
32'd14377: dataIn1 = 32'd216
; 
32'd14378: dataIn1 = 32'd223
; 
32'd14379: dataIn1 = 32'd232
; 
32'd14380: dataIn1 = 32'd234
; 
32'd14381: dataIn1 = 32'd238
; 
32'd14382: dataIn1 = 32'd247
; 
32'd14383: dataIn1 = 32'd256
; 
32'd14384: dataIn1 = 32'd285
; 
32'd14385: dataIn1 = 32'd315
; 
32'd14386: dataIn1 = 32'd339
; 
32'd14387: dataIn1 = 32'd341
; 
32'd14388: dataIn1 = 32'd346
; 
32'd14389: dataIn1 = 32'd353
; 
32'd14390: dataIn1 = 32'd359
; 
32'd14391: dataIn1 = 32'd360
; 
32'd14392: dataIn1 = 32'd391
; 
32'd14393: dataIn1 = 32'd475
; 
32'd14394: dataIn1 = 32'd485
; 
32'd14395: dataIn1 = 32'd508
; 
32'd14396: dataIn1 = 32'd510
; 
32'd14397: dataIn1 = 32'd533
; 
32'd14398: dataIn1 = 32'd543
; 
32'd14399: dataIn1 = 32'd553
; 
32'd14400: dataIn1 = 32'd597
; 
32'd14401: dataIn1 = 32'd604
; 
32'd14402: dataIn1 = 32'd610
; 
32'd14403: dataIn1 = 32'd636
; 
32'd14404: dataIn1 = 32'd639
; 
32'd14405: dataIn1 = 32'd641
; 
32'd14406: dataIn1 = 32'd666
; 
32'd14407: dataIn1 = 32'd674
; 
32'd14408: dataIn1 = 32'd704
; 
32'd14409: dataIn1 = 32'd724
; 
32'd14410: dataIn1 = 32'd732
; 
32'd14411: dataIn1 = 32'd738
; 
32'd14412: dataIn1 = 32'd740
; 
32'd14413: dataIn1 = 32'd773
; 
32'd14414: dataIn1 = 32'd791
; 
32'd14415: dataIn1 = 32'd793
; 
32'd14416: dataIn1 = 32'd799
; 
32'd14417: dataIn1 = 32'd161
; 
32'd14418: dataIn1 = 32'd167
; 
32'd14419: dataIn1 = 32'd169
; 
32'd14420: dataIn1 = 32'd183
; 
32'd14421: dataIn1 = 32'd187
; 
32'd14422: dataIn1 = 32'd222
; 
32'd14423: dataIn1 = 32'd237
; 
32'd14424: dataIn1 = 32'd251
; 
32'd14425: dataIn1 = 32'd256
; 
32'd14426: dataIn1 = 32'd311
; 
32'd14427: dataIn1 = 32'd344
; 
32'd14428: dataIn1 = 32'd365
; 
32'd14429: dataIn1 = 32'd368
; 
32'd14430: dataIn1 = 32'd370
; 
32'd14431: dataIn1 = 32'd396
; 
32'd14432: dataIn1 = 32'd412
; 
32'd14433: dataIn1 = 32'd445
; 
32'd14434: dataIn1 = 32'd471
; 
32'd14435: dataIn1 = 32'd486
; 
32'd14436: dataIn1 = 32'd522
; 
32'd14437: dataIn1 = 32'd545
; 
32'd14438: dataIn1 = 32'd546
; 
32'd14439: dataIn1 = 32'd580
; 
32'd14440: dataIn1 = 32'd584
; 
32'd14441: dataIn1 = 32'd594
; 
32'd14442: dataIn1 = 32'd599
; 
32'd14443: dataIn1 = 32'd603
; 
32'd14444: dataIn1 = 32'd607
; 
32'd14445: dataIn1 = 32'd649
; 
32'd14446: dataIn1 = 32'd674
; 
32'd14447: dataIn1 = 32'd676
; 
32'd14448: dataIn1 = 32'd684
; 
32'd14449: dataIn1 = 32'd725
; 
32'd14450: dataIn1 = 32'd729
; 
32'd14451: dataIn1 = 32'd777
; 
32'd14452: dataIn1 = 32'd787
; 
32'd14453: dataIn1 = 32'd177
; 
32'd14454: dataIn1 = 32'd179
; 
32'd14455: dataIn1 = 32'd193
; 
32'd14456: dataIn1 = 32'd199
; 
32'd14457: dataIn1 = 32'd202
; 
32'd14458: dataIn1 = 32'd233
; 
32'd14459: dataIn1 = 32'd250
; 
32'd14460: dataIn1 = 32'd265
; 
32'd14461: dataIn1 = 32'd271
; 
32'd14462: dataIn1 = 32'd308
; 
32'd14463: dataIn1 = 32'd314
; 
32'd14464: dataIn1 = 32'd329
; 
32'd14465: dataIn1 = 32'd349
; 
32'd14466: dataIn1 = 32'd367
; 
32'd14467: dataIn1 = 32'd372
; 
32'd14468: dataIn1 = 32'd389
; 
32'd14469: dataIn1 = 32'd400
; 
32'd14470: dataIn1 = 32'd409
; 
32'd14471: dataIn1 = 32'd420
; 
32'd14472: dataIn1 = 32'd435
; 
32'd14473: dataIn1 = 32'd448
; 
32'd14474: dataIn1 = 32'd449
; 
32'd14475: dataIn1 = 32'd454
; 
32'd14476: dataIn1 = 32'd455
; 
32'd14477: dataIn1 = 32'd460
; 
32'd14478: dataIn1 = 32'd465
; 
32'd14479: dataIn1 = 32'd494
; 
32'd14480: dataIn1 = 32'd495
; 
32'd14481: dataIn1 = 32'd521
; 
32'd14482: dataIn1 = 32'd575
; 
32'd14483: dataIn1 = 32'd584
; 
32'd14484: dataIn1 = 32'd609
; 
32'd14485: dataIn1 = 32'd619
; 
32'd14486: dataIn1 = 32'd650
; 
32'd14487: dataIn1 = 32'd659
; 
32'd14488: dataIn1 = 32'd688
; 
32'd14489: dataIn1 = 32'd697
; 
32'd14490: dataIn1 = 32'd707
; 
32'd14491: dataIn1 = 32'd708
; 
32'd14492: dataIn1 = 32'd710
; 
32'd14493: dataIn1 = 32'd755
; 
32'd14494: dataIn1 = 32'd766
; 
32'd14495: dataIn1 = 32'd791
; 
32'd14496: dataIn1 = 32'd154
; 
32'd14497: dataIn1 = 32'd182
; 
32'd14498: dataIn1 = 32'd191
; 
32'd14499: dataIn1 = 32'd260
; 
32'd14500: dataIn1 = 32'd263
; 
32'd14501: dataIn1 = 32'd288
; 
32'd14502: dataIn1 = 32'd302
; 
32'd14503: dataIn1 = 32'd315
; 
32'd14504: dataIn1 = 32'd331
; 
32'd14505: dataIn1 = 32'd338
; 
32'd14506: dataIn1 = 32'd399
; 
32'd14507: dataIn1 = 32'd418
; 
32'd14508: dataIn1 = 32'd423
; 
32'd14509: dataIn1 = 32'd438
; 
32'd14510: dataIn1 = 32'd448
; 
32'd14511: dataIn1 = 32'd456
; 
32'd14512: dataIn1 = 32'd458
; 
32'd14513: dataIn1 = 32'd490
; 
32'd14514: dataIn1 = 32'd510
; 
32'd14515: dataIn1 = 32'd514
; 
32'd14516: dataIn1 = 32'd525
; 
32'd14517: dataIn1 = 32'd526
; 
32'd14518: dataIn1 = 32'd540
; 
32'd14519: dataIn1 = 32'd562
; 
32'd14520: dataIn1 = 32'd563
; 
32'd14521: dataIn1 = 32'd602
; 
32'd14522: dataIn1 = 32'd616
; 
32'd14523: dataIn1 = 32'd712
; 
32'd14524: dataIn1 = 32'd744
; 
32'd14525: dataIn1 = 32'd790
; 
32'd14526: dataIn1 = 32'd798
; 
32'd14527: dataIn1 = 32'd159
; 
32'd14528: dataIn1 = 32'd161
; 
32'd14529: dataIn1 = 32'd168
; 
32'd14530: dataIn1 = 32'd172
; 
32'd14531: dataIn1 = 32'd207
; 
32'd14532: dataIn1 = 32'd224
; 
32'd14533: dataIn1 = 32'd240
; 
32'd14534: dataIn1 = 32'd255
; 
32'd14535: dataIn1 = 32'd271
; 
32'd14536: dataIn1 = 32'd275
; 
32'd14537: dataIn1 = 32'd290
; 
32'd14538: dataIn1 = 32'd320
; 
32'd14539: dataIn1 = 32'd328
; 
32'd14540: dataIn1 = 32'd342
; 
32'd14541: dataIn1 = 32'd376
; 
32'd14542: dataIn1 = 32'd384
; 
32'd14543: dataIn1 = 32'd420
; 
32'd14544: dataIn1 = 32'd436
; 
32'd14545: dataIn1 = 32'd439
; 
32'd14546: dataIn1 = 32'd472
; 
32'd14547: dataIn1 = 32'd474
; 
32'd14548: dataIn1 = 32'd481
; 
32'd14549: dataIn1 = 32'd489
; 
32'd14550: dataIn1 = 32'd563
; 
32'd14551: dataIn1 = 32'd564
; 
32'd14552: dataIn1 = 32'd576
; 
32'd14553: dataIn1 = 32'd616
; 
32'd14554: dataIn1 = 32'd627
; 
32'd14555: dataIn1 = 32'd636
; 
32'd14556: dataIn1 = 32'd681
; 
32'd14557: dataIn1 = 32'd692
; 
32'd14558: dataIn1 = 32'd693
; 
32'd14559: dataIn1 = 32'd695
; 
32'd14560: dataIn1 = 32'd703
; 
32'd14561: dataIn1 = 32'd712
; 
32'd14562: dataIn1 = 32'd713
; 
32'd14563: dataIn1 = 32'd727
; 
32'd14564: dataIn1 = 32'd728
; 
32'd14565: dataIn1 = 32'd758
; 
32'd14566: dataIn1 = 32'd765
; 
32'd14567: dataIn1 = 32'd773
; 
32'd14568: dataIn1 = 32'd781
; 
32'd14569: dataIn1 = 32'd160
; 
32'd14570: dataIn1 = 32'd161
; 
32'd14571: dataIn1 = 32'd177
; 
32'd14572: dataIn1 = 32'd201
; 
32'd14573: dataIn1 = 32'd235
; 
32'd14574: dataIn1 = 32'd272
; 
32'd14575: dataIn1 = 32'd282
; 
32'd14576: dataIn1 = 32'd291
; 
32'd14577: dataIn1 = 32'd298
; 
32'd14578: dataIn1 = 32'd363
; 
32'd14579: dataIn1 = 32'd392
; 
32'd14580: dataIn1 = 32'd397
; 
32'd14581: dataIn1 = 32'd424
; 
32'd14582: dataIn1 = 32'd425
; 
32'd14583: dataIn1 = 32'd427
; 
32'd14584: dataIn1 = 32'd433
; 
32'd14585: dataIn1 = 32'd451
; 
32'd14586: dataIn1 = 32'd489
; 
32'd14587: dataIn1 = 32'd492
; 
32'd14588: dataIn1 = 32'd495
; 
32'd14589: dataIn1 = 32'd501
; 
32'd14590: dataIn1 = 32'd507
; 
32'd14591: dataIn1 = 32'd547
; 
32'd14592: dataIn1 = 32'd568
; 
32'd14593: dataIn1 = 32'd589
; 
32'd14594: dataIn1 = 32'd605
; 
32'd14595: dataIn1 = 32'd610
; 
32'd14596: dataIn1 = 32'd618
; 
32'd14597: dataIn1 = 32'd634
; 
32'd14598: dataIn1 = 32'd652
; 
32'd14599: dataIn1 = 32'd679
; 
32'd14600: dataIn1 = 32'd685
; 
32'd14601: dataIn1 = 32'd687
; 
32'd14602: dataIn1 = 32'd700
; 
32'd14603: dataIn1 = 32'd721
; 
32'd14604: dataIn1 = 32'd741
; 
32'd14605: dataIn1 = 32'd187
; 
32'd14606: dataIn1 = 32'd210
; 
32'd14607: dataIn1 = 32'd211
; 
32'd14608: dataIn1 = 32'd213
; 
32'd14609: dataIn1 = 32'd217
; 
32'd14610: dataIn1 = 32'd243
; 
32'd14611: dataIn1 = 32'd245
; 
32'd14612: dataIn1 = 32'd254
; 
32'd14613: dataIn1 = 32'd269
; 
32'd14614: dataIn1 = 32'd293
; 
32'd14615: dataIn1 = 32'd297
; 
32'd14616: dataIn1 = 32'd300
; 
32'd14617: dataIn1 = 32'd346
; 
32'd14618: dataIn1 = 32'd354
; 
32'd14619: dataIn1 = 32'd358
; 
32'd14620: dataIn1 = 32'd362
; 
32'd14621: dataIn1 = 32'd384
; 
32'd14622: dataIn1 = 32'd395
; 
32'd14623: dataIn1 = 32'd445
; 
32'd14624: dataIn1 = 32'd456
; 
32'd14625: dataIn1 = 32'd461
; 
32'd14626: dataIn1 = 32'd463
; 
32'd14627: dataIn1 = 32'd478
; 
32'd14628: dataIn1 = 32'd500
; 
32'd14629: dataIn1 = 32'd504
; 
32'd14630: dataIn1 = 32'd510
; 
32'd14631: dataIn1 = 32'd517
; 
32'd14632: dataIn1 = 32'd552
; 
32'd14633: dataIn1 = 32'd565
; 
32'd14634: dataIn1 = 32'd585
; 
32'd14635: dataIn1 = 32'd591
; 
32'd14636: dataIn1 = 32'd622
; 
32'd14637: dataIn1 = 32'd651
; 
32'd14638: dataIn1 = 32'd670
; 
32'd14639: dataIn1 = 32'd693
; 
32'd14640: dataIn1 = 32'd717
; 
32'd14641: dataIn1 = 32'd724
; 
32'd14642: dataIn1 = 32'd739
; 
32'd14643: dataIn1 = 32'd745
; 
32'd14644: dataIn1 = 32'd760
; 
32'd14645: dataIn1 = 32'd798
; 
32'd14646: dataIn1 = 32'd212
; 
32'd14647: dataIn1 = 32'd243
; 
32'd14648: dataIn1 = 32'd276
; 
32'd14649: dataIn1 = 32'd297
; 
32'd14650: dataIn1 = 32'd326
; 
32'd14651: dataIn1 = 32'd338
; 
32'd14652: dataIn1 = 32'd346
; 
32'd14653: dataIn1 = 32'd366
; 
32'd14654: dataIn1 = 32'd367
; 
32'd14655: dataIn1 = 32'd420
; 
32'd14656: dataIn1 = 32'd425
; 
32'd14657: dataIn1 = 32'd458
; 
32'd14658: dataIn1 = 32'd529
; 
32'd14659: dataIn1 = 32'd534
; 
32'd14660: dataIn1 = 32'd567
; 
32'd14661: dataIn1 = 32'd584
; 
32'd14662: dataIn1 = 32'd596
; 
32'd14663: dataIn1 = 32'd609
; 
32'd14664: dataIn1 = 32'd610
; 
32'd14665: dataIn1 = 32'd614
; 
32'd14666: dataIn1 = 32'd615
; 
32'd14667: dataIn1 = 32'd647
; 
32'd14668: dataIn1 = 32'd674
; 
32'd14669: dataIn1 = 32'd695
; 
32'd14670: dataIn1 = 32'd727
; 
32'd14671: dataIn1 = 32'd744
; 
32'd14672: dataIn1 = 32'd761
; 
32'd14673: dataIn1 = 32'd766
; 
32'd14674: dataIn1 = 32'd785
; 
32'd14675: dataIn1 = 32'd788
; 
32'd14676: dataIn1 = 32'd792
; 
32'd14677: dataIn1 = 32'd796
; 
32'd14678: dataIn1 = 32'd159
; 
32'd14679: dataIn1 = 32'd193
; 
32'd14680: dataIn1 = 32'd200
; 
32'd14681: dataIn1 = 32'd214
; 
32'd14682: dataIn1 = 32'd215
; 
32'd14683: dataIn1 = 32'd270
; 
32'd14684: dataIn1 = 32'd282
; 
32'd14685: dataIn1 = 32'd312
; 
32'd14686: dataIn1 = 32'd323
; 
32'd14687: dataIn1 = 32'd341
; 
32'd14688: dataIn1 = 32'd370
; 
32'd14689: dataIn1 = 32'd384
; 
32'd14690: dataIn1 = 32'd385
; 
32'd14691: dataIn1 = 32'd417
; 
32'd14692: dataIn1 = 32'd426
; 
32'd14693: dataIn1 = 32'd445
; 
32'd14694: dataIn1 = 32'd468
; 
32'd14695: dataIn1 = 32'd476
; 
32'd14696: dataIn1 = 32'd478
; 
32'd14697: dataIn1 = 32'd480
; 
32'd14698: dataIn1 = 32'd481
; 
32'd14699: dataIn1 = 32'd508
; 
32'd14700: dataIn1 = 32'd515
; 
32'd14701: dataIn1 = 32'd516
; 
32'd14702: dataIn1 = 32'd567
; 
32'd14703: dataIn1 = 32'd572
; 
32'd14704: dataIn1 = 32'd578
; 
32'd14705: dataIn1 = 32'd593
; 
32'd14706: dataIn1 = 32'd624
; 
32'd14707: dataIn1 = 32'd669
; 
32'd14708: dataIn1 = 32'd680
; 
32'd14709: dataIn1 = 32'd683
; 
32'd14710: dataIn1 = 32'd694
; 
32'd14711: dataIn1 = 32'd706
; 
32'd14712: dataIn1 = 32'd740
; 
32'd14713: dataIn1 = 32'd770
; 
32'd14714: dataIn1 = 32'd789
; 
32'd14715: dataIn1 = 32'd790
; 
32'd14716: dataIn1 = 32'd210
; 
32'd14717: dataIn1 = 32'd235
; 
32'd14718: dataIn1 = 32'd260
; 
32'd14719: dataIn1 = 32'd293
; 
32'd14720: dataIn1 = 32'd296
; 
32'd14721: dataIn1 = 32'd317
; 
32'd14722: dataIn1 = 32'd341
; 
32'd14723: dataIn1 = 32'd353
; 
32'd14724: dataIn1 = 32'd362
; 
32'd14725: dataIn1 = 32'd369
; 
32'd14726: dataIn1 = 32'd392
; 
32'd14727: dataIn1 = 32'd411
; 
32'd14728: dataIn1 = 32'd423
; 
32'd14729: dataIn1 = 32'd498
; 
32'd14730: dataIn1 = 32'd500
; 
32'd14731: dataIn1 = 32'd505
; 
32'd14732: dataIn1 = 32'd508
; 
32'd14733: dataIn1 = 32'd511
; 
32'd14734: dataIn1 = 32'd518
; 
32'd14735: dataIn1 = 32'd528
; 
32'd14736: dataIn1 = 32'd529
; 
32'd14737: dataIn1 = 32'd555
; 
32'd14738: dataIn1 = 32'd559
; 
32'd14739: dataIn1 = 32'd569
; 
32'd14740: dataIn1 = 32'd573
; 
32'd14741: dataIn1 = 32'd575
; 
32'd14742: dataIn1 = 32'd579
; 
32'd14743: dataIn1 = 32'd581
; 
32'd14744: dataIn1 = 32'd587
; 
32'd14745: dataIn1 = 32'd589
; 
32'd14746: dataIn1 = 32'd607
; 
32'd14747: dataIn1 = 32'd615
; 
32'd14748: dataIn1 = 32'd627
; 
32'd14749: dataIn1 = 32'd672
; 
32'd14750: dataIn1 = 32'd673
; 
32'd14751: dataIn1 = 32'd700
; 
32'd14752: dataIn1 = 32'd705
; 
32'd14753: dataIn1 = 32'd732
; 
32'd14754: dataIn1 = 32'd733
; 
32'd14755: dataIn1 = 32'd761
; 
32'd14756: dataIn1 = 32'd766
; 
32'd14757: dataIn1 = 32'd793
; 
32'd14758: dataIn1 = 32'd796
; 
32'd14759: dataIn1 = 32'd171
; 
32'd14760: dataIn1 = 32'd192
; 
32'd14761: dataIn1 = 32'd220
; 
32'd14762: dataIn1 = 32'd246
; 
32'd14763: dataIn1 = 32'd279
; 
32'd14764: dataIn1 = 32'd295
; 
32'd14765: dataIn1 = 32'd338
; 
32'd14766: dataIn1 = 32'd344
; 
32'd14767: dataIn1 = 32'd353
; 
32'd14768: dataIn1 = 32'd357
; 
32'd14769: dataIn1 = 32'd380
; 
32'd14770: dataIn1 = 32'd396
; 
32'd14771: dataIn1 = 32'd397
; 
32'd14772: dataIn1 = 32'd399
; 
32'd14773: dataIn1 = 32'd417
; 
32'd14774: dataIn1 = 32'd428
; 
32'd14775: dataIn1 = 32'd473
; 
32'd14776: dataIn1 = 32'd496
; 
32'd14777: dataIn1 = 32'd514
; 
32'd14778: dataIn1 = 32'd517
; 
32'd14779: dataIn1 = 32'd572
; 
32'd14780: dataIn1 = 32'd597
; 
32'd14781: dataIn1 = 32'd641
; 
32'd14782: dataIn1 = 32'd651
; 
32'd14783: dataIn1 = 32'd655
; 
32'd14784: dataIn1 = 32'd656
; 
32'd14785: dataIn1 = 32'd671
; 
32'd14786: dataIn1 = 32'd677
; 
32'd14787: dataIn1 = 32'd681
; 
32'd14788: dataIn1 = 32'd716
; 
32'd14789: dataIn1 = 32'd719
; 
32'd14790: dataIn1 = 32'd724
; 
32'd14791: dataIn1 = 32'd736
; 
32'd14792: dataIn1 = 32'd767
; 
32'd14793: dataIn1 = 32'd772
; 
32'd14794: dataIn1 = 32'd774
; 
32'd14795: dataIn1 = 32'd795
; 
32'd14796: dataIn1 = 32'd797
; 
32'd14797: dataIn1 = 32'd216
; 
32'd14798: dataIn1 = 32'd240
; 
32'd14799: dataIn1 = 32'd245
; 
32'd14800: dataIn1 = 32'd249
; 
32'd14801: dataIn1 = 32'd271
; 
32'd14802: dataIn1 = 32'd272
; 
32'd14803: dataIn1 = 32'd288
; 
32'd14804: dataIn1 = 32'd345
; 
32'd14805: dataIn1 = 32'd348
; 
32'd14806: dataIn1 = 32'd364
; 
32'd14807: dataIn1 = 32'd392
; 
32'd14808: dataIn1 = 32'd395
; 
32'd14809: dataIn1 = 32'd413
; 
32'd14810: dataIn1 = 32'd432
; 
32'd14811: dataIn1 = 32'd442
; 
32'd14812: dataIn1 = 32'd462
; 
32'd14813: dataIn1 = 32'd495
; 
32'd14814: dataIn1 = 32'd509
; 
32'd14815: dataIn1 = 32'd533
; 
32'd14816: dataIn1 = 32'd543
; 
32'd14817: dataIn1 = 32'd560
; 
32'd14818: dataIn1 = 32'd577
; 
32'd14819: dataIn1 = 32'd581
; 
32'd14820: dataIn1 = 32'd613
; 
32'd14821: dataIn1 = 32'd614
; 
32'd14822: dataIn1 = 32'd624
; 
32'd14823: dataIn1 = 32'd669
; 
32'd14824: dataIn1 = 32'd698
; 
32'd14825: dataIn1 = 32'd734
; 
32'd14826: dataIn1 = 32'd742
; 
32'd14827: dataIn1 = 32'd767
; 
32'd14828: dataIn1 = 32'd776
; 
32'd14829: dataIn1 = 32'd779
; 
32'd14830: dataIn1 = 32'd787
; 
32'd14831: dataIn1 = 32'd188
; 
32'd14832: dataIn1 = 32'd197
; 
32'd14833: dataIn1 = 32'd213
; 
32'd14834: dataIn1 = 32'd215
; 
32'd14835: dataIn1 = 32'd253
; 
32'd14836: dataIn1 = 32'd285
; 
32'd14837: dataIn1 = 32'd306
; 
32'd14838: dataIn1 = 32'd344
; 
32'd14839: dataIn1 = 32'd353
; 
32'd14840: dataIn1 = 32'd371
; 
32'd14841: dataIn1 = 32'd380
; 
32'd14842: dataIn1 = 32'd406
; 
32'd14843: dataIn1 = 32'd412
; 
32'd14844: dataIn1 = 32'd460
; 
32'd14845: dataIn1 = 32'd466
; 
32'd14846: dataIn1 = 32'd512
; 
32'd14847: dataIn1 = 32'd516
; 
32'd14848: dataIn1 = 32'd528
; 
32'd14849: dataIn1 = 32'd539
; 
32'd14850: dataIn1 = 32'd567
; 
32'd14851: dataIn1 = 32'd573
; 
32'd14852: dataIn1 = 32'd587
; 
32'd14853: dataIn1 = 32'd590
; 
32'd14854: dataIn1 = 32'd591
; 
32'd14855: dataIn1 = 32'd604
; 
32'd14856: dataIn1 = 32'd616
; 
32'd14857: dataIn1 = 32'd621
; 
32'd14858: dataIn1 = 32'd623
; 
32'd14859: dataIn1 = 32'd646
; 
32'd14860: dataIn1 = 32'd668
; 
32'd14861: dataIn1 = 32'd678
; 
32'd14862: dataIn1 = 32'd701
; 
32'd14863: dataIn1 = 32'd741
; 
32'd14864: dataIn1 = 32'd743
; 
32'd14865: dataIn1 = 32'd745
; 
32'd14866: dataIn1 = 32'd751
; 
32'd14867: dataIn1 = 32'd763
; 
32'd14868: dataIn1 = 32'd770
; 
32'd14869: dataIn1 = 32'd774
; 
32'd14870: dataIn1 = 32'd778
; 
32'd14871: dataIn1 = 32'd780
; 
32'd14872: dataIn1 = 32'd171
; 
32'd14873: dataIn1 = 32'd215
; 
32'd14874: dataIn1 = 32'd221
; 
32'd14875: dataIn1 = 32'd279
; 
32'd14876: dataIn1 = 32'd297
; 
32'd14877: dataIn1 = 32'd310
; 
32'd14878: dataIn1 = 32'd313
; 
32'd14879: dataIn1 = 32'd329
; 
32'd14880: dataIn1 = 32'd339
; 
32'd14881: dataIn1 = 32'd361
; 
32'd14882: dataIn1 = 32'd438
; 
32'd14883: dataIn1 = 32'd440
; 
32'd14884: dataIn1 = 32'd451
; 
32'd14885: dataIn1 = 32'd461
; 
32'd14886: dataIn1 = 32'd485
; 
32'd14887: dataIn1 = 32'd516
; 
32'd14888: dataIn1 = 32'd520
; 
32'd14889: dataIn1 = 32'd525
; 
32'd14890: dataIn1 = 32'd533
; 
32'd14891: dataIn1 = 32'd536
; 
32'd14892: dataIn1 = 32'd537
; 
32'd14893: dataIn1 = 32'd563
; 
32'd14894: dataIn1 = 32'd572
; 
32'd14895: dataIn1 = 32'd595
; 
32'd14896: dataIn1 = 32'd596
; 
32'd14897: dataIn1 = 32'd615
; 
32'd14898: dataIn1 = 32'd632
; 
32'd14899: dataIn1 = 32'd663
; 
32'd14900: dataIn1 = 32'd669
; 
32'd14901: dataIn1 = 32'd695
; 
32'd14902: dataIn1 = 32'd699
; 
32'd14903: dataIn1 = 32'd719
; 
32'd14904: dataIn1 = 32'd780
; 
32'd14905: dataIn1 = 32'd797
; 
32'd14906: dataIn1 = 32'd175
; 
32'd14907: dataIn1 = 32'd178
; 
32'd14908: dataIn1 = 32'd191
; 
32'd14909: dataIn1 = 32'd193
; 
32'd14910: dataIn1 = 32'd208
; 
32'd14911: dataIn1 = 32'd214
; 
32'd14912: dataIn1 = 32'd261
; 
32'd14913: dataIn1 = 32'd273
; 
32'd14914: dataIn1 = 32'd281
; 
32'd14915: dataIn1 = 32'd291
; 
32'd14916: dataIn1 = 32'd295
; 
32'd14917: dataIn1 = 32'd336
; 
32'd14918: dataIn1 = 32'd342
; 
32'd14919: dataIn1 = 32'd343
; 
32'd14920: dataIn1 = 32'd344
; 
32'd14921: dataIn1 = 32'd363
; 
32'd14922: dataIn1 = 32'd372
; 
32'd14923: dataIn1 = 32'd387
; 
32'd14924: dataIn1 = 32'd389
; 
32'd14925: dataIn1 = 32'd391
; 
32'd14926: dataIn1 = 32'd403
; 
32'd14927: dataIn1 = 32'd404
; 
32'd14928: dataIn1 = 32'd421
; 
32'd14929: dataIn1 = 32'd438
; 
32'd14930: dataIn1 = 32'd439
; 
32'd14931: dataIn1 = 32'd445
; 
32'd14932: dataIn1 = 32'd454
; 
32'd14933: dataIn1 = 32'd475
; 
32'd14934: dataIn1 = 32'd497
; 
32'd14935: dataIn1 = 32'd500
; 
32'd14936: dataIn1 = 32'd536
; 
32'd14937: dataIn1 = 32'd578
; 
32'd14938: dataIn1 = 32'd595
; 
32'd14939: dataIn1 = 32'd603
; 
32'd14940: dataIn1 = 32'd604
; 
32'd14941: dataIn1 = 32'd608
; 
32'd14942: dataIn1 = 32'd612
; 
32'd14943: dataIn1 = 32'd628
; 
32'd14944: dataIn1 = 32'd646
; 
32'd14945: dataIn1 = 32'd653
; 
32'd14946: dataIn1 = 32'd665
; 
32'd14947: dataIn1 = 32'd668
; 
32'd14948: dataIn1 = 32'd679
; 
32'd14949: dataIn1 = 32'd686
; 
32'd14950: dataIn1 = 32'd689
; 
32'd14951: dataIn1 = 32'd705
; 
32'd14952: dataIn1 = 32'd733
; 
32'd14953: dataIn1 = 32'd759
; 
32'd14954: dataIn1 = 32'd776
; 
32'd14955: dataIn1 = 32'd778
; 
32'd14956: dataIn1 = 32'd788
; 
32'd14957: dataIn1 = 32'd225
; 
32'd14958: dataIn1 = 32'd227
; 
32'd14959: dataIn1 = 32'd228
; 
32'd14960: dataIn1 = 32'd238
; 
32'd14961: dataIn1 = 32'd243
; 
32'd14962: dataIn1 = 32'd246
; 
32'd14963: dataIn1 = 32'd254
; 
32'd14964: dataIn1 = 32'd264
; 
32'd14965: dataIn1 = 32'd304
; 
32'd14966: dataIn1 = 32'd330
; 
32'd14967: dataIn1 = 32'd336
; 
32'd14968: dataIn1 = 32'd350
; 
32'd14969: dataIn1 = 32'd353
; 
32'd14970: dataIn1 = 32'd358
; 
32'd14971: dataIn1 = 32'd368
; 
32'd14972: dataIn1 = 32'd376
; 
32'd14973: dataIn1 = 32'd393
; 
32'd14974: dataIn1 = 32'd433
; 
32'd14975: dataIn1 = 32'd442
; 
32'd14976: dataIn1 = 32'd456
; 
32'd14977: dataIn1 = 32'd470
; 
32'd14978: dataIn1 = 32'd472
; 
32'd14979: dataIn1 = 32'd476
; 
32'd14980: dataIn1 = 32'd482
; 
32'd14981: dataIn1 = 32'd517
; 
32'd14982: dataIn1 = 32'd526
; 
32'd14983: dataIn1 = 32'd531
; 
32'd14984: dataIn1 = 32'd539
; 
32'd14985: dataIn1 = 32'd555
; 
32'd14986: dataIn1 = 32'd594
; 
32'd14987: dataIn1 = 32'd604
; 
32'd14988: dataIn1 = 32'd607
; 
32'd14989: dataIn1 = 32'd609
; 
32'd14990: dataIn1 = 32'd620
; 
32'd14991: dataIn1 = 32'd623
; 
32'd14992: dataIn1 = 32'd625
; 
32'd14993: dataIn1 = 32'd648
; 
32'd14994: dataIn1 = 32'd663
; 
32'd14995: dataIn1 = 32'd670
; 
32'd14996: dataIn1 = 32'd678
; 
32'd14997: dataIn1 = 32'd694
; 
32'd14998: dataIn1 = 32'd703
; 
32'd14999: dataIn1 = 32'd715
; 
32'd15000: dataIn1 = 32'd730
; 
32'd15001: dataIn1 = 32'd781
; 
32'd15002: dataIn1 = 32'd171
; 
32'd15003: dataIn1 = 32'd179
; 
32'd15004: dataIn1 = 32'd181
; 
32'd15005: dataIn1 = 32'd219
; 
32'd15006: dataIn1 = 32'd303
; 
32'd15007: dataIn1 = 32'd315
; 
32'd15008: dataIn1 = 32'd319
; 
32'd15009: dataIn1 = 32'd322
; 
32'd15010: dataIn1 = 32'd339
; 
32'd15011: dataIn1 = 32'd402
; 
32'd15012: dataIn1 = 32'd436
; 
32'd15013: dataIn1 = 32'd452
; 
32'd15014: dataIn1 = 32'd462
; 
32'd15015: dataIn1 = 32'd471
; 
32'd15016: dataIn1 = 32'd519
; 
32'd15017: dataIn1 = 32'd547
; 
32'd15018: dataIn1 = 32'd569
; 
32'd15019: dataIn1 = 32'd589
; 
32'd15020: dataIn1 = 32'd667
; 
32'd15021: dataIn1 = 32'd670
; 
32'd15022: dataIn1 = 32'd675
; 
32'd15023: dataIn1 = 32'd679
; 
32'd15024: dataIn1 = 32'd681
; 
32'd15025: dataIn1 = 32'd704
; 
32'd15026: dataIn1 = 32'd741
; 
32'd15027: dataIn1 = 32'd749
; 
32'd15028: dataIn1 = 32'd752
; 
32'd15029: dataIn1 = 32'd765
; 
32'd15030: dataIn1 = 32'd773
; 
32'd15031: dataIn1 = 32'd777
; 
32'd15032: dataIn1 = 32'd784
; 
32'd15033: dataIn1 = 32'd787
; 
32'd15034: dataIn1 = 32'd172
; 
32'd15035: dataIn1 = 32'd177
; 
32'd15036: dataIn1 = 32'd180
; 
32'd15037: dataIn1 = 32'd187
; 
32'd15038: dataIn1 = 32'd226
; 
32'd15039: dataIn1 = 32'd229
; 
32'd15040: dataIn1 = 32'd248
; 
32'd15041: dataIn1 = 32'd252
; 
32'd15042: dataIn1 = 32'd256
; 
32'd15043: dataIn1 = 32'd280
; 
32'd15044: dataIn1 = 32'd291
; 
32'd15045: dataIn1 = 32'd306
; 
32'd15046: dataIn1 = 32'd310
; 
32'd15047: dataIn1 = 32'd371
; 
32'd15048: dataIn1 = 32'd378
; 
32'd15049: dataIn1 = 32'd398
; 
32'd15050: dataIn1 = 32'd430
; 
32'd15051: dataIn1 = 32'd447
; 
32'd15052: dataIn1 = 32'd448
; 
32'd15053: dataIn1 = 32'd467
; 
32'd15054: dataIn1 = 32'd477
; 
32'd15055: dataIn1 = 32'd485
; 
32'd15056: dataIn1 = 32'd516
; 
32'd15057: dataIn1 = 32'd518
; 
32'd15058: dataIn1 = 32'd526
; 
32'd15059: dataIn1 = 32'd545
; 
32'd15060: dataIn1 = 32'd577
; 
32'd15061: dataIn1 = 32'd589
; 
32'd15062: dataIn1 = 32'd591
; 
32'd15063: dataIn1 = 32'd604
; 
32'd15064: dataIn1 = 32'd606
; 
32'd15065: dataIn1 = 32'd610
; 
32'd15066: dataIn1 = 32'd612
; 
32'd15067: dataIn1 = 32'd620
; 
32'd15068: dataIn1 = 32'd632
; 
32'd15069: dataIn1 = 32'd656
; 
32'd15070: dataIn1 = 32'd679
; 
32'd15071: dataIn1 = 32'd684
; 
32'd15072: dataIn1 = 32'd718
; 
32'd15073: dataIn1 = 32'd737
; 
32'd15074: dataIn1 = 32'd790
; 
32'd15075: dataIn1 = 32'd177
; 
32'd15076: dataIn1 = 32'd187
; 
32'd15077: dataIn1 = 32'd199
; 
32'd15078: dataIn1 = 32'd210
; 
32'd15079: dataIn1 = 32'd211
; 
32'd15080: dataIn1 = 32'd225
; 
32'd15081: dataIn1 = 32'd247
; 
32'd15082: dataIn1 = 32'd258
; 
32'd15083: dataIn1 = 32'd268
; 
32'd15084: dataIn1 = 32'd295
; 
32'd15085: dataIn1 = 32'd316
; 
32'd15086: dataIn1 = 32'd324
; 
32'd15087: dataIn1 = 32'd351
; 
32'd15088: dataIn1 = 32'd368
; 
32'd15089: dataIn1 = 32'd381
; 
32'd15090: dataIn1 = 32'd409
; 
32'd15091: dataIn1 = 32'd414
; 
32'd15092: dataIn1 = 32'd477
; 
32'd15093: dataIn1 = 32'd485
; 
32'd15094: dataIn1 = 32'd497
; 
32'd15095: dataIn1 = 32'd510
; 
32'd15096: dataIn1 = 32'd515
; 
32'd15097: dataIn1 = 32'd518
; 
32'd15098: dataIn1 = 32'd527
; 
32'd15099: dataIn1 = 32'd539
; 
32'd15100: dataIn1 = 32'd546
; 
32'd15101: dataIn1 = 32'd553
; 
32'd15102: dataIn1 = 32'd582
; 
32'd15103: dataIn1 = 32'd585
; 
32'd15104: dataIn1 = 32'd587
; 
32'd15105: dataIn1 = 32'd605
; 
32'd15106: dataIn1 = 32'd607
; 
32'd15107: dataIn1 = 32'd627
; 
32'd15108: dataIn1 = 32'd630
; 
32'd15109: dataIn1 = 32'd642
; 
32'd15110: dataIn1 = 32'd646
; 
32'd15111: dataIn1 = 32'd648
; 
32'd15112: dataIn1 = 32'd650
; 
32'd15113: dataIn1 = 32'd656
; 
32'd15114: dataIn1 = 32'd687
; 
32'd15115: dataIn1 = 32'd690
; 
32'd15116: dataIn1 = 32'd694
; 
32'd15117: dataIn1 = 32'd699
; 
32'd15118: dataIn1 = 32'd706
; 
32'd15119: dataIn1 = 32'd714
; 
32'd15120: dataIn1 = 32'd734
; 
32'd15121: dataIn1 = 32'd187
; 
32'd15122: dataIn1 = 32'd218
; 
32'd15123: dataIn1 = 32'd221
; 
32'd15124: dataIn1 = 32'd223
; 
32'd15125: dataIn1 = 32'd240
; 
32'd15126: dataIn1 = 32'd281
; 
32'd15127: dataIn1 = 32'd285
; 
32'd15128: dataIn1 = 32'd286
; 
32'd15129: dataIn1 = 32'd318
; 
32'd15130: dataIn1 = 32'd320
; 
32'd15131: dataIn1 = 32'd349
; 
32'd15132: dataIn1 = 32'd364
; 
32'd15133: dataIn1 = 32'd377
; 
32'd15134: dataIn1 = 32'd397
; 
32'd15135: dataIn1 = 32'd399
; 
32'd15136: dataIn1 = 32'd408
; 
32'd15137: dataIn1 = 32'd411
; 
32'd15138: dataIn1 = 32'd428
; 
32'd15139: dataIn1 = 32'd470
; 
32'd15140: dataIn1 = 32'd476
; 
32'd15141: dataIn1 = 32'd511
; 
32'd15142: dataIn1 = 32'd523
; 
32'd15143: dataIn1 = 32'd524
; 
32'd15144: dataIn1 = 32'd546
; 
32'd15145: dataIn1 = 32'd599
; 
32'd15146: dataIn1 = 32'd613
; 
32'd15147: dataIn1 = 32'd615
; 
32'd15148: dataIn1 = 32'd623
; 
32'd15149: dataIn1 = 32'd625
; 
32'd15150: dataIn1 = 32'd631
; 
32'd15151: dataIn1 = 32'd635
; 
32'd15152: dataIn1 = 32'd641
; 
32'd15153: dataIn1 = 32'd661
; 
32'd15154: dataIn1 = 32'd694
; 
32'd15155: dataIn1 = 32'd756
; 
32'd15156: dataIn1 = 32'd800
; 
32'd15157: dataIn1 = 32'd208
; 
32'd15158: dataIn1 = 32'd218
; 
32'd15159: dataIn1 = 32'd220
; 
32'd15160: dataIn1 = 32'd230
; 
32'd15161: dataIn1 = 32'd249
; 
32'd15162: dataIn1 = 32'd267
; 
32'd15163: dataIn1 = 32'd269
; 
32'd15164: dataIn1 = 32'd278
; 
32'd15165: dataIn1 = 32'd292
; 
32'd15166: dataIn1 = 32'd294
; 
32'd15167: dataIn1 = 32'd299
; 
32'd15168: dataIn1 = 32'd325
; 
32'd15169: dataIn1 = 32'd333
; 
32'd15170: dataIn1 = 32'd372
; 
32'd15171: dataIn1 = 32'd373
; 
32'd15172: dataIn1 = 32'd385
; 
32'd15173: dataIn1 = 32'd418
; 
32'd15174: dataIn1 = 32'd420
; 
32'd15175: dataIn1 = 32'd433
; 
32'd15176: dataIn1 = 32'd443
; 
32'd15177: dataIn1 = 32'd454
; 
32'd15178: dataIn1 = 32'd455
; 
32'd15179: dataIn1 = 32'd468
; 
32'd15180: dataIn1 = 32'd470
; 
32'd15181: dataIn1 = 32'd479
; 
32'd15182: dataIn1 = 32'd481
; 
32'd15183: dataIn1 = 32'd521
; 
32'd15184: dataIn1 = 32'd541
; 
32'd15185: dataIn1 = 32'd587
; 
32'd15186: dataIn1 = 32'd588
; 
32'd15187: dataIn1 = 32'd598
; 
32'd15188: dataIn1 = 32'd609
; 
32'd15189: dataIn1 = 32'd635
; 
32'd15190: dataIn1 = 32'd649
; 
32'd15191: dataIn1 = 32'd654
; 
32'd15192: dataIn1 = 32'd681
; 
32'd15193: dataIn1 = 32'd682
; 
32'd15194: dataIn1 = 32'd691
; 
32'd15195: dataIn1 = 32'd709
; 
32'd15196: dataIn1 = 32'd733
; 
32'd15197: dataIn1 = 32'd736
; 
32'd15198: dataIn1 = 32'd742
; 
32'd15199: dataIn1 = 32'd743
; 
32'd15200: dataIn1 = 32'd748
; 
32'd15201: dataIn1 = 32'd750
; 
32'd15202: dataIn1 = 32'd781
; 
32'd15203: dataIn1 = 32'd171
; 
32'd15204: dataIn1 = 32'd198
; 
32'd15205: dataIn1 = 32'd201
; 
32'd15206: dataIn1 = 32'd239
; 
32'd15207: dataIn1 = 32'd242
; 
32'd15208: dataIn1 = 32'd244
; 
32'd15209: dataIn1 = 32'd296
; 
32'd15210: dataIn1 = 32'd313
; 
32'd15211: dataIn1 = 32'd333
; 
32'd15212: dataIn1 = 32'd342
; 
32'd15213: dataIn1 = 32'd355
; 
32'd15214: dataIn1 = 32'd378
; 
32'd15215: dataIn1 = 32'd381
; 
32'd15216: dataIn1 = 32'd403
; 
32'd15217: dataIn1 = 32'd408
; 
32'd15218: dataIn1 = 32'd433
; 
32'd15219: dataIn1 = 32'd446
; 
32'd15220: dataIn1 = 32'd449
; 
32'd15221: dataIn1 = 32'd457
; 
32'd15222: dataIn1 = 32'd474
; 
32'd15223: dataIn1 = 32'd482
; 
32'd15224: dataIn1 = 32'd516
; 
32'd15225: dataIn1 = 32'd530
; 
32'd15226: dataIn1 = 32'd536
; 
32'd15227: dataIn1 = 32'd543
; 
32'd15228: dataIn1 = 32'd546
; 
32'd15229: dataIn1 = 32'd580
; 
32'd15230: dataIn1 = 32'd591
; 
32'd15231: dataIn1 = 32'd596
; 
32'd15232: dataIn1 = 32'd601
; 
32'd15233: dataIn1 = 32'd650
; 
32'd15234: dataIn1 = 32'd661
; 
32'd15235: dataIn1 = 32'd675
; 
32'd15236: dataIn1 = 32'd690
; 
32'd15237: dataIn1 = 32'd695
; 
32'd15238: dataIn1 = 32'd715
; 
32'd15239: dataIn1 = 32'd742
; 
32'd15240: dataIn1 = 32'd748
; 
32'd15241: dataIn1 = 32'd765
; 
32'd15242: dataIn1 = 32'd769
; 
32'd15243: dataIn1 = 32'd779
; 
32'd15244: dataIn1 = 32'd175
; 
32'd15245: dataIn1 = 32'd177
; 
32'd15246: dataIn1 = 32'd190
; 
32'd15247: dataIn1 = 32'd191
; 
32'd15248: dataIn1 = 32'd202
; 
32'd15249: dataIn1 = 32'd206
; 
32'd15250: dataIn1 = 32'd247
; 
32'd15251: dataIn1 = 32'd258
; 
32'd15252: dataIn1 = 32'd293
; 
32'd15253: dataIn1 = 32'd297
; 
32'd15254: dataIn1 = 32'd320
; 
32'd15255: dataIn1 = 32'd348
; 
32'd15256: dataIn1 = 32'd361
; 
32'd15257: dataIn1 = 32'd389
; 
32'd15258: dataIn1 = 32'd436
; 
32'd15259: dataIn1 = 32'd468
; 
32'd15260: dataIn1 = 32'd471
; 
32'd15261: dataIn1 = 32'd498
; 
32'd15262: dataIn1 = 32'd499
; 
32'd15263: dataIn1 = 32'd504
; 
32'd15264: dataIn1 = 32'd510
; 
32'd15265: dataIn1 = 32'd548
; 
32'd15266: dataIn1 = 32'd557
; 
32'd15267: dataIn1 = 32'd560
; 
32'd15268: dataIn1 = 32'd629
; 
32'd15269: dataIn1 = 32'd631
; 
32'd15270: dataIn1 = 32'd645
; 
32'd15271: dataIn1 = 32'd662
; 
32'd15272: dataIn1 = 32'd670
; 
32'd15273: dataIn1 = 32'd671
; 
32'd15274: dataIn1 = 32'd675
; 
32'd15275: dataIn1 = 32'd686
; 
32'd15276: dataIn1 = 32'd706
; 
32'd15277: dataIn1 = 32'd760
; 
32'd15278: dataIn1 = 32'd767
; 
32'd15279: dataIn1 = 32'd182
; 
32'd15280: dataIn1 = 32'd219
; 
32'd15281: dataIn1 = 32'd236
; 
32'd15282: dataIn1 = 32'd238
; 
32'd15283: dataIn1 = 32'd282
; 
32'd15284: dataIn1 = 32'd296
; 
32'd15285: dataIn1 = 32'd307
; 
32'd15286: dataIn1 = 32'd311
; 
32'd15287: dataIn1 = 32'd354
; 
32'd15288: dataIn1 = 32'd376
; 
32'd15289: dataIn1 = 32'd435
; 
32'd15290: dataIn1 = 32'd463
; 
32'd15291: dataIn1 = 32'd475
; 
32'd15292: dataIn1 = 32'd544
; 
32'd15293: dataIn1 = 32'd546
; 
32'd15294: dataIn1 = 32'd551
; 
32'd15295: dataIn1 = 32'd588
; 
32'd15296: dataIn1 = 32'd610
; 
32'd15297: dataIn1 = 32'd620
; 
32'd15298: dataIn1 = 32'd635
; 
32'd15299: dataIn1 = 32'd636
; 
32'd15300: dataIn1 = 32'd640
; 
32'd15301: dataIn1 = 32'd642
; 
32'd15302: dataIn1 = 32'd646
; 
32'd15303: dataIn1 = 32'd670
; 
32'd15304: dataIn1 = 32'd707
; 
32'd15305: dataIn1 = 32'd723
; 
32'd15306: dataIn1 = 32'd746
; 
32'd15307: dataIn1 = 32'd769
; 
32'd15308: dataIn1 = 32'd776
; 
32'd15309: dataIn1 = 32'd794
; 
32'd15310: dataIn1 = 32'd182
; 
32'd15311: dataIn1 = 32'd216
; 
32'd15312: dataIn1 = 32'd226
; 
32'd15313: dataIn1 = 32'd233
; 
32'd15314: dataIn1 = 32'd234
; 
32'd15315: dataIn1 = 32'd237
; 
32'd15316: dataIn1 = 32'd251
; 
32'd15317: dataIn1 = 32'd273
; 
32'd15318: dataIn1 = 32'd354
; 
32'd15319: dataIn1 = 32'd377
; 
32'd15320: dataIn1 = 32'd415
; 
32'd15321: dataIn1 = 32'd455
; 
32'd15322: dataIn1 = 32'd461
; 
32'd15323: dataIn1 = 32'd473
; 
32'd15324: dataIn1 = 32'd499
; 
32'd15325: dataIn1 = 32'd516
; 
32'd15326: dataIn1 = 32'd523
; 
32'd15327: dataIn1 = 32'd569
; 
32'd15328: dataIn1 = 32'd619
; 
32'd15329: dataIn1 = 32'd648
; 
32'd15330: dataIn1 = 32'd655
; 
32'd15331: dataIn1 = 32'd657
; 
32'd15332: dataIn1 = 32'd659
; 
32'd15333: dataIn1 = 32'd663
; 
32'd15334: dataIn1 = 32'd669
; 
32'd15335: dataIn1 = 32'd689
; 
32'd15336: dataIn1 = 32'd690
; 
32'd15337: dataIn1 = 32'd695
; 
32'd15338: dataIn1 = 32'd715
; 
32'd15339: dataIn1 = 32'd733
; 
32'd15340: dataIn1 = 32'd739
; 
32'd15341: dataIn1 = 32'd757
; 
32'd15342: dataIn1 = 32'd788
; 
32'd15343: dataIn1 = 32'd791
; 
32'd15344: dataIn1 = 32'd211
; 
32'd15345: dataIn1 = 32'd218
; 
32'd15346: dataIn1 = 32'd225
; 
32'd15347: dataIn1 = 32'd233
; 
32'd15348: dataIn1 = 32'd249
; 
32'd15349: dataIn1 = 32'd279
; 
32'd15350: dataIn1 = 32'd299
; 
32'd15351: dataIn1 = 32'd314
; 
32'd15352: dataIn1 = 32'd316
; 
32'd15353: dataIn1 = 32'd322
; 
32'd15354: dataIn1 = 32'd323
; 
32'd15355: dataIn1 = 32'd341
; 
32'd15356: dataIn1 = 32'd351
; 
32'd15357: dataIn1 = 32'd372
; 
32'd15358: dataIn1 = 32'd386
; 
32'd15359: dataIn1 = 32'd388
; 
32'd15360: dataIn1 = 32'd418
; 
32'd15361: dataIn1 = 32'd421
; 
32'd15362: dataIn1 = 32'd422
; 
32'd15363: dataIn1 = 32'd431
; 
32'd15364: dataIn1 = 32'd462
; 
32'd15365: dataIn1 = 32'd463
; 
32'd15366: dataIn1 = 32'd466
; 
32'd15367: dataIn1 = 32'd470
; 
32'd15368: dataIn1 = 32'd472
; 
32'd15369: dataIn1 = 32'd475
; 
32'd15370: dataIn1 = 32'd487
; 
32'd15371: dataIn1 = 32'd525
; 
32'd15372: dataIn1 = 32'd536
; 
32'd15373: dataIn1 = 32'd549
; 
32'd15374: dataIn1 = 32'd586
; 
32'd15375: dataIn1 = 32'd603
; 
32'd15376: dataIn1 = 32'd609
; 
32'd15377: dataIn1 = 32'd616
; 
32'd15378: dataIn1 = 32'd618
; 
32'd15379: dataIn1 = 32'd626
; 
32'd15380: dataIn1 = 32'd642
; 
32'd15381: dataIn1 = 32'd659
; 
32'd15382: dataIn1 = 32'd672
; 
32'd15383: dataIn1 = 32'd691
; 
32'd15384: dataIn1 = 32'd710
; 
32'd15385: dataIn1 = 32'd711
; 
32'd15386: dataIn1 = 32'd719
; 
32'd15387: dataIn1 = 32'd735
; 
32'd15388: dataIn1 = 32'd738
; 
32'd15389: dataIn1 = 32'd746
; 
32'd15390: dataIn1 = 32'd764
; 
32'd15391: dataIn1 = 32'd780
; 
32'd15392: dataIn1 = 32'd782
; 
32'd15393: dataIn1 = 32'd191
; 
32'd15394: dataIn1 = 32'd193
; 
32'd15395: dataIn1 = 32'd201
; 
32'd15396: dataIn1 = 32'd205
; 
32'd15397: dataIn1 = 32'd208
; 
32'd15398: dataIn1 = 32'd225
; 
32'd15399: dataIn1 = 32'd243
; 
32'd15400: dataIn1 = 32'd248
; 
32'd15401: dataIn1 = 32'd249
; 
32'd15402: dataIn1 = 32'd259
; 
32'd15403: dataIn1 = 32'd276
; 
32'd15404: dataIn1 = 32'd280
; 
32'd15405: dataIn1 = 32'd316
; 
32'd15406: dataIn1 = 32'd329
; 
32'd15407: dataIn1 = 32'd358
; 
32'd15408: dataIn1 = 32'd359
; 
32'd15409: dataIn1 = 32'd371
; 
32'd15410: dataIn1 = 32'd381
; 
32'd15411: dataIn1 = 32'd398
; 
32'd15412: dataIn1 = 32'd423
; 
32'd15413: dataIn1 = 32'd444
; 
32'd15414: dataIn1 = 32'd472
; 
32'd15415: dataIn1 = 32'd483
; 
32'd15416: dataIn1 = 32'd489
; 
32'd15417: dataIn1 = 32'd535
; 
32'd15418: dataIn1 = 32'd552
; 
32'd15419: dataIn1 = 32'd559
; 
32'd15420: dataIn1 = 32'd578
; 
32'd15421: dataIn1 = 32'd638
; 
32'd15422: dataIn1 = 32'd658
; 
32'd15423: dataIn1 = 32'd659
; 
32'd15424: dataIn1 = 32'd664
; 
32'd15425: dataIn1 = 32'd691
; 
32'd15426: dataIn1 = 32'd697
; 
32'd15427: dataIn1 = 32'd703
; 
32'd15428: dataIn1 = 32'd735
; 
32'd15429: dataIn1 = 32'd771
; 
32'd15430: dataIn1 = 32'd781
; 
32'd15431: dataIn1 = 32'd786
; 
32'd15432: dataIn1 = 32'd181
; 
32'd15433: dataIn1 = 32'd188
; 
32'd15434: dataIn1 = 32'd223
; 
32'd15435: dataIn1 = 32'd224
; 
32'd15436: dataIn1 = 32'd272
; 
32'd15437: dataIn1 = 32'd292
; 
32'd15438: dataIn1 = 32'd326
; 
32'd15439: dataIn1 = 32'd333
; 
32'd15440: dataIn1 = 32'd343
; 
32'd15441: dataIn1 = 32'd344
; 
32'd15442: dataIn1 = 32'd349
; 
32'd15443: dataIn1 = 32'd375
; 
32'd15444: dataIn1 = 32'd386
; 
32'd15445: dataIn1 = 32'd395
; 
32'd15446: dataIn1 = 32'd486
; 
32'd15447: dataIn1 = 32'd496
; 
32'd15448: dataIn1 = 32'd504
; 
32'd15449: dataIn1 = 32'd510
; 
32'd15450: dataIn1 = 32'd518
; 
32'd15451: dataIn1 = 32'd536
; 
32'd15452: dataIn1 = 32'd548
; 
32'd15453: dataIn1 = 32'd563
; 
32'd15454: dataIn1 = 32'd569
; 
32'd15455: dataIn1 = 32'd573
; 
32'd15456: dataIn1 = 32'd585
; 
32'd15457: dataIn1 = 32'd589
; 
32'd15458: dataIn1 = 32'd595
; 
32'd15459: dataIn1 = 32'd602
; 
32'd15460: dataIn1 = 32'd619
; 
32'd15461: dataIn1 = 32'd629
; 
32'd15462: dataIn1 = 32'd656
; 
32'd15463: dataIn1 = 32'd659
; 
32'd15464: dataIn1 = 32'd667
; 
32'd15465: dataIn1 = 32'd671
; 
32'd15466: dataIn1 = 32'd677
; 
32'd15467: dataIn1 = 32'd679
; 
32'd15468: dataIn1 = 32'd681
; 
32'd15469: dataIn1 = 32'd683
; 
32'd15470: dataIn1 = 32'd687
; 
32'd15471: dataIn1 = 32'd703
; 
32'd15472: dataIn1 = 32'd732
; 
32'd15473: dataIn1 = 32'd769
; 
32'd15474: dataIn1 = 32'd774
; 
32'd15475: dataIn1 = 32'd787
; 
32'd15476: dataIn1 = 32'd195
; 
32'd15477: dataIn1 = 32'd203
; 
32'd15478: dataIn1 = 32'd205
; 
32'd15479: dataIn1 = 32'd242
; 
32'd15480: dataIn1 = 32'd276
; 
32'd15481: dataIn1 = 32'd302
; 
32'd15482: dataIn1 = 32'd312
; 
32'd15483: dataIn1 = 32'd316
; 
32'd15484: dataIn1 = 32'd365
; 
32'd15485: dataIn1 = 32'd374
; 
32'd15486: dataIn1 = 32'd397
; 
32'd15487: dataIn1 = 32'd398
; 
32'd15488: dataIn1 = 32'd407
; 
32'd15489: dataIn1 = 32'd408
; 
32'd15490: dataIn1 = 32'd433
; 
32'd15491: dataIn1 = 32'd485
; 
32'd15492: dataIn1 = 32'd504
; 
32'd15493: dataIn1 = 32'd516
; 
32'd15494: dataIn1 = 32'd547
; 
32'd15495: dataIn1 = 32'd553
; 
32'd15496: dataIn1 = 32'd578
; 
32'd15497: dataIn1 = 32'd583
; 
32'd15498: dataIn1 = 32'd600
; 
32'd15499: dataIn1 = 32'd606
; 
32'd15500: dataIn1 = 32'd656
; 
32'd15501: dataIn1 = 32'd665
; 
32'd15502: dataIn1 = 32'd733
; 
32'd15503: dataIn1 = 32'd746
; 
32'd15504: dataIn1 = 32'd756
; 
32'd15505: dataIn1 = 32'd768
; 
32'd15506: dataIn1 = 32'd180
; 
32'd15507: dataIn1 = 32'd190
; 
32'd15508: dataIn1 = 32'd202
; 
32'd15509: dataIn1 = 32'd222
; 
32'd15510: dataIn1 = 32'd229
; 
32'd15511: dataIn1 = 32'd242
; 
32'd15512: dataIn1 = 32'd257
; 
32'd15513: dataIn1 = 32'd276
; 
32'd15514: dataIn1 = 32'd290
; 
32'd15515: dataIn1 = 32'd291
; 
32'd15516: dataIn1 = 32'd314
; 
32'd15517: dataIn1 = 32'd331
; 
32'd15518: dataIn1 = 32'd379
; 
32'd15519: dataIn1 = 32'd406
; 
32'd15520: dataIn1 = 32'd408
; 
32'd15521: dataIn1 = 32'd429
; 
32'd15522: dataIn1 = 32'd452
; 
32'd15523: dataIn1 = 32'd499
; 
32'd15524: dataIn1 = 32'd508
; 
32'd15525: dataIn1 = 32'd511
; 
32'd15526: dataIn1 = 32'd547
; 
32'd15527: dataIn1 = 32'd595
; 
32'd15528: dataIn1 = 32'd605
; 
32'd15529: dataIn1 = 32'd609
; 
32'd15530: dataIn1 = 32'd627
; 
32'd15531: dataIn1 = 32'd643
; 
32'd15532: dataIn1 = 32'd651
; 
32'd15533: dataIn1 = 32'd655
; 
32'd15534: dataIn1 = 32'd676
; 
32'd15535: dataIn1 = 32'd689
; 
32'd15536: dataIn1 = 32'd719
; 
32'd15537: dataIn1 = 32'd722
; 
32'd15538: dataIn1 = 32'd724
; 
32'd15539: dataIn1 = 32'd749
; 
32'd15540: dataIn1 = 32'd760
; 
32'd15541: dataIn1 = 32'd761
; 
32'd15542: dataIn1 = 32'd769
; 
32'd15543: dataIn1 = 32'd771
; 
32'd15544: dataIn1 = 32'd786
; 
32'd15545: dataIn1 = 32'd799
; 
32'd15546: dataIn1 = 32'd186
; 
32'd15547: dataIn1 = 32'd201
; 
32'd15548: dataIn1 = 32'd209
; 
32'd15549: dataIn1 = 32'd237
; 
32'd15550: dataIn1 = 32'd243
; 
32'd15551: dataIn1 = 32'd264
; 
32'd15552: dataIn1 = 32'd266
; 
32'd15553: dataIn1 = 32'd295
; 
32'd15554: dataIn1 = 32'd318
; 
32'd15555: dataIn1 = 32'd351
; 
32'd15556: dataIn1 = 32'd399
; 
32'd15557: dataIn1 = 32'd404
; 
32'd15558: dataIn1 = 32'd426
; 
32'd15559: dataIn1 = 32'd431
; 
32'd15560: dataIn1 = 32'd432
; 
32'd15561: dataIn1 = 32'd457
; 
32'd15562: dataIn1 = 32'd465
; 
32'd15563: dataIn1 = 32'd471
; 
32'd15564: dataIn1 = 32'd479
; 
32'd15565: dataIn1 = 32'd488
; 
32'd15566: dataIn1 = 32'd517
; 
32'd15567: dataIn1 = 32'd533
; 
32'd15568: dataIn1 = 32'd546
; 
32'd15569: dataIn1 = 32'd562
; 
32'd15570: dataIn1 = 32'd575
; 
32'd15571: dataIn1 = 32'd601
; 
32'd15572: dataIn1 = 32'd619
; 
32'd15573: dataIn1 = 32'd620
; 
32'd15574: dataIn1 = 32'd663
; 
32'd15575: dataIn1 = 32'd740
; 
32'd15576: dataIn1 = 32'd751
; 
32'd15577: dataIn1 = 32'd774
; 
32'd15578: dataIn1 = 32'd190
; 
32'd15579: dataIn1 = 32'd216
; 
32'd15580: dataIn1 = 32'd240
; 
32'd15581: dataIn1 = 32'd247
; 
32'd15582: dataIn1 = 32'd254
; 
32'd15583: dataIn1 = 32'd259
; 
32'd15584: dataIn1 = 32'd308
; 
32'd15585: dataIn1 = 32'd322
; 
32'd15586: dataIn1 = 32'd382
; 
32'd15587: dataIn1 = 32'd492
; 
32'd15588: dataIn1 = 32'd539
; 
32'd15589: dataIn1 = 32'd541
; 
32'd15590: dataIn1 = 32'd548
; 
32'd15591: dataIn1 = 32'd563
; 
32'd15592: dataIn1 = 32'd597
; 
32'd15593: dataIn1 = 32'd644
; 
32'd15594: dataIn1 = 32'd688
; 
32'd15595: dataIn1 = 32'd698
; 
32'd15596: dataIn1 = 32'd736
; 
32'd15597: dataIn1 = 32'd754
; 
32'd15598: dataIn1 = 32'd760
; 
32'd15599: dataIn1 = 32'd773
; 
32'd15600: dataIn1 = 32'd776
; 
32'd15601: dataIn1 = 32'd794
; 
32'd15602: dataIn1 = 32'd799
; 
32'd15603: dataIn1 = 32'd217
; 
32'd15604: dataIn1 = 32'd243
; 
32'd15605: dataIn1 = 32'd263
; 
32'd15606: dataIn1 = 32'd281
; 
32'd15607: dataIn1 = 32'd294
; 
32'd15608: dataIn1 = 32'd297
; 
32'd15609: dataIn1 = 32'd304
; 
32'd15610: dataIn1 = 32'd359
; 
32'd15611: dataIn1 = 32'd378
; 
32'd15612: dataIn1 = 32'd380
; 
32'd15613: dataIn1 = 32'd398
; 
32'd15614: dataIn1 = 32'd410
; 
32'd15615: dataIn1 = 32'd412
; 
32'd15616: dataIn1 = 32'd420
; 
32'd15617: dataIn1 = 32'd428
; 
32'd15618: dataIn1 = 32'd429
; 
32'd15619: dataIn1 = 32'd432
; 
32'd15620: dataIn1 = 32'd454
; 
32'd15621: dataIn1 = 32'd466
; 
32'd15622: dataIn1 = 32'd481
; 
32'd15623: dataIn1 = 32'd504
; 
32'd15624: dataIn1 = 32'd565
; 
32'd15625: dataIn1 = 32'd574
; 
32'd15626: dataIn1 = 32'd581
; 
32'd15627: dataIn1 = 32'd606
; 
32'd15628: dataIn1 = 32'd617
; 
32'd15629: dataIn1 = 32'd666
; 
32'd15630: dataIn1 = 32'd678
; 
32'd15631: dataIn1 = 32'd702
; 
32'd15632: dataIn1 = 32'd730
; 
32'd15633: dataIn1 = 32'd758
; 
32'd15634: dataIn1 = 32'd763
; 
32'd15635: dataIn1 = 32'd768
; 
32'd15636: dataIn1 = 32'd798
; 
32'd15637: dataIn1 = 32'd204
; 
32'd15638: dataIn1 = 32'd223
; 
32'd15639: dataIn1 = 32'd232
; 
32'd15640: dataIn1 = 32'd249
; 
32'd15641: dataIn1 = 32'd265
; 
32'd15642: dataIn1 = 32'd300
; 
32'd15643: dataIn1 = 32'd310
; 
32'd15644: dataIn1 = 32'd355
; 
32'd15645: dataIn1 = 32'd373
; 
32'd15646: dataIn1 = 32'd376
; 
32'd15647: dataIn1 = 32'd379
; 
32'd15648: dataIn1 = 32'd399
; 
32'd15649: dataIn1 = 32'd402
; 
32'd15650: dataIn1 = 32'd404
; 
32'd15651: dataIn1 = 32'd408
; 
32'd15652: dataIn1 = 32'd411
; 
32'd15653: dataIn1 = 32'd459
; 
32'd15654: dataIn1 = 32'd462
; 
32'd15655: dataIn1 = 32'd464
; 
32'd15656: dataIn1 = 32'd471
; 
32'd15657: dataIn1 = 32'd472
; 
32'd15658: dataIn1 = 32'd491
; 
32'd15659: dataIn1 = 32'd502
; 
32'd15660: dataIn1 = 32'd525
; 
32'd15661: dataIn1 = 32'd545
; 
32'd15662: dataIn1 = 32'd552
; 
32'd15663: dataIn1 = 32'd557
; 
32'd15664: dataIn1 = 32'd591
; 
32'd15665: dataIn1 = 32'd596
; 
32'd15666: dataIn1 = 32'd603
; 
32'd15667: dataIn1 = 32'd614
; 
32'd15668: dataIn1 = 32'd618
; 
32'd15669: dataIn1 = 32'd645
; 
32'd15670: dataIn1 = 32'd661
; 
32'd15671: dataIn1 = 32'd665
; 
32'd15672: dataIn1 = 32'd672
; 
32'd15673: dataIn1 = 32'd682
; 
32'd15674: dataIn1 = 32'd693
; 
32'd15675: dataIn1 = 32'd719
; 
32'd15676: dataIn1 = 32'd724
; 
32'd15677: dataIn1 = 32'd736
; 
32'd15678: dataIn1 = 32'd771
; 
32'd15679: dataIn1 = 32'd782
; 
32'd15680: dataIn1 = 32'd800
; 
32'd15681: dataIn1 = 32'd185
; 
32'd15682: dataIn1 = 32'd205
; 
32'd15683: dataIn1 = 32'd224
; 
32'd15684: dataIn1 = 32'd231
; 
32'd15685: dataIn1 = 32'd292
; 
32'd15686: dataIn1 = 32'd305
; 
32'd15687: dataIn1 = 32'd315
; 
32'd15688: dataIn1 = 32'd317
; 
32'd15689: dataIn1 = 32'd318
; 
32'd15690: dataIn1 = 32'd340
; 
32'd15691: dataIn1 = 32'd347
; 
32'd15692: dataIn1 = 32'd350
; 
32'd15693: dataIn1 = 32'd351
; 
32'd15694: dataIn1 = 32'd363
; 
32'd15695: dataIn1 = 32'd419
; 
32'd15696: dataIn1 = 32'd421
; 
32'd15697: dataIn1 = 32'd443
; 
32'd15698: dataIn1 = 32'd451
; 
32'd15699: dataIn1 = 32'd462
; 
32'd15700: dataIn1 = 32'd504
; 
32'd15701: dataIn1 = 32'd515
; 
32'd15702: dataIn1 = 32'd530
; 
32'd15703: dataIn1 = 32'd531
; 
32'd15704: dataIn1 = 32'd569
; 
32'd15705: dataIn1 = 32'd593
; 
32'd15706: dataIn1 = 32'd603
; 
32'd15707: dataIn1 = 32'd667
; 
32'd15708: dataIn1 = 32'd698
; 
32'd15709: dataIn1 = 32'd725
; 
32'd15710: dataIn1 = 32'd730
; 
32'd15711: dataIn1 = 32'd741
; 
32'd15712: dataIn1 = 32'd748
; 
32'd15713: dataIn1 = 32'd777
; 
32'd15714: dataIn1 = 32'd779
; 
32'd15715: dataIn1 = 32'd781
; 
32'd15716: dataIn1 = 32'd783
; 
32'd15717: dataIn1 = 32'd785
; 
32'd15718: dataIn1 = 32'd794
; 
32'd15719: dataIn1 = 32'd796
; 
32'd15720: dataIn1 = 32'd209
; 
32'd15721: dataIn1 = 32'd265
; 
32'd15722: dataIn1 = 32'd272
; 
32'd15723: dataIn1 = 32'd278
; 
32'd15724: dataIn1 = 32'd295
; 
32'd15725: dataIn1 = 32'd319
; 
32'd15726: dataIn1 = 32'd330
; 
32'd15727: dataIn1 = 32'd334
; 
32'd15728: dataIn1 = 32'd337
; 
32'd15729: dataIn1 = 32'd339
; 
32'd15730: dataIn1 = 32'd351
; 
32'd15731: dataIn1 = 32'd362
; 
32'd15732: dataIn1 = 32'd378
; 
32'd15733: dataIn1 = 32'd406
; 
32'd15734: dataIn1 = 32'd424
; 
32'd15735: dataIn1 = 32'd449
; 
32'd15736: dataIn1 = 32'd457
; 
32'd15737: dataIn1 = 32'd500
; 
32'd15738: dataIn1 = 32'd532
; 
32'd15739: dataIn1 = 32'd535
; 
32'd15740: dataIn1 = 32'd558
; 
32'd15741: dataIn1 = 32'd569
; 
32'd15742: dataIn1 = 32'd572
; 
32'd15743: dataIn1 = 32'd580
; 
32'd15744: dataIn1 = 32'd607
; 
32'd15745: dataIn1 = 32'd630
; 
32'd15746: dataIn1 = 32'd643
; 
32'd15747: dataIn1 = 32'd658
; 
32'd15748: dataIn1 = 32'd667
; 
32'd15749: dataIn1 = 32'd681
; 
32'd15750: dataIn1 = 32'd733
; 
32'd15751: dataIn1 = 32'd742
; 
32'd15752: dataIn1 = 32'd768
; 
32'd15753: dataIn1 = 32'd774
; 
32'd15754: dataIn1 = 32'd787
; 
32'd15755: dataIn1 = 32'd192
; 
32'd15756: dataIn1 = 32'd220
; 
32'd15757: dataIn1 = 32'd222
; 
32'd15758: dataIn1 = 32'd237
; 
32'd15759: dataIn1 = 32'd239
; 
32'd15760: dataIn1 = 32'd279
; 
32'd15761: dataIn1 = 32'd303
; 
32'd15762: dataIn1 = 32'd319
; 
32'd15763: dataIn1 = 32'd333
; 
32'd15764: dataIn1 = 32'd337
; 
32'd15765: dataIn1 = 32'd384
; 
32'd15766: dataIn1 = 32'd427
; 
32'd15767: dataIn1 = 32'd441
; 
32'd15768: dataIn1 = 32'd443
; 
32'd15769: dataIn1 = 32'd449
; 
32'd15770: dataIn1 = 32'd461
; 
32'd15771: dataIn1 = 32'd463
; 
32'd15772: dataIn1 = 32'd467
; 
32'd15773: dataIn1 = 32'd475
; 
32'd15774: dataIn1 = 32'd480
; 
32'd15775: dataIn1 = 32'd515
; 
32'd15776: dataIn1 = 32'd520
; 
32'd15777: dataIn1 = 32'd534
; 
32'd15778: dataIn1 = 32'd545
; 
32'd15779: dataIn1 = 32'd559
; 
32'd15780: dataIn1 = 32'd570
; 
32'd15781: dataIn1 = 32'd574
; 
32'd15782: dataIn1 = 32'd582
; 
32'd15783: dataIn1 = 32'd593
; 
32'd15784: dataIn1 = 32'd594
; 
32'd15785: dataIn1 = 32'd630
; 
32'd15786: dataIn1 = 32'd706
; 
32'd15787: dataIn1 = 32'd717
; 
32'd15788: dataIn1 = 32'd726
; 
32'd15789: dataIn1 = 32'd775
; 
32'd15790: dataIn1 = 32'd776
; 
32'd15791: dataIn1 = 32'd785
; 
32'd15792: dataIn1 = 32'd786
; 
32'd15793: dataIn1 = 32'd793
; 
32'd15794: dataIn1 = 32'd196
; 
32'd15795: dataIn1 = 32'd205
; 
32'd15796: dataIn1 = 32'd218
; 
32'd15797: dataIn1 = 32'd225
; 
32'd15798: dataIn1 = 32'd265
; 
32'd15799: dataIn1 = 32'd310
; 
32'd15800: dataIn1 = 32'd341
; 
32'd15801: dataIn1 = 32'd344
; 
32'd15802: dataIn1 = 32'd351
; 
32'd15803: dataIn1 = 32'd356
; 
32'd15804: dataIn1 = 32'd364
; 
32'd15805: dataIn1 = 32'd370
; 
32'd15806: dataIn1 = 32'd371
; 
32'd15807: dataIn1 = 32'd387
; 
32'd15808: dataIn1 = 32'd391
; 
32'd15809: dataIn1 = 32'd443
; 
32'd15810: dataIn1 = 32'd458
; 
32'd15811: dataIn1 = 32'd464
; 
32'd15812: dataIn1 = 32'd485
; 
32'd15813: dataIn1 = 32'd486
; 
32'd15814: dataIn1 = 32'd493
; 
32'd15815: dataIn1 = 32'd497
; 
32'd15816: dataIn1 = 32'd510
; 
32'd15817: dataIn1 = 32'd516
; 
32'd15818: dataIn1 = 32'd527
; 
32'd15819: dataIn1 = 32'd532
; 
32'd15820: dataIn1 = 32'd546
; 
32'd15821: dataIn1 = 32'd551
; 
32'd15822: dataIn1 = 32'd584
; 
32'd15823: dataIn1 = 32'd589
; 
32'd15824: dataIn1 = 32'd598
; 
32'd15825: dataIn1 = 32'd614
; 
32'd15826: dataIn1 = 32'd663
; 
32'd15827: dataIn1 = 32'd696
; 
32'd15828: dataIn1 = 32'd709
; 
32'd15829: dataIn1 = 32'd712
; 
32'd15830: dataIn1 = 32'd721
; 
32'd15831: dataIn1 = 32'd724
; 
32'd15832: dataIn1 = 32'd734
; 
32'd15833: dataIn1 = 32'd748
; 
32'd15834: dataIn1 = 32'd749
; 
32'd15835: dataIn1 = 32'd759
; 
32'd15836: dataIn1 = 32'd246
; 
32'd15837: dataIn1 = 32'd296
; 
32'd15838: dataIn1 = 32'd322
; 
32'd15839: dataIn1 = 32'd365
; 
32'd15840: dataIn1 = 32'd371
; 
32'd15841: dataIn1 = 32'd387
; 
32'd15842: dataIn1 = 32'd411
; 
32'd15843: dataIn1 = 32'd414
; 
32'd15844: dataIn1 = 32'd416
; 
32'd15845: dataIn1 = 32'd474
; 
32'd15846: dataIn1 = 32'd484
; 
32'd15847: dataIn1 = 32'd489
; 
32'd15848: dataIn1 = 32'd498
; 
32'd15849: dataIn1 = 32'd523
; 
32'd15850: dataIn1 = 32'd542
; 
32'd15851: dataIn1 = 32'd565
; 
32'd15852: dataIn1 = 32'd576
; 
32'd15853: dataIn1 = 32'd583
; 
32'd15854: dataIn1 = 32'd586
; 
32'd15855: dataIn1 = 32'd588
; 
32'd15856: dataIn1 = 32'd609
; 
32'd15857: dataIn1 = 32'd617
; 
32'd15858: dataIn1 = 32'd622
; 
32'd15859: dataIn1 = 32'd632
; 
32'd15860: dataIn1 = 32'd645
; 
32'd15861: dataIn1 = 32'd652
; 
32'd15862: dataIn1 = 32'd664
; 
32'd15863: dataIn1 = 32'd666
; 
32'd15864: dataIn1 = 32'd728
; 
32'd15865: dataIn1 = 32'd735
; 
32'd15866: dataIn1 = 32'd776
; 
32'd15867: dataIn1 = 32'd200
; 
32'd15868: dataIn1 = 32'd207
; 
32'd15869: dataIn1 = 32'd350
; 
32'd15870: dataIn1 = 32'd354
; 
32'd15871: dataIn1 = 32'd439
; 
32'd15872: dataIn1 = 32'd464
; 
32'd15873: dataIn1 = 32'd469
; 
32'd15874: dataIn1 = 32'd480
; 
32'd15875: dataIn1 = 32'd502
; 
32'd15876: dataIn1 = 32'd514
; 
32'd15877: dataIn1 = 32'd570
; 
32'd15878: dataIn1 = 32'd657
; 
32'd15879: dataIn1 = 32'd683
; 
32'd15880: dataIn1 = 32'd687
; 
32'd15881: dataIn1 = 32'd692
; 
32'd15882: dataIn1 = 32'd700
; 
32'd15883: dataIn1 = 32'd702
; 
32'd15884: dataIn1 = 32'd724
; 
32'd15885: dataIn1 = 32'd738
; 
32'd15886: dataIn1 = 32'd742
; 
32'd15887: dataIn1 = 32'd772
; 
32'd15888: dataIn1 = 32'd796
; 
32'd15889: dataIn1 = 32'd799
; 
32'd15890: dataIn1 = 32'd200
; 
32'd15891: dataIn1 = 32'd225
; 
32'd15892: dataIn1 = 32'd261
; 
32'd15893: dataIn1 = 32'd290
; 
32'd15894: dataIn1 = 32'd304
; 
32'd15895: dataIn1 = 32'd339
; 
32'd15896: dataIn1 = 32'd396
; 
32'd15897: dataIn1 = 32'd403
; 
32'd15898: dataIn1 = 32'd423
; 
32'd15899: dataIn1 = 32'd429
; 
32'd15900: dataIn1 = 32'd441
; 
32'd15901: dataIn1 = 32'd453
; 
32'd15902: dataIn1 = 32'd470
; 
32'd15903: dataIn1 = 32'd488
; 
32'd15904: dataIn1 = 32'd525
; 
32'd15905: dataIn1 = 32'd535
; 
32'd15906: dataIn1 = 32'd569
; 
32'd15907: dataIn1 = 32'd589
; 
32'd15908: dataIn1 = 32'd591
; 
32'd15909: dataIn1 = 32'd598
; 
32'd15910: dataIn1 = 32'd610
; 
32'd15911: dataIn1 = 32'd639
; 
32'd15912: dataIn1 = 32'd654
; 
32'd15913: dataIn1 = 32'd655
; 
32'd15914: dataIn1 = 32'd658
; 
32'd15915: dataIn1 = 32'd665
; 
32'd15916: dataIn1 = 32'd671
; 
32'd15917: dataIn1 = 32'd680
; 
32'd15918: dataIn1 = 32'd681
; 
32'd15919: dataIn1 = 32'd690
; 
32'd15920: dataIn1 = 32'd727
; 
32'd15921: dataIn1 = 32'd796
; 
32'd15922: dataIn1 = 32'd194
; 
32'd15923: dataIn1 = 32'd202
; 
32'd15924: dataIn1 = 32'd203
; 
32'd15925: dataIn1 = 32'd206
; 
32'd15926: dataIn1 = 32'd213
; 
32'd15927: dataIn1 = 32'd224
; 
32'd15928: dataIn1 = 32'd238
; 
32'd15929: dataIn1 = 32'd243
; 
32'd15930: dataIn1 = 32'd260
; 
32'd15931: dataIn1 = 32'd271
; 
32'd15932: dataIn1 = 32'd274
; 
32'd15933: dataIn1 = 32'd331
; 
32'd15934: dataIn1 = 32'd336
; 
32'd15935: dataIn1 = 32'd374
; 
32'd15936: dataIn1 = 32'd391
; 
32'd15937: dataIn1 = 32'd397
; 
32'd15938: dataIn1 = 32'd416
; 
32'd15939: dataIn1 = 32'd446
; 
32'd15940: dataIn1 = 32'd447
; 
32'd15941: dataIn1 = 32'd491
; 
32'd15942: dataIn1 = 32'd496
; 
32'd15943: dataIn1 = 32'd519
; 
32'd15944: dataIn1 = 32'd560
; 
32'd15945: dataIn1 = 32'd569
; 
32'd15946: dataIn1 = 32'd606
; 
32'd15947: dataIn1 = 32'd623
; 
32'd15948: dataIn1 = 32'd638
; 
32'd15949: dataIn1 = 32'd680
; 
32'd15950: dataIn1 = 32'd720
; 
32'd15951: dataIn1 = 32'd736
; 
32'd15952: dataIn1 = 32'd737
; 
32'd15953: dataIn1 = 32'd759
; 
32'd15954: dataIn1 = 32'd760
; 
32'd15955: dataIn1 = 32'd780
; 
32'd15956: dataIn1 = 32'd786
; 
32'd15957: dataIn1 = 32'd791
; 
32'd15958: dataIn1 = 32'd203
; 
32'd15959: dataIn1 = 32'd212
; 
32'd15960: dataIn1 = 32'd215
; 
32'd15961: dataIn1 = 32'd237
; 
32'd15962: dataIn1 = 32'd274
; 
32'd15963: dataIn1 = 32'd308
; 
32'd15964: dataIn1 = 32'd309
; 
32'd15965: dataIn1 = 32'd322
; 
32'd15966: dataIn1 = 32'd330
; 
32'd15967: dataIn1 = 32'd376
; 
32'd15968: dataIn1 = 32'd385
; 
32'd15969: dataIn1 = 32'd392
; 
32'd15970: dataIn1 = 32'd417
; 
32'd15971: dataIn1 = 32'd433
; 
32'd15972: dataIn1 = 32'd464
; 
32'd15973: dataIn1 = 32'd495
; 
32'd15974: dataIn1 = 32'd508
; 
32'd15975: dataIn1 = 32'd547
; 
32'd15976: dataIn1 = 32'd567
; 
32'd15977: dataIn1 = 32'd570
; 
32'd15978: dataIn1 = 32'd577
; 
32'd15979: dataIn1 = 32'd598
; 
32'd15980: dataIn1 = 32'd607
; 
32'd15981: dataIn1 = 32'd622
; 
32'd15982: dataIn1 = 32'd631
; 
32'd15983: dataIn1 = 32'd634
; 
32'd15984: dataIn1 = 32'd648
; 
32'd15985: dataIn1 = 32'd686
; 
32'd15986: dataIn1 = 32'd693
; 
32'd15987: dataIn1 = 32'd703
; 
32'd15988: dataIn1 = 32'd720
; 
32'd15989: dataIn1 = 32'd762
; 
32'd15990: dataIn1 = 32'd773
; 
32'd15991: dataIn1 = 32'd196
; 
32'd15992: dataIn1 = 32'd198
; 
32'd15993: dataIn1 = 32'd205
; 
32'd15994: dataIn1 = 32'd209
; 
32'd15995: dataIn1 = 32'd223
; 
32'd15996: dataIn1 = 32'd246
; 
32'd15997: dataIn1 = 32'd250
; 
32'd15998: dataIn1 = 32'd254
; 
32'd15999: dataIn1 = 32'd291
; 
32'd16000: dataIn1 = 32'd292
; 
32'd16001: dataIn1 = 32'd347
; 
32'd16002: dataIn1 = 32'd354
; 
32'd16003: dataIn1 = 32'd355
; 
32'd16004: dataIn1 = 32'd356
; 
32'd16005: dataIn1 = 32'd365
; 
32'd16006: dataIn1 = 32'd371
; 
32'd16007: dataIn1 = 32'd383
; 
32'd16008: dataIn1 = 32'd392
; 
32'd16009: dataIn1 = 32'd399
; 
32'd16010: dataIn1 = 32'd404
; 
32'd16011: dataIn1 = 32'd413
; 
32'd16012: dataIn1 = 32'd430
; 
32'd16013: dataIn1 = 32'd438
; 
32'd16014: dataIn1 = 32'd459
; 
32'd16015: dataIn1 = 32'd467
; 
32'd16016: dataIn1 = 32'd520
; 
32'd16017: dataIn1 = 32'd524
; 
32'd16018: dataIn1 = 32'd529
; 
32'd16019: dataIn1 = 32'd544
; 
32'd16020: dataIn1 = 32'd554
; 
32'd16021: dataIn1 = 32'd573
; 
32'd16022: dataIn1 = 32'd593
; 
32'd16023: dataIn1 = 32'd608
; 
32'd16024: dataIn1 = 32'd628
; 
32'd16025: dataIn1 = 32'd685
; 
32'd16026: dataIn1 = 32'd716
; 
32'd16027: dataIn1 = 32'd717
; 
32'd16028: dataIn1 = 32'd721
; 
32'd16029: dataIn1 = 32'd732
; 
32'd16030: dataIn1 = 32'd733
; 
32'd16031: dataIn1 = 32'd740
; 
32'd16032: dataIn1 = 32'd765
; 
32'd16033: dataIn1 = 32'd770
; 
32'd16034: dataIn1 = 32'd774
; 
32'd16035: dataIn1 = 32'd799
; 
32'd16036: dataIn1 = 32'd800
; 
32'd16037: dataIn1 = 32'd201
; 
32'd16038: dataIn1 = 32'd225
; 
32'd16039: dataIn1 = 32'd231
; 
32'd16040: dataIn1 = 32'd278
; 
32'd16041: dataIn1 = 32'd321
; 
32'd16042: dataIn1 = 32'd333
; 
32'd16043: dataIn1 = 32'd337
; 
32'd16044: dataIn1 = 32'd339
; 
32'd16045: dataIn1 = 32'd352
; 
32'd16046: dataIn1 = 32'd414
; 
32'd16047: dataIn1 = 32'd426
; 
32'd16048: dataIn1 = 32'd431
; 
32'd16049: dataIn1 = 32'd495
; 
32'd16050: dataIn1 = 32'd496
; 
32'd16051: dataIn1 = 32'd509
; 
32'd16052: dataIn1 = 32'd512
; 
32'd16053: dataIn1 = 32'd523
; 
32'd16054: dataIn1 = 32'd531
; 
32'd16055: dataIn1 = 32'd553
; 
32'd16056: dataIn1 = 32'd560
; 
32'd16057: dataIn1 = 32'd592
; 
32'd16058: dataIn1 = 32'd593
; 
32'd16059: dataIn1 = 32'd604
; 
32'd16060: dataIn1 = 32'd612
; 
32'd16061: dataIn1 = 32'd613
; 
32'd16062: dataIn1 = 32'd644
; 
32'd16063: dataIn1 = 32'd657
; 
32'd16064: dataIn1 = 32'd670
; 
32'd16065: dataIn1 = 32'd708
; 
32'd16066: dataIn1 = 32'd710
; 
32'd16067: dataIn1 = 32'd714
; 
32'd16068: dataIn1 = 32'd715
; 
32'd16069: dataIn1 = 32'd727
; 
32'd16070: dataIn1 = 32'd730
; 
32'd16071: dataIn1 = 32'd755
; 
32'd16072: dataIn1 = 32'd784
; 
32'd16073: dataIn1 = 32'd800
; 
32'd16074: dataIn1 = 32'd199
; 
32'd16075: dataIn1 = 32'd203
; 
32'd16076: dataIn1 = 32'd235
; 
32'd16077: dataIn1 = 32'd265
; 
32'd16078: dataIn1 = 32'd294
; 
32'd16079: dataIn1 = 32'd314
; 
32'd16080: dataIn1 = 32'd338
; 
32'd16081: dataIn1 = 32'd378
; 
32'd16082: dataIn1 = 32'd380
; 
32'd16083: dataIn1 = 32'd394
; 
32'd16084: dataIn1 = 32'd430
; 
32'd16085: dataIn1 = 32'd436
; 
32'd16086: dataIn1 = 32'd444
; 
32'd16087: dataIn1 = 32'd458
; 
32'd16088: dataIn1 = 32'd477
; 
32'd16089: dataIn1 = 32'd506
; 
32'd16090: dataIn1 = 32'd515
; 
32'd16091: dataIn1 = 32'd528
; 
32'd16092: dataIn1 = 32'd534
; 
32'd16093: dataIn1 = 32'd547
; 
32'd16094: dataIn1 = 32'd555
; 
32'd16095: dataIn1 = 32'd558
; 
32'd16096: dataIn1 = 32'd568
; 
32'd16097: dataIn1 = 32'd571
; 
32'd16098: dataIn1 = 32'd601
; 
32'd16099: dataIn1 = 32'd620
; 
32'd16100: dataIn1 = 32'd642
; 
32'd16101: dataIn1 = 32'd647
; 
32'd16102: dataIn1 = 32'd666
; 
32'd16103: dataIn1 = 32'd670
; 
32'd16104: dataIn1 = 32'd691
; 
32'd16105: dataIn1 = 32'd731
; 
32'd16106: dataIn1 = 32'd744
; 
32'd16107: dataIn1 = 32'd755
; 
32'd16108: dataIn1 = 32'd782
; 
32'd16109: dataIn1 = 32'd783
; 
32'd16110: dataIn1 = 32'd791
; 
32'd16111: dataIn1 = 32'd196
; 
32'd16112: dataIn1 = 32'd201
; 
32'd16113: dataIn1 = 32'd204
; 
32'd16114: dataIn1 = 32'd216
; 
32'd16115: dataIn1 = 32'd236
; 
32'd16116: dataIn1 = 32'd284
; 
32'd16117: dataIn1 = 32'd287
; 
32'd16118: dataIn1 = 32'd372
; 
32'd16119: dataIn1 = 32'd383
; 
32'd16120: dataIn1 = 32'd401
; 
32'd16121: dataIn1 = 32'd445
; 
32'd16122: dataIn1 = 32'd446
; 
32'd16123: dataIn1 = 32'd463
; 
32'd16124: dataIn1 = 32'd465
; 
32'd16125: dataIn1 = 32'd466
; 
32'd16126: dataIn1 = 32'd543
; 
32'd16127: dataIn1 = 32'd545
; 
32'd16128: dataIn1 = 32'd550
; 
32'd16129: dataIn1 = 32'd566
; 
32'd16130: dataIn1 = 32'd595
; 
32'd16131: dataIn1 = 32'd613
; 
32'd16132: dataIn1 = 32'd631
; 
32'd16133: dataIn1 = 32'd634
; 
32'd16134: dataIn1 = 32'd639
; 
32'd16135: dataIn1 = 32'd662
; 
32'd16136: dataIn1 = 32'd669
; 
32'd16137: dataIn1 = 32'd672
; 
32'd16138: dataIn1 = 32'd685
; 
32'd16139: dataIn1 = 32'd695
; 
32'd16140: dataIn1 = 32'd704
; 
32'd16141: dataIn1 = 32'd722
; 
32'd16142: dataIn1 = 32'd772
; 
32'd16143: dataIn1 = 32'd773
; 
32'd16144: dataIn1 = 32'd794
; 
32'd16145: dataIn1 = 32'd206
; 
32'd16146: dataIn1 = 32'd213
; 
32'd16147: dataIn1 = 32'd219
; 
32'd16148: dataIn1 = 32'd220
; 
32'd16149: dataIn1 = 32'd221
; 
32'd16150: dataIn1 = 32'd237
; 
32'd16151: dataIn1 = 32'd247
; 
32'd16152: dataIn1 = 32'd262
; 
32'd16153: dataIn1 = 32'd287
; 
32'd16154: dataIn1 = 32'd306
; 
32'd16155: dataIn1 = 32'd313
; 
32'd16156: dataIn1 = 32'd323
; 
32'd16157: dataIn1 = 32'd348
; 
32'd16158: dataIn1 = 32'd356
; 
32'd16159: dataIn1 = 32'd381
; 
32'd16160: dataIn1 = 32'd388
; 
32'd16161: dataIn1 = 32'd393
; 
32'd16162: dataIn1 = 32'd426
; 
32'd16163: dataIn1 = 32'd431
; 
32'd16164: dataIn1 = 32'd492
; 
32'd16165: dataIn1 = 32'd494
; 
32'd16166: dataIn1 = 32'd535
; 
32'd16167: dataIn1 = 32'd572
; 
32'd16168: dataIn1 = 32'd575
; 
32'd16169: dataIn1 = 32'd576
; 
32'd16170: dataIn1 = 32'd598
; 
32'd16171: dataIn1 = 32'd605
; 
32'd16172: dataIn1 = 32'd637
; 
32'd16173: dataIn1 = 32'd679
; 
32'd16174: dataIn1 = 32'd681
; 
32'd16175: dataIn1 = 32'd737
; 
32'd16176: dataIn1 = 32'd740
; 
32'd16177: dataIn1 = 32'd744
; 
32'd16178: dataIn1 = 32'd797
; 
32'd16179: dataIn1 = 32'd206
; 
32'd16180: dataIn1 = 32'd211
; 
32'd16181: dataIn1 = 32'd212
; 
32'd16182: dataIn1 = 32'd261
; 
32'd16183: dataIn1 = 32'd262
; 
32'd16184: dataIn1 = 32'd293
; 
32'd16185: dataIn1 = 32'd303
; 
32'd16186: dataIn1 = 32'd340
; 
32'd16187: dataIn1 = 32'd378
; 
32'd16188: dataIn1 = 32'd382
; 
32'd16189: dataIn1 = 32'd390
; 
32'd16190: dataIn1 = 32'd395
; 
32'd16191: dataIn1 = 32'd397
; 
32'd16192: dataIn1 = 32'd399
; 
32'd16193: dataIn1 = 32'd404
; 
32'd16194: dataIn1 = 32'd419
; 
32'd16195: dataIn1 = 32'd422
; 
32'd16196: dataIn1 = 32'd459
; 
32'd16197: dataIn1 = 32'd478
; 
32'd16198: dataIn1 = 32'd498
; 
32'd16199: dataIn1 = 32'd500
; 
32'd16200: dataIn1 = 32'd533
; 
32'd16201: dataIn1 = 32'd535
; 
32'd16202: dataIn1 = 32'd564
; 
32'd16203: dataIn1 = 32'd571
; 
32'd16204: dataIn1 = 32'd594
; 
32'd16205: dataIn1 = 32'd621
; 
32'd16206: dataIn1 = 32'd625
; 
32'd16207: dataIn1 = 32'd648
; 
32'd16208: dataIn1 = 32'd659
; 
32'd16209: dataIn1 = 32'd663
; 
32'd16210: dataIn1 = 32'd669
; 
32'd16211: dataIn1 = 32'd678
; 
32'd16212: dataIn1 = 32'd688
; 
32'd16213: dataIn1 = 32'd699
; 
32'd16214: dataIn1 = 32'd702
; 
32'd16215: dataIn1 = 32'd729
; 
32'd16216: dataIn1 = 32'd740
; 
32'd16217: dataIn1 = 32'd742
; 
32'd16218: dataIn1 = 32'd760
; 
32'd16219: dataIn1 = 32'd765
; 
32'd16220: dataIn1 = 32'd771
; 
32'd16221: dataIn1 = 32'd773
; 
32'd16222: dataIn1 = 32'd778
; 
32'd16223: dataIn1 = 32'd212
; 
32'd16224: dataIn1 = 32'd213
; 
32'd16225: dataIn1 = 32'd220
; 
32'd16226: dataIn1 = 32'd239
; 
32'd16227: dataIn1 = 32'd263
; 
32'd16228: dataIn1 = 32'd286
; 
32'd16229: dataIn1 = 32'd287
; 
32'd16230: dataIn1 = 32'd310
; 
32'd16231: dataIn1 = 32'd312
; 
32'd16232: dataIn1 = 32'd323
; 
32'd16233: dataIn1 = 32'd336
; 
32'd16234: dataIn1 = 32'd344
; 
32'd16235: dataIn1 = 32'd380
; 
32'd16236: dataIn1 = 32'd384
; 
32'd16237: dataIn1 = 32'd393
; 
32'd16238: dataIn1 = 32'd402
; 
32'd16239: dataIn1 = 32'd415
; 
32'd16240: dataIn1 = 32'd432
; 
32'd16241: dataIn1 = 32'd440
; 
32'd16242: dataIn1 = 32'd442
; 
32'd16243: dataIn1 = 32'd443
; 
32'd16244: dataIn1 = 32'd475
; 
32'd16245: dataIn1 = 32'd496
; 
32'd16246: dataIn1 = 32'd510
; 
32'd16247: dataIn1 = 32'd512
; 
32'd16248: dataIn1 = 32'd519
; 
32'd16249: dataIn1 = 32'd529
; 
32'd16250: dataIn1 = 32'd567
; 
32'd16251: dataIn1 = 32'd616
; 
32'd16252: dataIn1 = 32'd622
; 
32'd16253: dataIn1 = 32'd641
; 
32'd16254: dataIn1 = 32'd670
; 
32'd16255: dataIn1 = 32'd675
; 
32'd16256: dataIn1 = 32'd681
; 
32'd16257: dataIn1 = 32'd698
; 
32'd16258: dataIn1 = 32'd725
; 
32'd16259: dataIn1 = 32'd729
; 
32'd16260: dataIn1 = 32'd733
; 
32'd16261: dataIn1 = 32'd736
; 
32'd16262: dataIn1 = 32'd738
; 
32'd16263: dataIn1 = 32'd741
; 
32'd16264: dataIn1 = 32'd742
; 
32'd16265: dataIn1 = 32'd749
; 
32'd16266: dataIn1 = 32'd796
; 
32'd16267: dataIn1 = 32'd212
; 
32'd16268: dataIn1 = 32'd232
; 
32'd16269: dataIn1 = 32'd239
; 
32'd16270: dataIn1 = 32'd241
; 
32'd16271: dataIn1 = 32'd256
; 
32'd16272: dataIn1 = 32'd257
; 
32'd16273: dataIn1 = 32'd275
; 
32'd16274: dataIn1 = 32'd309
; 
32'd16275: dataIn1 = 32'd350
; 
32'd16276: dataIn1 = 32'd392
; 
32'd16277: dataIn1 = 32'd415
; 
32'd16278: dataIn1 = 32'd418
; 
32'd16279: dataIn1 = 32'd422
; 
32'd16280: dataIn1 = 32'd429
; 
32'd16281: dataIn1 = 32'd432
; 
32'd16282: dataIn1 = 32'd442
; 
32'd16283: dataIn1 = 32'd456
; 
32'd16284: dataIn1 = 32'd467
; 
32'd16285: dataIn1 = 32'd475
; 
32'd16286: dataIn1 = 32'd502
; 
32'd16287: dataIn1 = 32'd515
; 
32'd16288: dataIn1 = 32'd541
; 
32'd16289: dataIn1 = 32'd542
; 
32'd16290: dataIn1 = 32'd550
; 
32'd16291: dataIn1 = 32'd558
; 
32'd16292: dataIn1 = 32'd584
; 
32'd16293: dataIn1 = 32'd625
; 
32'd16294: dataIn1 = 32'd628
; 
32'd16295: dataIn1 = 32'd635
; 
32'd16296: dataIn1 = 32'd648
; 
32'd16297: dataIn1 = 32'd679
; 
32'd16298: dataIn1 = 32'd683
; 
32'd16299: dataIn1 = 32'd707
; 
32'd16300: dataIn1 = 32'd748
; 
32'd16301: dataIn1 = 32'd750
; 
32'd16302: dataIn1 = 32'd758
; 
32'd16303: dataIn1 = 32'd775
; 
32'd16304: dataIn1 = 32'd779
; 
32'd16305: dataIn1 = 32'd784
; 
32'd16306: dataIn1 = 32'd798
; 
32'd16307: dataIn1 = 32'd213
; 
32'd16308: dataIn1 = 32'd253
; 
32'd16309: dataIn1 = 32'd257
; 
32'd16310: dataIn1 = 32'd286
; 
32'd16311: dataIn1 = 32'd295
; 
32'd16312: dataIn1 = 32'd308
; 
32'd16313: dataIn1 = 32'd327
; 
32'd16314: dataIn1 = 32'd331
; 
32'd16315: dataIn1 = 32'd354
; 
32'd16316: dataIn1 = 32'd358
; 
32'd16317: dataIn1 = 32'd360
; 
32'd16318: dataIn1 = 32'd377
; 
32'd16319: dataIn1 = 32'd396
; 
32'd16320: dataIn1 = 32'd423
; 
32'd16321: dataIn1 = 32'd427
; 
32'd16322: dataIn1 = 32'd436
; 
32'd16323: dataIn1 = 32'd478
; 
32'd16324: dataIn1 = 32'd486
; 
32'd16325: dataIn1 = 32'd510
; 
32'd16326: dataIn1 = 32'd511
; 
32'd16327: dataIn1 = 32'd515
; 
32'd16328: dataIn1 = 32'd527
; 
32'd16329: dataIn1 = 32'd558
; 
32'd16330: dataIn1 = 32'd562
; 
32'd16331: dataIn1 = 32'd569
; 
32'd16332: dataIn1 = 32'd600
; 
32'd16333: dataIn1 = 32'd628
; 
32'd16334: dataIn1 = 32'd636
; 
32'd16335: dataIn1 = 32'd638
; 
32'd16336: dataIn1 = 32'd651
; 
32'd16337: dataIn1 = 32'd683
; 
32'd16338: dataIn1 = 32'd699
; 
32'd16339: dataIn1 = 32'd770
; 
32'd16340: dataIn1 = 32'd783
; 
32'd16341: dataIn1 = 32'd243
; 
32'd16342: dataIn1 = 32'd246
; 
32'd16343: dataIn1 = 32'd278
; 
32'd16344: dataIn1 = 32'd285
; 
32'd16345: dataIn1 = 32'd307
; 
32'd16346: dataIn1 = 32'd312
; 
32'd16347: dataIn1 = 32'd331
; 
32'd16348: dataIn1 = 32'd384
; 
32'd16349: dataIn1 = 32'd399
; 
32'd16350: dataIn1 = 32'd402
; 
32'd16351: dataIn1 = 32'd408
; 
32'd16352: dataIn1 = 32'd418
; 
32'd16353: dataIn1 = 32'd422
; 
32'd16354: dataIn1 = 32'd424
; 
32'd16355: dataIn1 = 32'd427
; 
32'd16356: dataIn1 = 32'd442
; 
32'd16357: dataIn1 = 32'd459
; 
32'd16358: dataIn1 = 32'd482
; 
32'd16359: dataIn1 = 32'd488
; 
32'd16360: dataIn1 = 32'd495
; 
32'd16361: dataIn1 = 32'd497
; 
32'd16362: dataIn1 = 32'd500
; 
32'd16363: dataIn1 = 32'd508
; 
32'd16364: dataIn1 = 32'd559
; 
32'd16365: dataIn1 = 32'd561
; 
32'd16366: dataIn1 = 32'd562
; 
32'd16367: dataIn1 = 32'd571
; 
32'd16368: dataIn1 = 32'd595
; 
32'd16369: dataIn1 = 32'd629
; 
32'd16370: dataIn1 = 32'd647
; 
32'd16371: dataIn1 = 32'd687
; 
32'd16372: dataIn1 = 32'd706
; 
32'd16373: dataIn1 = 32'd726
; 
32'd16374: dataIn1 = 32'd757
; 
32'd16375: dataIn1 = 32'd761
; 
32'd16376: dataIn1 = 32'd205
; 
32'd16377: dataIn1 = 32'd210
; 
32'd16378: dataIn1 = 32'd214
; 
32'd16379: dataIn1 = 32'd222
; 
32'd16380: dataIn1 = 32'd224
; 
32'd16381: dataIn1 = 32'd253
; 
32'd16382: dataIn1 = 32'd257
; 
32'd16383: dataIn1 = 32'd264
; 
32'd16384: dataIn1 = 32'd280
; 
32'd16385: dataIn1 = 32'd287
; 
32'd16386: dataIn1 = 32'd327
; 
32'd16387: dataIn1 = 32'd376
; 
32'd16388: dataIn1 = 32'd397
; 
32'd16389: dataIn1 = 32'd425
; 
32'd16390: dataIn1 = 32'd427
; 
32'd16391: dataIn1 = 32'd431
; 
32'd16392: dataIn1 = 32'd446
; 
32'd16393: dataIn1 = 32'd465
; 
32'd16394: dataIn1 = 32'd488
; 
32'd16395: dataIn1 = 32'd494
; 
32'd16396: dataIn1 = 32'd511
; 
32'd16397: dataIn1 = 32'd515
; 
32'd16398: dataIn1 = 32'd527
; 
32'd16399: dataIn1 = 32'd545
; 
32'd16400: dataIn1 = 32'd649
; 
32'd16401: dataIn1 = 32'd663
; 
32'd16402: dataIn1 = 32'd675
; 
32'd16403: dataIn1 = 32'd691
; 
32'd16404: dataIn1 = 32'd709
; 
32'd16405: dataIn1 = 32'd716
; 
32'd16406: dataIn1 = 32'd724
; 
32'd16407: dataIn1 = 32'd734
; 
32'd16408: dataIn1 = 32'd747
; 
32'd16409: dataIn1 = 32'd760
; 
32'd16410: dataIn1 = 32'd763
; 
32'd16411: dataIn1 = 32'd222
; 
32'd16412: dataIn1 = 32'd241
; 
32'd16413: dataIn1 = 32'd320
; 
32'd16414: dataIn1 = 32'd343
; 
32'd16415: dataIn1 = 32'd344
; 
32'd16416: dataIn1 = 32'd356
; 
32'd16417: dataIn1 = 32'd357
; 
32'd16418: dataIn1 = 32'd361
; 
32'd16419: dataIn1 = 32'd382
; 
32'd16420: dataIn1 = 32'd405
; 
32'd16421: dataIn1 = 32'd407
; 
32'd16422: dataIn1 = 32'd411
; 
32'd16423: dataIn1 = 32'd418
; 
32'd16424: dataIn1 = 32'd450
; 
32'd16425: dataIn1 = 32'd466
; 
32'd16426: dataIn1 = 32'd469
; 
32'd16427: dataIn1 = 32'd477
; 
32'd16428: dataIn1 = 32'd486
; 
32'd16429: dataIn1 = 32'd497
; 
32'd16430: dataIn1 = 32'd501
; 
32'd16431: dataIn1 = 32'd521
; 
32'd16432: dataIn1 = 32'd545
; 
32'd16433: dataIn1 = 32'd550
; 
32'd16434: dataIn1 = 32'd553
; 
32'd16435: dataIn1 = 32'd557
; 
32'd16436: dataIn1 = 32'd562
; 
32'd16437: dataIn1 = 32'd578
; 
32'd16438: dataIn1 = 32'd580
; 
32'd16439: dataIn1 = 32'd598
; 
32'd16440: dataIn1 = 32'd606
; 
32'd16441: dataIn1 = 32'd611
; 
32'd16442: dataIn1 = 32'd627
; 
32'd16443: dataIn1 = 32'd646
; 
32'd16444: dataIn1 = 32'd658
; 
32'd16445: dataIn1 = 32'd670
; 
32'd16446: dataIn1 = 32'd676
; 
32'd16447: dataIn1 = 32'd687
; 
32'd16448: dataIn1 = 32'd695
; 
32'd16449: dataIn1 = 32'd713
; 
32'd16450: dataIn1 = 32'd722
; 
32'd16451: dataIn1 = 32'd724
; 
32'd16452: dataIn1 = 32'd754
; 
32'd16453: dataIn1 = 32'd791
; 
32'd16454: dataIn1 = 32'd241
; 
32'd16455: dataIn1 = 32'd249
; 
32'd16456: dataIn1 = 32'd260
; 
32'd16457: dataIn1 = 32'd280
; 
32'd16458: dataIn1 = 32'd294
; 
32'd16459: dataIn1 = 32'd301
; 
32'd16460: dataIn1 = 32'd317
; 
32'd16461: dataIn1 = 32'd321
; 
32'd16462: dataIn1 = 32'd323
; 
32'd16463: dataIn1 = 32'd324
; 
32'd16464: dataIn1 = 32'd327
; 
32'd16465: dataIn1 = 32'd352
; 
32'd16466: dataIn1 = 32'd364
; 
32'd16467: dataIn1 = 32'd369
; 
32'd16468: dataIn1 = 32'd383
; 
32'd16469: dataIn1 = 32'd390
; 
32'd16470: dataIn1 = 32'd406
; 
32'd16471: dataIn1 = 32'd417
; 
32'd16472: dataIn1 = 32'd438
; 
32'd16473: dataIn1 = 32'd439
; 
32'd16474: dataIn1 = 32'd462
; 
32'd16475: dataIn1 = 32'd468
; 
32'd16476: dataIn1 = 32'd477
; 
32'd16477: dataIn1 = 32'd495
; 
32'd16478: dataIn1 = 32'd497
; 
32'd16479: dataIn1 = 32'd506
; 
32'd16480: dataIn1 = 32'd519
; 
32'd16481: dataIn1 = 32'd575
; 
32'd16482: dataIn1 = 32'd605
; 
32'd16483: dataIn1 = 32'd623
; 
32'd16484: dataIn1 = 32'd630
; 
32'd16485: dataIn1 = 32'd643
; 
32'd16486: dataIn1 = 32'd667
; 
32'd16487: dataIn1 = 32'd691
; 
32'd16488: dataIn1 = 32'd712
; 
32'd16489: dataIn1 = 32'd743
; 
32'd16490: dataIn1 = 32'd755
; 
32'd16491: dataIn1 = 32'd760
; 
32'd16492: dataIn1 = 32'd778
; 
32'd16493: dataIn1 = 32'd780
; 
32'd16494: dataIn1 = 32'd797
; 
32'd16495: dataIn1 = 32'd256
; 
32'd16496: dataIn1 = 32'd262
; 
32'd16497: dataIn1 = 32'd269
; 
32'd16498: dataIn1 = 32'd316
; 
32'd16499: dataIn1 = 32'd356
; 
32'd16500: dataIn1 = 32'd359
; 
32'd16501: dataIn1 = 32'd367
; 
32'd16502: dataIn1 = 32'd375
; 
32'd16503: dataIn1 = 32'd411
; 
32'd16504: dataIn1 = 32'd423
; 
32'd16505: dataIn1 = 32'd445
; 
32'd16506: dataIn1 = 32'd451
; 
32'd16507: dataIn1 = 32'd453
; 
32'd16508: dataIn1 = 32'd461
; 
32'd16509: dataIn1 = 32'd487
; 
32'd16510: dataIn1 = 32'd491
; 
32'd16511: dataIn1 = 32'd509
; 
32'd16512: dataIn1 = 32'd528
; 
32'd16513: dataIn1 = 32'd532
; 
32'd16514: dataIn1 = 32'd557
; 
32'd16515: dataIn1 = 32'd561
; 
32'd16516: dataIn1 = 32'd569
; 
32'd16517: dataIn1 = 32'd572
; 
32'd16518: dataIn1 = 32'd578
; 
32'd16519: dataIn1 = 32'd583
; 
32'd16520: dataIn1 = 32'd585
; 
32'd16521: dataIn1 = 32'd586
; 
32'd16522: dataIn1 = 32'd595
; 
32'd16523: dataIn1 = 32'd653
; 
32'd16524: dataIn1 = 32'd678
; 
32'd16525: dataIn1 = 32'd684
; 
32'd16526: dataIn1 = 32'd702
; 
32'd16527: dataIn1 = 32'd747
; 
32'd16528: dataIn1 = 32'd778
; 
32'd16529: dataIn1 = 32'd781
; 
32'd16530: dataIn1 = 32'd262
; 
32'd16531: dataIn1 = 32'd295
; 
32'd16532: dataIn1 = 32'd311
; 
32'd16533: dataIn1 = 32'd315
; 
32'd16534: dataIn1 = 32'd317
; 
32'd16535: dataIn1 = 32'd323
; 
32'd16536: dataIn1 = 32'd325
; 
32'd16537: dataIn1 = 32'd333
; 
32'd16538: dataIn1 = 32'd347
; 
32'd16539: dataIn1 = 32'd361
; 
32'd16540: dataIn1 = 32'd370
; 
32'd16541: dataIn1 = 32'd379
; 
32'd16542: dataIn1 = 32'd386
; 
32'd16543: dataIn1 = 32'd401
; 
32'd16544: dataIn1 = 32'd416
; 
32'd16545: dataIn1 = 32'd456
; 
32'd16546: dataIn1 = 32'd465
; 
32'd16547: dataIn1 = 32'd535
; 
32'd16548: dataIn1 = 32'd554
; 
32'd16549: dataIn1 = 32'd568
; 
32'd16550: dataIn1 = 32'd581
; 
32'd16551: dataIn1 = 32'd586
; 
32'd16552: dataIn1 = 32'd607
; 
32'd16553: dataIn1 = 32'd612
; 
32'd16554: dataIn1 = 32'd623
; 
32'd16555: dataIn1 = 32'd625
; 
32'd16556: dataIn1 = 32'd661
; 
32'd16557: dataIn1 = 32'd665
; 
32'd16558: dataIn1 = 32'd674
; 
32'd16559: dataIn1 = 32'd739
; 
32'd16560: dataIn1 = 32'd740
; 
32'd16561: dataIn1 = 32'd741
; 
32'd16562: dataIn1 = 32'd774
; 
32'd16563: dataIn1 = 32'd776
; 
32'd16564: dataIn1 = 32'd208
; 
32'd16565: dataIn1 = 32'd239
; 
32'd16566: dataIn1 = 32'd257
; 
32'd16567: dataIn1 = 32'd277
; 
32'd16568: dataIn1 = 32'd297
; 
32'd16569: dataIn1 = 32'd300
; 
32'd16570: dataIn1 = 32'd324
; 
32'd16571: dataIn1 = 32'd340
; 
32'd16572: dataIn1 = 32'd341
; 
32'd16573: dataIn1 = 32'd371
; 
32'd16574: dataIn1 = 32'd375
; 
32'd16575: dataIn1 = 32'd378
; 
32'd16576: dataIn1 = 32'd396
; 
32'd16577: dataIn1 = 32'd407
; 
32'd16578: dataIn1 = 32'd456
; 
32'd16579: dataIn1 = 32'd471
; 
32'd16580: dataIn1 = 32'd479
; 
32'd16581: dataIn1 = 32'd486
; 
32'd16582: dataIn1 = 32'd490
; 
32'd16583: dataIn1 = 32'd503
; 
32'd16584: dataIn1 = 32'd566
; 
32'd16585: dataIn1 = 32'd587
; 
32'd16586: dataIn1 = 32'd640
; 
32'd16587: dataIn1 = 32'd679
; 
32'd16588: dataIn1 = 32'd699
; 
32'd16589: dataIn1 = 32'd710
; 
32'd16590: dataIn1 = 32'd738
; 
32'd16591: dataIn1 = 32'd743
; 
32'd16592: dataIn1 = 32'd752
; 
32'd16593: dataIn1 = 32'd755
; 
32'd16594: dataIn1 = 32'd786
; 
32'd16595: dataIn1 = 32'd227
; 
32'd16596: dataIn1 = 32'd267
; 
32'd16597: dataIn1 = 32'd286
; 
32'd16598: dataIn1 = 32'd311
; 
32'd16599: dataIn1 = 32'd319
; 
32'd16600: dataIn1 = 32'd327
; 
32'd16601: dataIn1 = 32'd360
; 
32'd16602: dataIn1 = 32'd374
; 
32'd16603: dataIn1 = 32'd377
; 
32'd16604: dataIn1 = 32'd379
; 
32'd16605: dataIn1 = 32'd419
; 
32'd16606: dataIn1 = 32'd427
; 
32'd16607: dataIn1 = 32'd441
; 
32'd16608: dataIn1 = 32'd449
; 
32'd16609: dataIn1 = 32'd456
; 
32'd16610: dataIn1 = 32'd475
; 
32'd16611: dataIn1 = 32'd489
; 
32'd16612: dataIn1 = 32'd490
; 
32'd16613: dataIn1 = 32'd497
; 
32'd16614: dataIn1 = 32'd515
; 
32'd16615: dataIn1 = 32'd525
; 
32'd16616: dataIn1 = 32'd544
; 
32'd16617: dataIn1 = 32'd593
; 
32'd16618: dataIn1 = 32'd595
; 
32'd16619: dataIn1 = 32'd602
; 
32'd16620: dataIn1 = 32'd647
; 
32'd16621: dataIn1 = 32'd651
; 
32'd16622: dataIn1 = 32'd656
; 
32'd16623: dataIn1 = 32'd657
; 
32'd16624: dataIn1 = 32'd673
; 
32'd16625: dataIn1 = 32'd701
; 
32'd16626: dataIn1 = 32'd717
; 
32'd16627: dataIn1 = 32'd740
; 
32'd16628: dataIn1 = 32'd751
; 
32'd16629: dataIn1 = 32'd772
; 
32'd16630: dataIn1 = 32'd791
; 
32'd16631: dataIn1 = 32'd794
; 
32'd16632: dataIn1 = 32'd796
; 
32'd16633: dataIn1 = 32'd221
; 
32'd16634: dataIn1 = 32'd274
; 
32'd16635: dataIn1 = 32'd275
; 
32'd16636: dataIn1 = 32'd301
; 
32'd16637: dataIn1 = 32'd320
; 
32'd16638: dataIn1 = 32'd351
; 
32'd16639: dataIn1 = 32'd353
; 
32'd16640: dataIn1 = 32'd358
; 
32'd16641: dataIn1 = 32'd365
; 
32'd16642: dataIn1 = 32'd366
; 
32'd16643: dataIn1 = 32'd389
; 
32'd16644: dataIn1 = 32'd394
; 
32'd16645: dataIn1 = 32'd420
; 
32'd16646: dataIn1 = 32'd424
; 
32'd16647: dataIn1 = 32'd456
; 
32'd16648: dataIn1 = 32'd478
; 
32'd16649: dataIn1 = 32'd489
; 
32'd16650: dataIn1 = 32'd514
; 
32'd16651: dataIn1 = 32'd535
; 
32'd16652: dataIn1 = 32'd540
; 
32'd16653: dataIn1 = 32'd552
; 
32'd16654: dataIn1 = 32'd568
; 
32'd16655: dataIn1 = 32'd583
; 
32'd16656: dataIn1 = 32'd591
; 
32'd16657: dataIn1 = 32'd603
; 
32'd16658: dataIn1 = 32'd607
; 
32'd16659: dataIn1 = 32'd628
; 
32'd16660: dataIn1 = 32'd652
; 
32'd16661: dataIn1 = 32'd655
; 
32'd16662: dataIn1 = 32'd687
; 
32'd16663: dataIn1 = 32'd703
; 
32'd16664: dataIn1 = 32'd743
; 
32'd16665: dataIn1 = 32'd746
; 
32'd16666: dataIn1 = 32'd771
; 
32'd16667: dataIn1 = 32'd775
; 
32'd16668: dataIn1 = 32'd779
; 
32'd16669: dataIn1 = 32'd788
; 
32'd16670: dataIn1 = 32'd241
; 
32'd16671: dataIn1 = 32'd250
; 
32'd16672: dataIn1 = 32'd263
; 
32'd16673: dataIn1 = 32'd272
; 
32'd16674: dataIn1 = 32'd286
; 
32'd16675: dataIn1 = 32'd304
; 
32'd16676: dataIn1 = 32'd410
; 
32'd16677: dataIn1 = 32'd429
; 
32'd16678: dataIn1 = 32'd437
; 
32'd16679: dataIn1 = 32'd475
; 
32'd16680: dataIn1 = 32'd479
; 
32'd16681: dataIn1 = 32'd489
; 
32'd16682: dataIn1 = 32'd491
; 
32'd16683: dataIn1 = 32'd515
; 
32'd16684: dataIn1 = 32'd524
; 
32'd16685: dataIn1 = 32'd558
; 
32'd16686: dataIn1 = 32'd586
; 
32'd16687: dataIn1 = 32'd590
; 
32'd16688: dataIn1 = 32'd640
; 
32'd16689: dataIn1 = 32'd652
; 
32'd16690: dataIn1 = 32'd654
; 
32'd16691: dataIn1 = 32'd660
; 
32'd16692: dataIn1 = 32'd661
; 
32'd16693: dataIn1 = 32'd683
; 
32'd16694: dataIn1 = 32'd719
; 
32'd16695: dataIn1 = 32'd738
; 
32'd16696: dataIn1 = 32'd758
; 
32'd16697: dataIn1 = 32'd763
; 
32'd16698: dataIn1 = 32'd789
; 
32'd16699: dataIn1 = 32'd231
; 
32'd16700: dataIn1 = 32'd247
; 
32'd16701: dataIn1 = 32'd264
; 
32'd16702: dataIn1 = 32'd268
; 
32'd16703: dataIn1 = 32'd271
; 
32'd16704: dataIn1 = 32'd292
; 
32'd16705: dataIn1 = 32'd301
; 
32'd16706: dataIn1 = 32'd324
; 
32'd16707: dataIn1 = 32'd353
; 
32'd16708: dataIn1 = 32'd355
; 
32'd16709: dataIn1 = 32'd368
; 
32'd16710: dataIn1 = 32'd381
; 
32'd16711: dataIn1 = 32'd396
; 
32'd16712: dataIn1 = 32'd414
; 
32'd16713: dataIn1 = 32'd415
; 
32'd16714: dataIn1 = 32'd421
; 
32'd16715: dataIn1 = 32'd433
; 
32'd16716: dataIn1 = 32'd445
; 
32'd16717: dataIn1 = 32'd457
; 
32'd16718: dataIn1 = 32'd459
; 
32'd16719: dataIn1 = 32'd466
; 
32'd16720: dataIn1 = 32'd524
; 
32'd16721: dataIn1 = 32'd528
; 
32'd16722: dataIn1 = 32'd531
; 
32'd16723: dataIn1 = 32'd539
; 
32'd16724: dataIn1 = 32'd547
; 
32'd16725: dataIn1 = 32'd550
; 
32'd16726: dataIn1 = 32'd565
; 
32'd16727: dataIn1 = 32'd583
; 
32'd16728: dataIn1 = 32'd640
; 
32'd16729: dataIn1 = 32'd647
; 
32'd16730: dataIn1 = 32'd663
; 
32'd16731: dataIn1 = 32'd696
; 
32'd16732: dataIn1 = 32'd700
; 
32'd16733: dataIn1 = 32'd750
; 
32'd16734: dataIn1 = 32'd767
; 
32'd16735: dataIn1 = 32'd774
; 
32'd16736: dataIn1 = 32'd781
; 
32'd16737: dataIn1 = 32'd782
; 
32'd16738: dataIn1 = 32'd783
; 
32'd16739: dataIn1 = 32'd282
; 
32'd16740: dataIn1 = 32'd285
; 
32'd16741: dataIn1 = 32'd319
; 
32'd16742: dataIn1 = 32'd333
; 
32'd16743: dataIn1 = 32'd364
; 
32'd16744: dataIn1 = 32'd396
; 
32'd16745: dataIn1 = 32'd397
; 
32'd16746: dataIn1 = 32'd398
; 
32'd16747: dataIn1 = 32'd412
; 
32'd16748: dataIn1 = 32'd413
; 
32'd16749: dataIn1 = 32'd428
; 
32'd16750: dataIn1 = 32'd434
; 
32'd16751: dataIn1 = 32'd436
; 
32'd16752: dataIn1 = 32'd438
; 
32'd16753: dataIn1 = 32'd456
; 
32'd16754: dataIn1 = 32'd494
; 
32'd16755: dataIn1 = 32'd508
; 
32'd16756: dataIn1 = 32'd526
; 
32'd16757: dataIn1 = 32'd555
; 
32'd16758: dataIn1 = 32'd573
; 
32'd16759: dataIn1 = 32'd588
; 
32'd16760: dataIn1 = 32'd620
; 
32'd16761: dataIn1 = 32'd645
; 
32'd16762: dataIn1 = 32'd680
; 
32'd16763: dataIn1 = 32'd701
; 
32'd16764: dataIn1 = 32'd728
; 
32'd16765: dataIn1 = 32'd758
; 
32'd16766: dataIn1 = 32'd768
; 
32'd16767: dataIn1 = 32'd781
; 
32'd16768: dataIn1 = 32'd226
; 
32'd16769: dataIn1 = 32'd247
; 
32'd16770: dataIn1 = 32'd294
; 
32'd16771: dataIn1 = 32'd296
; 
32'd16772: dataIn1 = 32'd310
; 
32'd16773: dataIn1 = 32'd315
; 
32'd16774: dataIn1 = 32'd324
; 
32'd16775: dataIn1 = 32'd326
; 
32'd16776: dataIn1 = 32'd341
; 
32'd16777: dataIn1 = 32'd346
; 
32'd16778: dataIn1 = 32'd361
; 
32'd16779: dataIn1 = 32'd377
; 
32'd16780: dataIn1 = 32'd387
; 
32'd16781: dataIn1 = 32'd408
; 
32'd16782: dataIn1 = 32'd412
; 
32'd16783: dataIn1 = 32'd415
; 
32'd16784: dataIn1 = 32'd428
; 
32'd16785: dataIn1 = 32'd441
; 
32'd16786: dataIn1 = 32'd443
; 
32'd16787: dataIn1 = 32'd479
; 
32'd16788: dataIn1 = 32'd493
; 
32'd16789: dataIn1 = 32'd500
; 
32'd16790: dataIn1 = 32'd507
; 
32'd16791: dataIn1 = 32'd531
; 
32'd16792: dataIn1 = 32'd544
; 
32'd16793: dataIn1 = 32'd548
; 
32'd16794: dataIn1 = 32'd564
; 
32'd16795: dataIn1 = 32'd600
; 
32'd16796: dataIn1 = 32'd601
; 
32'd16797: dataIn1 = 32'd627
; 
32'd16798: dataIn1 = 32'd663
; 
32'd16799: dataIn1 = 32'd666
; 
32'd16800: dataIn1 = 32'd692
; 
32'd16801: dataIn1 = 32'd693
; 
32'd16802: dataIn1 = 32'd710
; 
32'd16803: dataIn1 = 32'd781
; 
32'd16804: dataIn1 = 32'd790
; 
32'd16805: dataIn1 = 32'd217
; 
32'd16806: dataIn1 = 32'd230
; 
32'd16807: dataIn1 = 32'd254
; 
32'd16808: dataIn1 = 32'd258
; 
32'd16809: dataIn1 = 32'd264
; 
32'd16810: dataIn1 = 32'd267
; 
32'd16811: dataIn1 = 32'd292
; 
32'd16812: dataIn1 = 32'd325
; 
32'd16813: dataIn1 = 32'd328
; 
32'd16814: dataIn1 = 32'd330
; 
32'd16815: dataIn1 = 32'd351
; 
32'd16816: dataIn1 = 32'd356
; 
32'd16817: dataIn1 = 32'd435
; 
32'd16818: dataIn1 = 32'd445
; 
32'd16819: dataIn1 = 32'd451
; 
32'd16820: dataIn1 = 32'd453
; 
32'd16821: dataIn1 = 32'd464
; 
32'd16822: dataIn1 = 32'd507
; 
32'd16823: dataIn1 = 32'd510
; 
32'd16824: dataIn1 = 32'd529
; 
32'd16825: dataIn1 = 32'd567
; 
32'd16826: dataIn1 = 32'd572
; 
32'd16827: dataIn1 = 32'd582
; 
32'd16828: dataIn1 = 32'd585
; 
32'd16829: dataIn1 = 32'd611
; 
32'd16830: dataIn1 = 32'd616
; 
32'd16831: dataIn1 = 32'd624
; 
32'd16832: dataIn1 = 32'd691
; 
32'd16833: dataIn1 = 32'd718
; 
32'd16834: dataIn1 = 32'd751
; 
32'd16835: dataIn1 = 32'd775
; 
32'd16836: dataIn1 = 32'd783
; 
32'd16837: dataIn1 = 32'd793
; 
32'd16838: dataIn1 = 32'd226
; 
32'd16839: dataIn1 = 32'd247
; 
32'd16840: dataIn1 = 32'd287
; 
32'd16841: dataIn1 = 32'd290
; 
32'd16842: dataIn1 = 32'd321
; 
32'd16843: dataIn1 = 32'd360
; 
32'd16844: dataIn1 = 32'd377
; 
32'd16845: dataIn1 = 32'd381
; 
32'd16846: dataIn1 = 32'd394
; 
32'd16847: dataIn1 = 32'd401
; 
32'd16848: dataIn1 = 32'd438
; 
32'd16849: dataIn1 = 32'd439
; 
32'd16850: dataIn1 = 32'd442
; 
32'd16851: dataIn1 = 32'd459
; 
32'd16852: dataIn1 = 32'd486
; 
32'd16853: dataIn1 = 32'd491
; 
32'd16854: dataIn1 = 32'd494
; 
32'd16855: dataIn1 = 32'd499
; 
32'd16856: dataIn1 = 32'd510
; 
32'd16857: dataIn1 = 32'd576
; 
32'd16858: dataIn1 = 32'd579
; 
32'd16859: dataIn1 = 32'd586
; 
32'd16860: dataIn1 = 32'd587
; 
32'd16861: dataIn1 = 32'd597
; 
32'd16862: dataIn1 = 32'd610
; 
32'd16863: dataIn1 = 32'd629
; 
32'd16864: dataIn1 = 32'd633
; 
32'd16865: dataIn1 = 32'd649
; 
32'd16866: dataIn1 = 32'd655
; 
32'd16867: dataIn1 = 32'd688
; 
32'd16868: dataIn1 = 32'd707
; 
32'd16869: dataIn1 = 32'd709
; 
32'd16870: dataIn1 = 32'd720
; 
32'd16871: dataIn1 = 32'd743
; 
32'd16872: dataIn1 = 32'd759
; 
32'd16873: dataIn1 = 32'd761
; 
32'd16874: dataIn1 = 32'd763
; 
32'd16875: dataIn1 = 32'd764
; 
32'd16876: dataIn1 = 32'd778
; 
32'd16877: dataIn1 = 32'd783
; 
32'd16878: dataIn1 = 32'd794
; 
32'd16879: dataIn1 = 32'd256
; 
32'd16880: dataIn1 = 32'd265
; 
32'd16881: dataIn1 = 32'd269
; 
32'd16882: dataIn1 = 32'd291
; 
32'd16883: dataIn1 = 32'd311
; 
32'd16884: dataIn1 = 32'd326
; 
32'd16885: dataIn1 = 32'd329
; 
32'd16886: dataIn1 = 32'd331
; 
32'd16887: dataIn1 = 32'd334
; 
32'd16888: dataIn1 = 32'd352
; 
32'd16889: dataIn1 = 32'd358
; 
32'd16890: dataIn1 = 32'd363
; 
32'd16891: dataIn1 = 32'd372
; 
32'd16892: dataIn1 = 32'd374
; 
32'd16893: dataIn1 = 32'd381
; 
32'd16894: dataIn1 = 32'd397
; 
32'd16895: dataIn1 = 32'd401
; 
32'd16896: dataIn1 = 32'd408
; 
32'd16897: dataIn1 = 32'd449
; 
32'd16898: dataIn1 = 32'd459
; 
32'd16899: dataIn1 = 32'd487
; 
32'd16900: dataIn1 = 32'd526
; 
32'd16901: dataIn1 = 32'd532
; 
32'd16902: dataIn1 = 32'd534
; 
32'd16903: dataIn1 = 32'd560
; 
32'd16904: dataIn1 = 32'd567
; 
32'd16905: dataIn1 = 32'd574
; 
32'd16906: dataIn1 = 32'd597
; 
32'd16907: dataIn1 = 32'd624
; 
32'd16908: dataIn1 = 32'd637
; 
32'd16909: dataIn1 = 32'd721
; 
32'd16910: dataIn1 = 32'd741
; 
32'd16911: dataIn1 = 32'd752
; 
32'd16912: dataIn1 = 32'd763
; 
32'd16913: dataIn1 = 32'd774
; 
32'd16914: dataIn1 = 32'd783
; 
32'd16915: dataIn1 = 32'd797
; 
32'd16916: dataIn1 = 32'd223
; 
32'd16917: dataIn1 = 32'd233
; 
32'd16918: dataIn1 = 32'd255
; 
32'd16919: dataIn1 = 32'd287
; 
32'd16920: dataIn1 = 32'd304
; 
32'd16921: dataIn1 = 32'd330
; 
32'd16922: dataIn1 = 32'd341
; 
32'd16923: dataIn1 = 32'd347
; 
32'd16924: dataIn1 = 32'd356
; 
32'd16925: dataIn1 = 32'd369
; 
32'd16926: dataIn1 = 32'd377
; 
32'd16927: dataIn1 = 32'd385
; 
32'd16928: dataIn1 = 32'd390
; 
32'd16929: dataIn1 = 32'd403
; 
32'd16930: dataIn1 = 32'd406
; 
32'd16931: dataIn1 = 32'd410
; 
32'd16932: dataIn1 = 32'd411
; 
32'd16933: dataIn1 = 32'd419
; 
32'd16934: dataIn1 = 32'd430
; 
32'd16935: dataIn1 = 32'd433
; 
32'd16936: dataIn1 = 32'd446
; 
32'd16937: dataIn1 = 32'd469
; 
32'd16938: dataIn1 = 32'd474
; 
32'd16939: dataIn1 = 32'd478
; 
32'd16940: dataIn1 = 32'd483
; 
32'd16941: dataIn1 = 32'd505
; 
32'd16942: dataIn1 = 32'd539
; 
32'd16943: dataIn1 = 32'd541
; 
32'd16944: dataIn1 = 32'd555
; 
32'd16945: dataIn1 = 32'd575
; 
32'd16946: dataIn1 = 32'd583
; 
32'd16947: dataIn1 = 32'd618
; 
32'd16948: dataIn1 = 32'd647
; 
32'd16949: dataIn1 = 32'd665
; 
32'd16950: dataIn1 = 32'd667
; 
32'd16951: dataIn1 = 32'd680
; 
32'd16952: dataIn1 = 32'd708
; 
32'd16953: dataIn1 = 32'd713
; 
32'd16954: dataIn1 = 32'd724
; 
32'd16955: dataIn1 = 32'd733
; 
32'd16956: dataIn1 = 32'd739
; 
32'd16957: dataIn1 = 32'd742
; 
32'd16958: dataIn1 = 32'd746
; 
32'd16959: dataIn1 = 32'd753
; 
32'd16960: dataIn1 = 32'd788
; 
32'd16961: dataIn1 = 32'd793
; 
32'd16962: dataIn1 = 32'd238
; 
32'd16963: dataIn1 = 32'd242
; 
32'd16964: dataIn1 = 32'd249
; 
32'd16965: dataIn1 = 32'd275
; 
32'd16966: dataIn1 = 32'd291
; 
32'd16967: dataIn1 = 32'd319
; 
32'd16968: dataIn1 = 32'd323
; 
32'd16969: dataIn1 = 32'd327
; 
32'd16970: dataIn1 = 32'd353
; 
32'd16971: dataIn1 = 32'd386
; 
32'd16972: dataIn1 = 32'd388
; 
32'd16973: dataIn1 = 32'd392
; 
32'd16974: dataIn1 = 32'd405
; 
32'd16975: dataIn1 = 32'd406
; 
32'd16976: dataIn1 = 32'd423
; 
32'd16977: dataIn1 = 32'd442
; 
32'd16978: dataIn1 = 32'd450
; 
32'd16979: dataIn1 = 32'd510
; 
32'd16980: dataIn1 = 32'd519
; 
32'd16981: dataIn1 = 32'd526
; 
32'd16982: dataIn1 = 32'd547
; 
32'd16983: dataIn1 = 32'd582
; 
32'd16984: dataIn1 = 32'd589
; 
32'd16985: dataIn1 = 32'd643
; 
32'd16986: dataIn1 = 32'd661
; 
32'd16987: dataIn1 = 32'd682
; 
32'd16988: dataIn1 = 32'd702
; 
32'd16989: dataIn1 = 32'd707
; 
32'd16990: dataIn1 = 32'd722
; 
32'd16991: dataIn1 = 32'd749
; 
32'd16992: dataIn1 = 32'd764
; 
32'd16993: dataIn1 = 32'd223
; 
32'd16994: dataIn1 = 32'd233
; 
32'd16995: dataIn1 = 32'd246
; 
32'd16996: dataIn1 = 32'd247
; 
32'd16997: dataIn1 = 32'd248
; 
32'd16998: dataIn1 = 32'd277
; 
32'd16999: dataIn1 = 32'd297
; 
32'd17000: dataIn1 = 32'd345
; 
32'd17001: dataIn1 = 32'd361
; 
32'd17002: dataIn1 = 32'd371
; 
32'd17003: dataIn1 = 32'd373
; 
32'd17004: dataIn1 = 32'd380
; 
32'd17005: dataIn1 = 32'd404
; 
32'd17006: dataIn1 = 32'd429
; 
32'd17007: dataIn1 = 32'd440
; 
32'd17008: dataIn1 = 32'd464
; 
32'd17009: dataIn1 = 32'd511
; 
32'd17010: dataIn1 = 32'd517
; 
32'd17011: dataIn1 = 32'd561
; 
32'd17012: dataIn1 = 32'd577
; 
32'd17013: dataIn1 = 32'd578
; 
32'd17014: dataIn1 = 32'd594
; 
32'd17015: dataIn1 = 32'd615
; 
32'd17016: dataIn1 = 32'd625
; 
32'd17017: dataIn1 = 32'd629
; 
32'd17018: dataIn1 = 32'd635
; 
32'd17019: dataIn1 = 32'd640
; 
32'd17020: dataIn1 = 32'd646
; 
32'd17021: dataIn1 = 32'd671
; 
32'd17022: dataIn1 = 32'd679
; 
32'd17023: dataIn1 = 32'd719
; 
32'd17024: dataIn1 = 32'd724
; 
32'd17025: dataIn1 = 32'd734
; 
32'd17026: dataIn1 = 32'd763
; 
32'd17027: dataIn1 = 32'd766
; 
32'd17028: dataIn1 = 32'd769
; 
32'd17029: dataIn1 = 32'd790
; 
32'd17030: dataIn1 = 32'd791
; 
32'd17031: dataIn1 = 32'd795
; 
32'd17032: dataIn1 = 32'd233
; 
32'd17033: dataIn1 = 32'd271
; 
32'd17034: dataIn1 = 32'd283
; 
32'd17035: dataIn1 = 32'd285
; 
32'd17036: dataIn1 = 32'd309
; 
32'd17037: dataIn1 = 32'd355
; 
32'd17038: dataIn1 = 32'd380
; 
32'd17039: dataIn1 = 32'd383
; 
32'd17040: dataIn1 = 32'd386
; 
32'd17041: dataIn1 = 32'd397
; 
32'd17042: dataIn1 = 32'd405
; 
32'd17043: dataIn1 = 32'd422
; 
32'd17044: dataIn1 = 32'd446
; 
32'd17045: dataIn1 = 32'd476
; 
32'd17046: dataIn1 = 32'd481
; 
32'd17047: dataIn1 = 32'd482
; 
32'd17048: dataIn1 = 32'd488
; 
32'd17049: dataIn1 = 32'd519
; 
32'd17050: dataIn1 = 32'd535
; 
32'd17051: dataIn1 = 32'd540
; 
32'd17052: dataIn1 = 32'd552
; 
32'd17053: dataIn1 = 32'd583
; 
32'd17054: dataIn1 = 32'd586
; 
32'd17055: dataIn1 = 32'd594
; 
32'd17056: dataIn1 = 32'd602
; 
32'd17057: dataIn1 = 32'd604
; 
32'd17058: dataIn1 = 32'd617
; 
32'd17059: dataIn1 = 32'd619
; 
32'd17060: dataIn1 = 32'd630
; 
32'd17061: dataIn1 = 32'd656
; 
32'd17062: dataIn1 = 32'd664
; 
32'd17063: dataIn1 = 32'd679
; 
32'd17064: dataIn1 = 32'd691
; 
32'd17065: dataIn1 = 32'd714
; 
32'd17066: dataIn1 = 32'd716
; 
32'd17067: dataIn1 = 32'd723
; 
32'd17068: dataIn1 = 32'd730
; 
32'd17069: dataIn1 = 32'd735
; 
32'd17070: dataIn1 = 32'd763
; 
32'd17071: dataIn1 = 32'd794
; 
32'd17072: dataIn1 = 32'd235
; 
32'd17073: dataIn1 = 32'd239
; 
32'd17074: dataIn1 = 32'd240
; 
32'd17075: dataIn1 = 32'd241
; 
32'd17076: dataIn1 = 32'd245
; 
32'd17077: dataIn1 = 32'd258
; 
32'd17078: dataIn1 = 32'd279
; 
32'd17079: dataIn1 = 32'd290
; 
32'd17080: dataIn1 = 32'd294
; 
32'd17081: dataIn1 = 32'd297
; 
32'd17082: dataIn1 = 32'd300
; 
32'd17083: dataIn1 = 32'd333
; 
32'd17084: dataIn1 = 32'd365
; 
32'd17085: dataIn1 = 32'd368
; 
32'd17086: dataIn1 = 32'd374
; 
32'd17087: dataIn1 = 32'd380
; 
32'd17088: dataIn1 = 32'd393
; 
32'd17089: dataIn1 = 32'd421
; 
32'd17090: dataIn1 = 32'd431
; 
32'd17091: dataIn1 = 32'd452
; 
32'd17092: dataIn1 = 32'd471
; 
32'd17093: dataIn1 = 32'd507
; 
32'd17094: dataIn1 = 32'd508
; 
32'd17095: dataIn1 = 32'd516
; 
32'd17096: dataIn1 = 32'd517
; 
32'd17097: dataIn1 = 32'd524
; 
32'd17098: dataIn1 = 32'd581
; 
32'd17099: dataIn1 = 32'd597
; 
32'd17100: dataIn1 = 32'd636
; 
32'd17101: dataIn1 = 32'd638
; 
32'd17102: dataIn1 = 32'd639
; 
32'd17103: dataIn1 = 32'd652
; 
32'd17104: dataIn1 = 32'd672
; 
32'd17105: dataIn1 = 32'd688
; 
32'd17106: dataIn1 = 32'd693
; 
32'd17107: dataIn1 = 32'd698
; 
32'd17108: dataIn1 = 32'd746
; 
32'd17109: dataIn1 = 32'd752
; 
32'd17110: dataIn1 = 32'd799
; 
32'd17111: dataIn1 = 32'd254
; 
32'd17112: dataIn1 = 32'd283
; 
32'd17113: dataIn1 = 32'd288
; 
32'd17114: dataIn1 = 32'd309
; 
32'd17115: dataIn1 = 32'd320
; 
32'd17116: dataIn1 = 32'd372
; 
32'd17117: dataIn1 = 32'd383
; 
32'd17118: dataIn1 = 32'd393
; 
32'd17119: dataIn1 = 32'd419
; 
32'd17120: dataIn1 = 32'd421
; 
32'd17121: dataIn1 = 32'd441
; 
32'd17122: dataIn1 = 32'd447
; 
32'd17123: dataIn1 = 32'd452
; 
32'd17124: dataIn1 = 32'd473
; 
32'd17125: dataIn1 = 32'd493
; 
32'd17126: dataIn1 = 32'd500
; 
32'd17127: dataIn1 = 32'd501
; 
32'd17128: dataIn1 = 32'd509
; 
32'd17129: dataIn1 = 32'd534
; 
32'd17130: dataIn1 = 32'd547
; 
32'd17131: dataIn1 = 32'd585
; 
32'd17132: dataIn1 = 32'd589
; 
32'd17133: dataIn1 = 32'd593
; 
32'd17134: dataIn1 = 32'd600
; 
32'd17135: dataIn1 = 32'd603
; 
32'd17136: dataIn1 = 32'd637
; 
32'd17137: dataIn1 = 32'd649
; 
32'd17138: dataIn1 = 32'd654
; 
32'd17139: dataIn1 = 32'd683
; 
32'd17140: dataIn1 = 32'd701
; 
32'd17141: dataIn1 = 32'd704
; 
32'd17142: dataIn1 = 32'd754
; 
32'd17143: dataIn1 = 32'd792
; 
32'd17144: dataIn1 = 32'd797
; 
32'd17145: dataIn1 = 32'd252
; 
32'd17146: dataIn1 = 32'd265
; 
32'd17147: dataIn1 = 32'd275
; 
32'd17148: dataIn1 = 32'd294
; 
32'd17149: dataIn1 = 32'd310
; 
32'd17150: dataIn1 = 32'd323
; 
32'd17151: dataIn1 = 32'd340
; 
32'd17152: dataIn1 = 32'd382
; 
32'd17153: dataIn1 = 32'd399
; 
32'd17154: dataIn1 = 32'd403
; 
32'd17155: dataIn1 = 32'd445
; 
32'd17156: dataIn1 = 32'd487
; 
32'd17157: dataIn1 = 32'd492
; 
32'd17158: dataIn1 = 32'd493
; 
32'd17159: dataIn1 = 32'd495
; 
32'd17160: dataIn1 = 32'd498
; 
32'd17161: dataIn1 = 32'd532
; 
32'd17162: dataIn1 = 32'd537
; 
32'd17163: dataIn1 = 32'd554
; 
32'd17164: dataIn1 = 32'd575
; 
32'd17165: dataIn1 = 32'd579
; 
32'd17166: dataIn1 = 32'd589
; 
32'd17167: dataIn1 = 32'd629
; 
32'd17168: dataIn1 = 32'd631
; 
32'd17169: dataIn1 = 32'd635
; 
32'd17170: dataIn1 = 32'd658
; 
32'd17171: dataIn1 = 32'd684
; 
32'd17172: dataIn1 = 32'd686
; 
32'd17173: dataIn1 = 32'd715
; 
32'd17174: dataIn1 = 32'd722
; 
32'd17175: dataIn1 = 32'd724
; 
32'd17176: dataIn1 = 32'd730
; 
32'd17177: dataIn1 = 32'd751
; 
32'd17178: dataIn1 = 32'd768
; 
32'd17179: dataIn1 = 32'd799
; 
32'd17180: dataIn1 = 32'd244
; 
32'd17181: dataIn1 = 32'd253
; 
32'd17182: dataIn1 = 32'd272
; 
32'd17183: dataIn1 = 32'd283
; 
32'd17184: dataIn1 = 32'd293
; 
32'd17185: dataIn1 = 32'd324
; 
32'd17186: dataIn1 = 32'd330
; 
32'd17187: dataIn1 = 32'd351
; 
32'd17188: dataIn1 = 32'd362
; 
32'd17189: dataIn1 = 32'd370
; 
32'd17190: dataIn1 = 32'd406
; 
32'd17191: dataIn1 = 32'd413
; 
32'd17192: dataIn1 = 32'd437
; 
32'd17193: dataIn1 = 32'd446
; 
32'd17194: dataIn1 = 32'd451
; 
32'd17195: dataIn1 = 32'd478
; 
32'd17196: dataIn1 = 32'd484
; 
32'd17197: dataIn1 = 32'd542
; 
32'd17198: dataIn1 = 32'd550
; 
32'd17199: dataIn1 = 32'd557
; 
32'd17200: dataIn1 = 32'd562
; 
32'd17201: dataIn1 = 32'd571
; 
32'd17202: dataIn1 = 32'd588
; 
32'd17203: dataIn1 = 32'd593
; 
32'd17204: dataIn1 = 32'd680
; 
32'd17205: dataIn1 = 32'd683
; 
32'd17206: dataIn1 = 32'd687
; 
32'd17207: dataIn1 = 32'd688
; 
32'd17208: dataIn1 = 32'd695
; 
32'd17209: dataIn1 = 32'd700
; 
32'd17210: dataIn1 = 32'd727
; 
32'd17211: dataIn1 = 32'd728
; 
32'd17212: dataIn1 = 32'd747
; 
32'd17213: dataIn1 = 32'd763
; 
32'd17214: dataIn1 = 32'd765
; 
32'd17215: dataIn1 = 32'd766
; 
32'd17216: dataIn1 = 32'd786
; 
32'd17217: dataIn1 = 32'd790
; 
32'd17218: dataIn1 = 32'd241
; 
32'd17219: dataIn1 = 32'd242
; 
32'd17220: dataIn1 = 32'd310
; 
32'd17221: dataIn1 = 32'd340
; 
32'd17222: dataIn1 = 32'd344
; 
32'd17223: dataIn1 = 32'd364
; 
32'd17224: dataIn1 = 32'd370
; 
32'd17225: dataIn1 = 32'd385
; 
32'd17226: dataIn1 = 32'd439
; 
32'd17227: dataIn1 = 32'd445
; 
32'd17228: dataIn1 = 32'd477
; 
32'd17229: dataIn1 = 32'd491
; 
32'd17230: dataIn1 = 32'd497
; 
32'd17231: dataIn1 = 32'd519
; 
32'd17232: dataIn1 = 32'd523
; 
32'd17233: dataIn1 = 32'd550
; 
32'd17234: dataIn1 = 32'd556
; 
32'd17235: dataIn1 = 32'd580
; 
32'd17236: dataIn1 = 32'd581
; 
32'd17237: dataIn1 = 32'd594
; 
32'd17238: dataIn1 = 32'd608
; 
32'd17239: dataIn1 = 32'd612
; 
32'd17240: dataIn1 = 32'd632
; 
32'd17241: dataIn1 = 32'd634
; 
32'd17242: dataIn1 = 32'd645
; 
32'd17243: dataIn1 = 32'd648
; 
32'd17244: dataIn1 = 32'd675
; 
32'd17245: dataIn1 = 32'd676
; 
32'd17246: dataIn1 = 32'd700
; 
32'd17247: dataIn1 = 32'd701
; 
32'd17248: dataIn1 = 32'd710
; 
32'd17249: dataIn1 = 32'd711
; 
32'd17250: dataIn1 = 32'd739
; 
32'd17251: dataIn1 = 32'd754
; 
32'd17252: dataIn1 = 32'd774
; 
32'd17253: dataIn1 = 32'd793
; 
32'd17254: dataIn1 = 32'd251
; 
32'd17255: dataIn1 = 32'd274
; 
32'd17256: dataIn1 = 32'd280
; 
32'd17257: dataIn1 = 32'd281
; 
32'd17258: dataIn1 = 32'd291
; 
32'd17259: dataIn1 = 32'd292
; 
32'd17260: dataIn1 = 32'd334
; 
32'd17261: dataIn1 = 32'd347
; 
32'd17262: dataIn1 = 32'd357
; 
32'd17263: dataIn1 = 32'd364
; 
32'd17264: dataIn1 = 32'd368
; 
32'd17265: dataIn1 = 32'd381
; 
32'd17266: dataIn1 = 32'd383
; 
32'd17267: dataIn1 = 32'd434
; 
32'd17268: dataIn1 = 32'd440
; 
32'd17269: dataIn1 = 32'd458
; 
32'd17270: dataIn1 = 32'd484
; 
32'd17271: dataIn1 = 32'd489
; 
32'd17272: dataIn1 = 32'd532
; 
32'd17273: dataIn1 = 32'd542
; 
32'd17274: dataIn1 = 32'd558
; 
32'd17275: dataIn1 = 32'd571
; 
32'd17276: dataIn1 = 32'd577
; 
32'd17277: dataIn1 = 32'd580
; 
32'd17278: dataIn1 = 32'd584
; 
32'd17279: dataIn1 = 32'd593
; 
32'd17280: dataIn1 = 32'd603
; 
32'd17281: dataIn1 = 32'd625
; 
32'd17282: dataIn1 = 32'd626
; 
32'd17283: dataIn1 = 32'd640
; 
32'd17284: dataIn1 = 32'd651
; 
32'd17285: dataIn1 = 32'd666
; 
32'd17286: dataIn1 = 32'd704
; 
32'd17287: dataIn1 = 32'd731
; 
32'd17288: dataIn1 = 32'd762
; 
32'd17289: dataIn1 = 32'd768
; 
32'd17290: dataIn1 = 32'd793
; 
32'd17291: dataIn1 = 32'd231
; 
32'd17292: dataIn1 = 32'd232
; 
32'd17293: dataIn1 = 32'd234
; 
32'd17294: dataIn1 = 32'd239
; 
32'd17295: dataIn1 = 32'd243
; 
32'd17296: dataIn1 = 32'd244
; 
32'd17297: dataIn1 = 32'd263
; 
32'd17298: dataIn1 = 32'd264
; 
32'd17299: dataIn1 = 32'd314
; 
32'd17300: dataIn1 = 32'd320
; 
32'd17301: dataIn1 = 32'd321
; 
32'd17302: dataIn1 = 32'd340
; 
32'd17303: dataIn1 = 32'd346
; 
32'd17304: dataIn1 = 32'd354
; 
32'd17305: dataIn1 = 32'd356
; 
32'd17306: dataIn1 = 32'd365
; 
32'd17307: dataIn1 = 32'd376
; 
32'd17308: dataIn1 = 32'd387
; 
32'd17309: dataIn1 = 32'd403
; 
32'd17310: dataIn1 = 32'd411
; 
32'd17311: dataIn1 = 32'd416
; 
32'd17312: dataIn1 = 32'd427
; 
32'd17313: dataIn1 = 32'd431
; 
32'd17314: dataIn1 = 32'd432
; 
32'd17315: dataIn1 = 32'd453
; 
32'd17316: dataIn1 = 32'd454
; 
32'd17317: dataIn1 = 32'd474
; 
32'd17318: dataIn1 = 32'd495
; 
32'd17319: dataIn1 = 32'd508
; 
32'd17320: dataIn1 = 32'd514
; 
32'd17321: dataIn1 = 32'd524
; 
32'd17322: dataIn1 = 32'd534
; 
32'd17323: dataIn1 = 32'd538
; 
32'd17324: dataIn1 = 32'd543
; 
32'd17325: dataIn1 = 32'd558
; 
32'd17326: dataIn1 = 32'd597
; 
32'd17327: dataIn1 = 32'd612
; 
32'd17328: dataIn1 = 32'd623
; 
32'd17329: dataIn1 = 32'd631
; 
32'd17330: dataIn1 = 32'd653
; 
32'd17331: dataIn1 = 32'd678
; 
32'd17332: dataIn1 = 32'd685
; 
32'd17333: dataIn1 = 32'd689
; 
32'd17334: dataIn1 = 32'd698
; 
32'd17335: dataIn1 = 32'd735
; 
32'd17336: dataIn1 = 32'd737
; 
32'd17337: dataIn1 = 32'd743
; 
32'd17338: dataIn1 = 32'd746
; 
32'd17339: dataIn1 = 32'd768
; 
32'd17340: dataIn1 = 32'd785
; 
32'd17341: dataIn1 = 32'd245
; 
32'd17342: dataIn1 = 32'd247
; 
32'd17343: dataIn1 = 32'd258
; 
32'd17344: dataIn1 = 32'd265
; 
32'd17345: dataIn1 = 32'd270
; 
32'd17346: dataIn1 = 32'd284
; 
32'd17347: dataIn1 = 32'd290
; 
32'd17348: dataIn1 = 32'd301
; 
32'd17349: dataIn1 = 32'd323
; 
32'd17350: dataIn1 = 32'd343
; 
32'd17351: dataIn1 = 32'd352
; 
32'd17352: dataIn1 = 32'd373
; 
32'd17353: dataIn1 = 32'd390
; 
32'd17354: dataIn1 = 32'd429
; 
32'd17355: dataIn1 = 32'd440
; 
32'd17356: dataIn1 = 32'd442
; 
32'd17357: dataIn1 = 32'd444
; 
32'd17358: dataIn1 = 32'd447
; 
32'd17359: dataIn1 = 32'd450
; 
32'd17360: dataIn1 = 32'd466
; 
32'd17361: dataIn1 = 32'd531
; 
32'd17362: dataIn1 = 32'd610
; 
32'd17363: dataIn1 = 32'd638
; 
32'd17364: dataIn1 = 32'd646
; 
32'd17365: dataIn1 = 32'd653
; 
32'd17366: dataIn1 = 32'd673
; 
32'd17367: dataIn1 = 32'd737
; 
32'd17368: dataIn1 = 32'd742
; 
32'd17369: dataIn1 = 32'd746
; 
32'd17370: dataIn1 = 32'd748
; 
32'd17371: dataIn1 = 32'd757
; 
32'd17372: dataIn1 = 32'd759
; 
32'd17373: dataIn1 = 32'd764
; 
32'd17374: dataIn1 = 32'd788
; 
32'd17375: dataIn1 = 32'd264
; 
32'd17376: dataIn1 = 32'd266
; 
32'd17377: dataIn1 = 32'd276
; 
32'd17378: dataIn1 = 32'd303
; 
32'd17379: dataIn1 = 32'd317
; 
32'd17380: dataIn1 = 32'd334
; 
32'd17381: dataIn1 = 32'd345
; 
32'd17382: dataIn1 = 32'd351
; 
32'd17383: dataIn1 = 32'd379
; 
32'd17384: dataIn1 = 32'd381
; 
32'd17385: dataIn1 = 32'd408
; 
32'd17386: dataIn1 = 32'd426
; 
32'd17387: dataIn1 = 32'd436
; 
32'd17388: dataIn1 = 32'd450
; 
32'd17389: dataIn1 = 32'd466
; 
32'd17390: dataIn1 = 32'd475
; 
32'd17391: dataIn1 = 32'd504
; 
32'd17392: dataIn1 = 32'd572
; 
32'd17393: dataIn1 = 32'd594
; 
32'd17394: dataIn1 = 32'd608
; 
32'd17395: dataIn1 = 32'd622
; 
32'd17396: dataIn1 = 32'd625
; 
32'd17397: dataIn1 = 32'd637
; 
32'd17398: dataIn1 = 32'd721
; 
32'd17399: dataIn1 = 32'd731
; 
32'd17400: dataIn1 = 32'd735
; 
32'd17401: dataIn1 = 32'd749
; 
32'd17402: dataIn1 = 32'd753
; 
32'd17403: dataIn1 = 32'd758
; 
32'd17404: dataIn1 = 32'd254
; 
32'd17405: dataIn1 = 32'd266
; 
32'd17406: dataIn1 = 32'd305
; 
32'd17407: dataIn1 = 32'd319
; 
32'd17408: dataIn1 = 32'd340
; 
32'd17409: dataIn1 = 32'd348
; 
32'd17410: dataIn1 = 32'd401
; 
32'd17411: dataIn1 = 32'd402
; 
32'd17412: dataIn1 = 32'd403
; 
32'd17413: dataIn1 = 32'd409
; 
32'd17414: dataIn1 = 32'd451
; 
32'd17415: dataIn1 = 32'd469
; 
32'd17416: dataIn1 = 32'd474
; 
32'd17417: dataIn1 = 32'd480
; 
32'd17418: dataIn1 = 32'd497
; 
32'd17419: dataIn1 = 32'd501
; 
32'd17420: dataIn1 = 32'd512
; 
32'd17421: dataIn1 = 32'd513
; 
32'd17422: dataIn1 = 32'd523
; 
32'd17423: dataIn1 = 32'd567
; 
32'd17424: dataIn1 = 32'd584
; 
32'd17425: dataIn1 = 32'd585
; 
32'd17426: dataIn1 = 32'd593
; 
32'd17427: dataIn1 = 32'd599
; 
32'd17428: dataIn1 = 32'd602
; 
32'd17429: dataIn1 = 32'd604
; 
32'd17430: dataIn1 = 32'd605
; 
32'd17431: dataIn1 = 32'd620
; 
32'd17432: dataIn1 = 32'd622
; 
32'd17433: dataIn1 = 32'd650
; 
32'd17434: dataIn1 = 32'd660
; 
32'd17435: dataIn1 = 32'd745
; 
32'd17436: dataIn1 = 32'd763
; 
32'd17437: dataIn1 = 32'd768
; 
32'd17438: dataIn1 = 32'd774
; 
32'd17439: dataIn1 = 32'd789
; 
32'd17440: dataIn1 = 32'd244
; 
32'd17441: dataIn1 = 32'd286
; 
32'd17442: dataIn1 = 32'd335
; 
32'd17443: dataIn1 = 32'd343
; 
32'd17444: dataIn1 = 32'd394
; 
32'd17445: dataIn1 = 32'd413
; 
32'd17446: dataIn1 = 32'd423
; 
32'd17447: dataIn1 = 32'd431
; 
32'd17448: dataIn1 = 32'd443
; 
32'd17449: dataIn1 = 32'd458
; 
32'd17450: dataIn1 = 32'd459
; 
32'd17451: dataIn1 = 32'd462
; 
32'd17452: dataIn1 = 32'd464
; 
32'd17453: dataIn1 = 32'd474
; 
32'd17454: dataIn1 = 32'd484
; 
32'd17455: dataIn1 = 32'd487
; 
32'd17456: dataIn1 = 32'd531
; 
32'd17457: dataIn1 = 32'd640
; 
32'd17458: dataIn1 = 32'd685
; 
32'd17459: dataIn1 = 32'd715
; 
32'd17460: dataIn1 = 32'd716
; 
32'd17461: dataIn1 = 32'd718
; 
32'd17462: dataIn1 = 32'd739
; 
32'd17463: dataIn1 = 32'd747
; 
32'd17464: dataIn1 = 32'd774
; 
32'd17465: dataIn1 = 32'd777
; 
32'd17466: dataIn1 = 32'd785
; 
32'd17467: dataIn1 = 32'd794
; 
32'd17468: dataIn1 = 32'd247
; 
32'd17469: dataIn1 = 32'd253
; 
32'd17470: dataIn1 = 32'd274
; 
32'd17471: dataIn1 = 32'd282
; 
32'd17472: dataIn1 = 32'd307
; 
32'd17473: dataIn1 = 32'd319
; 
32'd17474: dataIn1 = 32'd329
; 
32'd17475: dataIn1 = 32'd364
; 
32'd17476: dataIn1 = 32'd366
; 
32'd17477: dataIn1 = 32'd377
; 
32'd17478: dataIn1 = 32'd387
; 
32'd17479: dataIn1 = 32'd395
; 
32'd17480: dataIn1 = 32'd408
; 
32'd17481: dataIn1 = 32'd412
; 
32'd17482: dataIn1 = 32'd433
; 
32'd17483: dataIn1 = 32'd434
; 
32'd17484: dataIn1 = 32'd445
; 
32'd17485: dataIn1 = 32'd451
; 
32'd17486: dataIn1 = 32'd460
; 
32'd17487: dataIn1 = 32'd474
; 
32'd17488: dataIn1 = 32'd475
; 
32'd17489: dataIn1 = 32'd486
; 
32'd17490: dataIn1 = 32'd495
; 
32'd17491: dataIn1 = 32'd498
; 
32'd17492: dataIn1 = 32'd501
; 
32'd17493: dataIn1 = 32'd510
; 
32'd17494: dataIn1 = 32'd524
; 
32'd17495: dataIn1 = 32'd530
; 
32'd17496: dataIn1 = 32'd541
; 
32'd17497: dataIn1 = 32'd543
; 
32'd17498: dataIn1 = 32'd550
; 
32'd17499: dataIn1 = 32'd561
; 
32'd17500: dataIn1 = 32'd580
; 
32'd17501: dataIn1 = 32'd587
; 
32'd17502: dataIn1 = 32'd603
; 
32'd17503: dataIn1 = 32'd604
; 
32'd17504: dataIn1 = 32'd614
; 
32'd17505: dataIn1 = 32'd622
; 
32'd17506: dataIn1 = 32'd630
; 
32'd17507: dataIn1 = 32'd631
; 
32'd17508: dataIn1 = 32'd634
; 
32'd17509: dataIn1 = 32'd660
; 
32'd17510: dataIn1 = 32'd671
; 
32'd17511: dataIn1 = 32'd695
; 
32'd17512: dataIn1 = 32'd702
; 
32'd17513: dataIn1 = 32'd728
; 
32'd17514: dataIn1 = 32'd752
; 
32'd17515: dataIn1 = 32'd772
; 
32'd17516: dataIn1 = 32'd777
; 
32'd17517: dataIn1 = 32'd778
; 
32'd17518: dataIn1 = 32'd786
; 
32'd17519: dataIn1 = 32'd796
; 
32'd17520: dataIn1 = 32'd246
; 
32'd17521: dataIn1 = 32'd259
; 
32'd17522: dataIn1 = 32'd272
; 
32'd17523: dataIn1 = 32'd312
; 
32'd17524: dataIn1 = 32'd324
; 
32'd17525: dataIn1 = 32'd335
; 
32'd17526: dataIn1 = 32'd337
; 
32'd17527: dataIn1 = 32'd347
; 
32'd17528: dataIn1 = 32'd365
; 
32'd17529: dataIn1 = 32'd372
; 
32'd17530: dataIn1 = 32'd395
; 
32'd17531: dataIn1 = 32'd416
; 
32'd17532: dataIn1 = 32'd425
; 
32'd17533: dataIn1 = 32'd467
; 
32'd17534: dataIn1 = 32'd492
; 
32'd17535: dataIn1 = 32'd497
; 
32'd17536: dataIn1 = 32'd500
; 
32'd17537: dataIn1 = 32'd561
; 
32'd17538: dataIn1 = 32'd595
; 
32'd17539: dataIn1 = 32'd647
; 
32'd17540: dataIn1 = 32'd663
; 
32'd17541: dataIn1 = 32'd682
; 
32'd17542: dataIn1 = 32'd693
; 
32'd17543: dataIn1 = 32'd695
; 
32'd17544: dataIn1 = 32'd734
; 
32'd17545: dataIn1 = 32'd767
; 
32'd17546: dataIn1 = 32'd789
; 
32'd17547: dataIn1 = 32'd795
; 
32'd17548: dataIn1 = 32'd242
; 
32'd17549: dataIn1 = 32'd253
; 
32'd17550: dataIn1 = 32'd260
; 
32'd17551: dataIn1 = 32'd262
; 
32'd17552: dataIn1 = 32'd316
; 
32'd17553: dataIn1 = 32'd332
; 
32'd17554: dataIn1 = 32'd333
; 
32'd17555: dataIn1 = 32'd360
; 
32'd17556: dataIn1 = 32'd386
; 
32'd17557: dataIn1 = 32'd404
; 
32'd17558: dataIn1 = 32'd409
; 
32'd17559: dataIn1 = 32'd410
; 
32'd17560: dataIn1 = 32'd438
; 
32'd17561: dataIn1 = 32'd487
; 
32'd17562: dataIn1 = 32'd496
; 
32'd17563: dataIn1 = 32'd545
; 
32'd17564: dataIn1 = 32'd577
; 
32'd17565: dataIn1 = 32'd607
; 
32'd17566: dataIn1 = 32'd614
; 
32'd17567: dataIn1 = 32'd622
; 
32'd17568: dataIn1 = 32'd628
; 
32'd17569: dataIn1 = 32'd633
; 
32'd17570: dataIn1 = 32'd665
; 
32'd17571: dataIn1 = 32'd675
; 
32'd17572: dataIn1 = 32'd682
; 
32'd17573: dataIn1 = 32'd688
; 
32'd17574: dataIn1 = 32'd716
; 
32'd17575: dataIn1 = 32'd720
; 
32'd17576: dataIn1 = 32'd726
; 
32'd17577: dataIn1 = 32'd737
; 
32'd17578: dataIn1 = 32'd740
; 
32'd17579: dataIn1 = 32'd780
; 
32'd17580: dataIn1 = 32'd254
; 
32'd17581: dataIn1 = 32'd263
; 
32'd17582: dataIn1 = 32'd266
; 
32'd17583: dataIn1 = 32'd285
; 
32'd17584: dataIn1 = 32'd291
; 
32'd17585: dataIn1 = 32'd336
; 
32'd17586: dataIn1 = 32'd358
; 
32'd17587: dataIn1 = 32'd364
; 
32'd17588: dataIn1 = 32'd392
; 
32'd17589: dataIn1 = 32'd411
; 
32'd17590: dataIn1 = 32'd415
; 
32'd17591: dataIn1 = 32'd428
; 
32'd17592: dataIn1 = 32'd520
; 
32'd17593: dataIn1 = 32'd549
; 
32'd17594: dataIn1 = 32'd555
; 
32'd17595: dataIn1 = 32'd628
; 
32'd17596: dataIn1 = 32'd635
; 
32'd17597: dataIn1 = 32'd638
; 
32'd17598: dataIn1 = 32'd640
; 
32'd17599: dataIn1 = 32'd646
; 
32'd17600: dataIn1 = 32'd654
; 
32'd17601: dataIn1 = 32'd666
; 
32'd17602: dataIn1 = 32'd685
; 
32'd17603: dataIn1 = 32'd692
; 
32'd17604: dataIn1 = 32'd736
; 
32'd17605: dataIn1 = 32'd738
; 
32'd17606: dataIn1 = 32'd739
; 
32'd17607: dataIn1 = 32'd746
; 
32'd17608: dataIn1 = 32'd748
; 
32'd17609: dataIn1 = 32'd758
; 
32'd17610: dataIn1 = 32'd760
; 
32'd17611: dataIn1 = 32'd777
; 
32'd17612: dataIn1 = 32'd787
; 
32'd17613: dataIn1 = 32'd261
; 
32'd17614: dataIn1 = 32'd285
; 
32'd17615: dataIn1 = 32'd296
; 
32'd17616: dataIn1 = 32'd311
; 
32'd17617: dataIn1 = 32'd325
; 
32'd17618: dataIn1 = 32'd328
; 
32'd17619: dataIn1 = 32'd351
; 
32'd17620: dataIn1 = 32'd372
; 
32'd17621: dataIn1 = 32'd392
; 
32'd17622: dataIn1 = 32'd412
; 
32'd17623: dataIn1 = 32'd423
; 
32'd17624: dataIn1 = 32'd431
; 
32'd17625: dataIn1 = 32'd435
; 
32'd17626: dataIn1 = 32'd465
; 
32'd17627: dataIn1 = 32'd467
; 
32'd17628: dataIn1 = 32'd491
; 
32'd17629: dataIn1 = 32'd574
; 
32'd17630: dataIn1 = 32'd611
; 
32'd17631: dataIn1 = 32'd616
; 
32'd17632: dataIn1 = 32'd624
; 
32'd17633: dataIn1 = 32'd668
; 
32'd17634: dataIn1 = 32'd669
; 
32'd17635: dataIn1 = 32'd672
; 
32'd17636: dataIn1 = 32'd678
; 
32'd17637: dataIn1 = 32'd692
; 
32'd17638: dataIn1 = 32'd700
; 
32'd17639: dataIn1 = 32'd705
; 
32'd17640: dataIn1 = 32'd786
; 
32'd17641: dataIn1 = 32'd252
; 
32'd17642: dataIn1 = 32'd254
; 
32'd17643: dataIn1 = 32'd284
; 
32'd17644: dataIn1 = 32'd295
; 
32'd17645: dataIn1 = 32'd301
; 
32'd17646: dataIn1 = 32'd344
; 
32'd17647: dataIn1 = 32'd345
; 
32'd17648: dataIn1 = 32'd353
; 
32'd17649: dataIn1 = 32'd372
; 
32'd17650: dataIn1 = 32'd384
; 
32'd17651: dataIn1 = 32'd402
; 
32'd17652: dataIn1 = 32'd428
; 
32'd17653: dataIn1 = 32'd451
; 
32'd17654: dataIn1 = 32'd463
; 
32'd17655: dataIn1 = 32'd472
; 
32'd17656: dataIn1 = 32'd503
; 
32'd17657: dataIn1 = 32'd511
; 
32'd17658: dataIn1 = 32'd530
; 
32'd17659: dataIn1 = 32'd544
; 
32'd17660: dataIn1 = 32'd551
; 
32'd17661: dataIn1 = 32'd565
; 
32'd17662: dataIn1 = 32'd567
; 
32'd17663: dataIn1 = 32'd617
; 
32'd17664: dataIn1 = 32'd630
; 
32'd17665: dataIn1 = 32'd636
; 
32'd17666: dataIn1 = 32'd653
; 
32'd17667: dataIn1 = 32'd679
; 
32'd17668: dataIn1 = 32'd683
; 
32'd17669: dataIn1 = 32'd685
; 
32'd17670: dataIn1 = 32'd706
; 
32'd17671: dataIn1 = 32'd729
; 
32'd17672: dataIn1 = 32'd744
; 
32'd17673: dataIn1 = 32'd775
; 
32'd17674: dataIn1 = 32'd778
; 
32'd17675: dataIn1 = 32'd782
; 
32'd17676: dataIn1 = 32'd790
; 
32'd17677: dataIn1 = 32'd800
; 
32'd17678: dataIn1 = 32'd261
; 
32'd17679: dataIn1 = 32'd269
; 
32'd17680: dataIn1 = 32'd271
; 
32'd17681: dataIn1 = 32'd284
; 
32'd17682: dataIn1 = 32'd375
; 
32'd17683: dataIn1 = 32'd379
; 
32'd17684: dataIn1 = 32'd386
; 
32'd17685: dataIn1 = 32'd397
; 
32'd17686: dataIn1 = 32'd402
; 
32'd17687: dataIn1 = 32'd415
; 
32'd17688: dataIn1 = 32'd450
; 
32'd17689: dataIn1 = 32'd465
; 
32'd17690: dataIn1 = 32'd513
; 
32'd17691: dataIn1 = 32'd542
; 
32'd17692: dataIn1 = 32'd547
; 
32'd17693: dataIn1 = 32'd575
; 
32'd17694: dataIn1 = 32'd581
; 
32'd17695: dataIn1 = 32'd582
; 
32'd17696: dataIn1 = 32'd603
; 
32'd17697: dataIn1 = 32'd643
; 
32'd17698: dataIn1 = 32'd680
; 
32'd17699: dataIn1 = 32'd681
; 
32'd17700: dataIn1 = 32'd682
; 
32'd17701: dataIn1 = 32'd698
; 
32'd17702: dataIn1 = 32'd705
; 
32'd17703: dataIn1 = 32'd714
; 
32'd17704: dataIn1 = 32'd723
; 
32'd17705: dataIn1 = 32'd744
; 
32'd17706: dataIn1 = 32'd759
; 
32'd17707: dataIn1 = 32'd763
; 
32'd17708: dataIn1 = 32'd782
; 
32'd17709: dataIn1 = 32'd792
; 
32'd17710: dataIn1 = 32'd793
; 
32'd17711: dataIn1 = 32'd286
; 
32'd17712: dataIn1 = 32'd296
; 
32'd17713: dataIn1 = 32'd303
; 
32'd17714: dataIn1 = 32'd341
; 
32'd17715: dataIn1 = 32'd376
; 
32'd17716: dataIn1 = 32'd423
; 
32'd17717: dataIn1 = 32'd431
; 
32'd17718: dataIn1 = 32'd487
; 
32'd17719: dataIn1 = 32'd504
; 
32'd17720: dataIn1 = 32'd518
; 
32'd17721: dataIn1 = 32'd525
; 
32'd17722: dataIn1 = 32'd549
; 
32'd17723: dataIn1 = 32'd573
; 
32'd17724: dataIn1 = 32'd637
; 
32'd17725: dataIn1 = 32'd655
; 
32'd17726: dataIn1 = 32'd666
; 
32'd17727: dataIn1 = 32'd694
; 
32'd17728: dataIn1 = 32'd697
; 
32'd17729: dataIn1 = 32'd729
; 
32'd17730: dataIn1 = 32'd738
; 
32'd17731: dataIn1 = 32'd759
; 
32'd17732: dataIn1 = 32'd761
; 
32'd17733: dataIn1 = 32'd769
; 
32'd17734: dataIn1 = 32'd788
; 
32'd17735: dataIn1 = 32'd269
; 
32'd17736: dataIn1 = 32'd285
; 
32'd17737: dataIn1 = 32'd286
; 
32'd17738: dataIn1 = 32'd312
; 
32'd17739: dataIn1 = 32'd354
; 
32'd17740: dataIn1 = 32'd383
; 
32'd17741: dataIn1 = 32'd418
; 
32'd17742: dataIn1 = 32'd422
; 
32'd17743: dataIn1 = 32'd436
; 
32'd17744: dataIn1 = 32'd442
; 
32'd17745: dataIn1 = 32'd443
; 
32'd17746: dataIn1 = 32'd449
; 
32'd17747: dataIn1 = 32'd451
; 
32'd17748: dataIn1 = 32'd471
; 
32'd17749: dataIn1 = 32'd488
; 
32'd17750: dataIn1 = 32'd490
; 
32'd17751: dataIn1 = 32'd508
; 
32'd17752: dataIn1 = 32'd524
; 
32'd17753: dataIn1 = 32'd572
; 
32'd17754: dataIn1 = 32'd582
; 
32'd17755: dataIn1 = 32'd599
; 
32'd17756: dataIn1 = 32'd612
; 
32'd17757: dataIn1 = 32'd624
; 
32'd17758: dataIn1 = 32'd639
; 
32'd17759: dataIn1 = 32'd642
; 
32'd17760: dataIn1 = 32'd649
; 
32'd17761: dataIn1 = 32'd659
; 
32'd17762: dataIn1 = 32'd681
; 
32'd17763: dataIn1 = 32'd765
; 
32'd17764: dataIn1 = 32'd787
; 
32'd17765: dataIn1 = 32'd793
; 
32'd17766: dataIn1 = 32'd794
; 
32'd17767: dataIn1 = 32'd246
; 
32'd17768: dataIn1 = 32'd265
; 
32'd17769: dataIn1 = 32'd280
; 
32'd17770: dataIn1 = 32'd306
; 
32'd17771: dataIn1 = 32'd314
; 
32'd17772: dataIn1 = 32'd380
; 
32'd17773: dataIn1 = 32'd407
; 
32'd17774: dataIn1 = 32'd432
; 
32'd17775: dataIn1 = 32'd445
; 
32'd17776: dataIn1 = 32'd453
; 
32'd17777: dataIn1 = 32'd523
; 
32'd17778: dataIn1 = 32'd535
; 
32'd17779: dataIn1 = 32'd539
; 
32'd17780: dataIn1 = 32'd540
; 
32'd17781: dataIn1 = 32'd564
; 
32'd17782: dataIn1 = 32'd569
; 
32'd17783: dataIn1 = 32'd570
; 
32'd17784: dataIn1 = 32'd577
; 
32'd17785: dataIn1 = 32'd584
; 
32'd17786: dataIn1 = 32'd592
; 
32'd17787: dataIn1 = 32'd599
; 
32'd17788: dataIn1 = 32'd622
; 
32'd17789: dataIn1 = 32'd630
; 
32'd17790: dataIn1 = 32'd665
; 
32'd17791: dataIn1 = 32'd677
; 
32'd17792: dataIn1 = 32'd728
; 
32'd17793: dataIn1 = 32'd738
; 
32'd17794: dataIn1 = 32'd742
; 
32'd17795: dataIn1 = 32'd746
; 
32'd17796: dataIn1 = 32'd755
; 
32'd17797: dataIn1 = 32'd762
; 
32'd17798: dataIn1 = 32'd791
; 
32'd17799: dataIn1 = 32'd800
; 
32'd17800: dataIn1 = 32'd263
; 
32'd17801: dataIn1 = 32'd276
; 
32'd17802: dataIn1 = 32'd313
; 
32'd17803: dataIn1 = 32'd322
; 
32'd17804: dataIn1 = 32'd339
; 
32'd17805: dataIn1 = 32'd341
; 
32'd17806: dataIn1 = 32'd355
; 
32'd17807: dataIn1 = 32'd369
; 
32'd17808: dataIn1 = 32'd375
; 
32'd17809: dataIn1 = 32'd389
; 
32'd17810: dataIn1 = 32'd429
; 
32'd17811: dataIn1 = 32'd443
; 
32'd17812: dataIn1 = 32'd455
; 
32'd17813: dataIn1 = 32'd463
; 
32'd17814: dataIn1 = 32'd495
; 
32'd17815: dataIn1 = 32'd503
; 
32'd17816: dataIn1 = 32'd505
; 
32'd17817: dataIn1 = 32'd525
; 
32'd17818: dataIn1 = 32'd532
; 
32'd17819: dataIn1 = 32'd536
; 
32'd17820: dataIn1 = 32'd537
; 
32'd17821: dataIn1 = 32'd540
; 
32'd17822: dataIn1 = 32'd588
; 
32'd17823: dataIn1 = 32'd598
; 
32'd17824: dataIn1 = 32'd602
; 
32'd17825: dataIn1 = 32'd623
; 
32'd17826: dataIn1 = 32'd624
; 
32'd17827: dataIn1 = 32'd627
; 
32'd17828: dataIn1 = 32'd641
; 
32'd17829: dataIn1 = 32'd645
; 
32'd17830: dataIn1 = 32'd648
; 
32'd17831: dataIn1 = 32'd658
; 
32'd17832: dataIn1 = 32'd676
; 
32'd17833: dataIn1 = 32'd678
; 
32'd17834: dataIn1 = 32'd686
; 
32'd17835: dataIn1 = 32'd708
; 
32'd17836: dataIn1 = 32'd709
; 
32'd17837: dataIn1 = 32'd726
; 
32'd17838: dataIn1 = 32'd738
; 
32'd17839: dataIn1 = 32'd793
; 
32'd17840: dataIn1 = 32'd253
; 
32'd17841: dataIn1 = 32'd258
; 
32'd17842: dataIn1 = 32'd271
; 
32'd17843: dataIn1 = 32'd318
; 
32'd17844: dataIn1 = 32'd324
; 
32'd17845: dataIn1 = 32'd338
; 
32'd17846: dataIn1 = 32'd370
; 
32'd17847: dataIn1 = 32'd373
; 
32'd17848: dataIn1 = 32'd403
; 
32'd17849: dataIn1 = 32'd404
; 
32'd17850: dataIn1 = 32'd414
; 
32'd17851: dataIn1 = 32'd420
; 
32'd17852: dataIn1 = 32'd468
; 
32'd17853: dataIn1 = 32'd477
; 
32'd17854: dataIn1 = 32'd481
; 
32'd17855: dataIn1 = 32'd491
; 
32'd17856: dataIn1 = 32'd501
; 
32'd17857: dataIn1 = 32'd504
; 
32'd17858: dataIn1 = 32'd539
; 
32'd17859: dataIn1 = 32'd542
; 
32'd17860: dataIn1 = 32'd543
; 
32'd17861: dataIn1 = 32'd550
; 
32'd17862: dataIn1 = 32'd561
; 
32'd17863: dataIn1 = 32'd563
; 
32'd17864: dataIn1 = 32'd568
; 
32'd17865: dataIn1 = 32'd571
; 
32'd17866: dataIn1 = 32'd601
; 
32'd17867: dataIn1 = 32'd605
; 
32'd17868: dataIn1 = 32'd621
; 
32'd17869: dataIn1 = 32'd664
; 
32'd17870: dataIn1 = 32'd677
; 
32'd17871: dataIn1 = 32'd697
; 
32'd17872: dataIn1 = 32'd699
; 
32'd17873: dataIn1 = 32'd703
; 
32'd17874: dataIn1 = 32'd725
; 
32'd17875: dataIn1 = 32'd755
; 
32'd17876: dataIn1 = 32'd757
; 
32'd17877: dataIn1 = 32'd759
; 
32'd17878: dataIn1 = 32'd773
; 
32'd17879: dataIn1 = 32'd775
; 
32'd17880: dataIn1 = 32'd246
; 
32'd17881: dataIn1 = 32'd253
; 
32'd17882: dataIn1 = 32'd279
; 
32'd17883: dataIn1 = 32'd322
; 
32'd17884: dataIn1 = 32'd326
; 
32'd17885: dataIn1 = 32'd358
; 
32'd17886: dataIn1 = 32'd371
; 
32'd17887: dataIn1 = 32'd392
; 
32'd17888: dataIn1 = 32'd420
; 
32'd17889: dataIn1 = 32'd422
; 
32'd17890: dataIn1 = 32'd437
; 
32'd17891: dataIn1 = 32'd477
; 
32'd17892: dataIn1 = 32'd496
; 
32'd17893: dataIn1 = 32'd517
; 
32'd17894: dataIn1 = 32'd519
; 
32'd17895: dataIn1 = 32'd559
; 
32'd17896: dataIn1 = 32'd586
; 
32'd17897: dataIn1 = 32'd587
; 
32'd17898: dataIn1 = 32'd592
; 
32'd17899: dataIn1 = 32'd611
; 
32'd17900: dataIn1 = 32'd624
; 
32'd17901: dataIn1 = 32'd633
; 
32'd17902: dataIn1 = 32'd652
; 
32'd17903: dataIn1 = 32'd657
; 
32'd17904: dataIn1 = 32'd662
; 
32'd17905: dataIn1 = 32'd699
; 
32'd17906: dataIn1 = 32'd715
; 
32'd17907: dataIn1 = 32'd721
; 
32'd17908: dataIn1 = 32'd738
; 
32'd17909: dataIn1 = 32'd765
; 
32'd17910: dataIn1 = 32'd783
; 
32'd17911: dataIn1 = 32'd285
; 
32'd17912: dataIn1 = 32'd299
; 
32'd17913: dataIn1 = 32'd304
; 
32'd17914: dataIn1 = 32'd328
; 
32'd17915: dataIn1 = 32'd346
; 
32'd17916: dataIn1 = 32'd375
; 
32'd17917: dataIn1 = 32'd378
; 
32'd17918: dataIn1 = 32'd390
; 
32'd17919: dataIn1 = 32'd401
; 
32'd17920: dataIn1 = 32'd403
; 
32'd17921: dataIn1 = 32'd405
; 
32'd17922: dataIn1 = 32'd408
; 
32'd17923: dataIn1 = 32'd409
; 
32'd17924: dataIn1 = 32'd423
; 
32'd17925: dataIn1 = 32'd448
; 
32'd17926: dataIn1 = 32'd449
; 
32'd17927: dataIn1 = 32'd478
; 
32'd17928: dataIn1 = 32'd495
; 
32'd17929: dataIn1 = 32'd507
; 
32'd17930: dataIn1 = 32'd522
; 
32'd17931: dataIn1 = 32'd538
; 
32'd17932: dataIn1 = 32'd540
; 
32'd17933: dataIn1 = 32'd563
; 
32'd17934: dataIn1 = 32'd588
; 
32'd17935: dataIn1 = 32'd597
; 
32'd17936: dataIn1 = 32'd607
; 
32'd17937: dataIn1 = 32'd629
; 
32'd17938: dataIn1 = 32'd633
; 
32'd17939: dataIn1 = 32'd645
; 
32'd17940: dataIn1 = 32'd657
; 
32'd17941: dataIn1 = 32'd660
; 
32'd17942: dataIn1 = 32'd687
; 
32'd17943: dataIn1 = 32'd716
; 
32'd17944: dataIn1 = 32'd726
; 
32'd17945: dataIn1 = 32'd740
; 
32'd17946: dataIn1 = 32'd745
; 
32'd17947: dataIn1 = 32'd752
; 
32'd17948: dataIn1 = 32'd785
; 
32'd17949: dataIn1 = 32'd790
; 
32'd17950: dataIn1 = 32'd792
; 
32'd17951: dataIn1 = 32'd262
; 
32'd17952: dataIn1 = 32'd287
; 
32'd17953: dataIn1 = 32'd307
; 
32'd17954: dataIn1 = 32'd342
; 
32'd17955: dataIn1 = 32'd346
; 
32'd17956: dataIn1 = 32'd355
; 
32'd17957: dataIn1 = 32'd357
; 
32'd17958: dataIn1 = 32'd376
; 
32'd17959: dataIn1 = 32'd406
; 
32'd17960: dataIn1 = 32'd433
; 
32'd17961: dataIn1 = 32'd469
; 
32'd17962: dataIn1 = 32'd474
; 
32'd17963: dataIn1 = 32'd502
; 
32'd17964: dataIn1 = 32'd530
; 
32'd17965: dataIn1 = 32'd536
; 
32'd17966: dataIn1 = 32'd552
; 
32'd17967: dataIn1 = 32'd556
; 
32'd17968: dataIn1 = 32'd559
; 
32'd17969: dataIn1 = 32'd562
; 
32'd17970: dataIn1 = 32'd582
; 
32'd17971: dataIn1 = 32'd590
; 
32'd17972: dataIn1 = 32'd599
; 
32'd17973: dataIn1 = 32'd666
; 
32'd17974: dataIn1 = 32'd699
; 
32'd17975: dataIn1 = 32'd710
; 
32'd17976: dataIn1 = 32'd723
; 
32'd17977: dataIn1 = 32'd743
; 
32'd17978: dataIn1 = 32'd754
; 
32'd17979: dataIn1 = 32'd760
; 
32'd17980: dataIn1 = 32'd779
; 
32'd17981: dataIn1 = 32'd785
; 
32'd17982: dataIn1 = 32'd786
; 
32'd17983: dataIn1 = 32'd790
; 
32'd17984: dataIn1 = 32'd278
; 
32'd17985: dataIn1 = 32'd284
; 
32'd17986: dataIn1 = 32'd302
; 
32'd17987: dataIn1 = 32'd314
; 
32'd17988: dataIn1 = 32'd322
; 
32'd17989: dataIn1 = 32'd347
; 
32'd17990: dataIn1 = 32'd350
; 
32'd17991: dataIn1 = 32'd381
; 
32'd17992: dataIn1 = 32'd414
; 
32'd17993: dataIn1 = 32'd417
; 
32'd17994: dataIn1 = 32'd466
; 
32'd17995: dataIn1 = 32'd490
; 
32'd17996: dataIn1 = 32'd491
; 
32'd17997: dataIn1 = 32'd497
; 
32'd17998: dataIn1 = 32'd516
; 
32'd17999: dataIn1 = 32'd547
; 
32'd18000: dataIn1 = 32'd549
; 
32'd18001: dataIn1 = 32'd587
; 
32'd18002: dataIn1 = 32'd592
; 
32'd18003: dataIn1 = 32'd647
; 
32'd18004: dataIn1 = 32'd658
; 
32'd18005: dataIn1 = 32'd662
; 
32'd18006: dataIn1 = 32'd665
; 
32'd18007: dataIn1 = 32'd668
; 
32'd18008: dataIn1 = 32'd680
; 
32'd18009: dataIn1 = 32'd701
; 
32'd18010: dataIn1 = 32'd703
; 
32'd18011: dataIn1 = 32'd706
; 
32'd18012: dataIn1 = 32'd712
; 
32'd18013: dataIn1 = 32'd748
; 
32'd18014: dataIn1 = 32'd783
; 
32'd18015: dataIn1 = 32'd794
; 
32'd18016: dataIn1 = 32'd799
; 
32'd18017: dataIn1 = 32'd800
; 
32'd18018: dataIn1 = 32'd253
; 
32'd18019: dataIn1 = 32'd269
; 
32'd18020: dataIn1 = 32'd271
; 
32'd18021: dataIn1 = 32'd288
; 
32'd18022: dataIn1 = 32'd309
; 
32'd18023: dataIn1 = 32'd316
; 
32'd18024: dataIn1 = 32'd318
; 
32'd18025: dataIn1 = 32'd333
; 
32'd18026: dataIn1 = 32'd348
; 
32'd18027: dataIn1 = 32'd362
; 
32'd18028: dataIn1 = 32'd366
; 
32'd18029: dataIn1 = 32'd387
; 
32'd18030: dataIn1 = 32'd436
; 
32'd18031: dataIn1 = 32'd438
; 
32'd18032: dataIn1 = 32'd457
; 
32'd18033: dataIn1 = 32'd510
; 
32'd18034: dataIn1 = 32'd537
; 
32'd18035: dataIn1 = 32'd566
; 
32'd18036: dataIn1 = 32'd582
; 
32'd18037: dataIn1 = 32'd585
; 
32'd18038: dataIn1 = 32'd647
; 
32'd18039: dataIn1 = 32'd675
; 
32'd18040: dataIn1 = 32'd686
; 
32'd18041: dataIn1 = 32'd687
; 
32'd18042: dataIn1 = 32'd690
; 
32'd18043: dataIn1 = 32'd694
; 
32'd18044: dataIn1 = 32'd695
; 
32'd18045: dataIn1 = 32'd704
; 
32'd18046: dataIn1 = 32'd732
; 
32'd18047: dataIn1 = 32'd745
; 
32'd18048: dataIn1 = 32'd747
; 
32'd18049: dataIn1 = 32'd752
; 
32'd18050: dataIn1 = 32'd763
; 
32'd18051: dataIn1 = 32'd788
; 
32'd18052: dataIn1 = 32'd790
; 
32'd18053: dataIn1 = 32'd285
; 
32'd18054: dataIn1 = 32'd307
; 
32'd18055: dataIn1 = 32'd314
; 
32'd18056: dataIn1 = 32'd336
; 
32'd18057: dataIn1 = 32'd348
; 
32'd18058: dataIn1 = 32'd350
; 
32'd18059: dataIn1 = 32'd358
; 
32'd18060: dataIn1 = 32'd360
; 
32'd18061: dataIn1 = 32'd364
; 
32'd18062: dataIn1 = 32'd369
; 
32'd18063: dataIn1 = 32'd434
; 
32'd18064: dataIn1 = 32'd453
; 
32'd18065: dataIn1 = 32'd454
; 
32'd18066: dataIn1 = 32'd465
; 
32'd18067: dataIn1 = 32'd485
; 
32'd18068: dataIn1 = 32'd495
; 
32'd18069: dataIn1 = 32'd516
; 
32'd18070: dataIn1 = 32'd517
; 
32'd18071: dataIn1 = 32'd535
; 
32'd18072: dataIn1 = 32'd540
; 
32'd18073: dataIn1 = 32'd547
; 
32'd18074: dataIn1 = 32'd560
; 
32'd18075: dataIn1 = 32'd574
; 
32'd18076: dataIn1 = 32'd579
; 
32'd18077: dataIn1 = 32'd627
; 
32'd18078: dataIn1 = 32'd634
; 
32'd18079: dataIn1 = 32'd638
; 
32'd18080: dataIn1 = 32'd684
; 
32'd18081: dataIn1 = 32'd702
; 
32'd18082: dataIn1 = 32'd736
; 
32'd18083: dataIn1 = 32'd756
; 
32'd18084: dataIn1 = 32'd764
; 
32'd18085: dataIn1 = 32'd784
; 
32'd18086: dataIn1 = 32'd789
; 
32'd18087: dataIn1 = 32'd263
; 
32'd18088: dataIn1 = 32'd265
; 
32'd18089: dataIn1 = 32'd283
; 
32'd18090: dataIn1 = 32'd285
; 
32'd18091: dataIn1 = 32'd305
; 
32'd18092: dataIn1 = 32'd394
; 
32'd18093: dataIn1 = 32'd405
; 
32'd18094: dataIn1 = 32'd421
; 
32'd18095: dataIn1 = 32'd430
; 
32'd18096: dataIn1 = 32'd468
; 
32'd18097: dataIn1 = 32'd512
; 
32'd18098: dataIn1 = 32'd540
; 
32'd18099: dataIn1 = 32'd543
; 
32'd18100: dataIn1 = 32'd548
; 
32'd18101: dataIn1 = 32'd587
; 
32'd18102: dataIn1 = 32'd599
; 
32'd18103: dataIn1 = 32'd621
; 
32'd18104: dataIn1 = 32'd623
; 
32'd18105: dataIn1 = 32'd631
; 
32'd18106: dataIn1 = 32'd638
; 
32'd18107: dataIn1 = 32'd650
; 
32'd18108: dataIn1 = 32'd652
; 
32'd18109: dataIn1 = 32'd663
; 
32'd18110: dataIn1 = 32'd674
; 
32'd18111: dataIn1 = 32'd685
; 
32'd18112: dataIn1 = 32'd697
; 
32'd18113: dataIn1 = 32'd699
; 
32'd18114: dataIn1 = 32'd714
; 
32'd18115: dataIn1 = 32'd727
; 
32'd18116: dataIn1 = 32'd728
; 
32'd18117: dataIn1 = 32'd732
; 
32'd18118: dataIn1 = 32'd754
; 
32'd18119: dataIn1 = 32'd762
; 
32'd18120: dataIn1 = 32'd767
; 
32'd18121: dataIn1 = 32'd780
; 
32'd18122: dataIn1 = 32'd290
; 
32'd18123: dataIn1 = 32'd297
; 
32'd18124: dataIn1 = 32'd303
; 
32'd18125: dataIn1 = 32'd343
; 
32'd18126: dataIn1 = 32'd363
; 
32'd18127: dataIn1 = 32'd374
; 
32'd18128: dataIn1 = 32'd386
; 
32'd18129: dataIn1 = 32'd399
; 
32'd18130: dataIn1 = 32'd402
; 
32'd18131: dataIn1 = 32'd440
; 
32'd18132: dataIn1 = 32'd453
; 
32'd18133: dataIn1 = 32'd474
; 
32'd18134: dataIn1 = 32'd505
; 
32'd18135: dataIn1 = 32'd508
; 
32'd18136: dataIn1 = 32'd537
; 
32'd18137: dataIn1 = 32'd551
; 
32'd18138: dataIn1 = 32'd571
; 
32'd18139: dataIn1 = 32'd603
; 
32'd18140: dataIn1 = 32'd604
; 
32'd18141: dataIn1 = 32'd609
; 
32'd18142: dataIn1 = 32'd621
; 
32'd18143: dataIn1 = 32'd630
; 
32'd18144: dataIn1 = 32'd663
; 
32'd18145: dataIn1 = 32'd666
; 
32'd18146: dataIn1 = 32'd676
; 
32'd18147: dataIn1 = 32'd694
; 
32'd18148: dataIn1 = 32'd716
; 
32'd18149: dataIn1 = 32'd720
; 
32'd18150: dataIn1 = 32'd725
; 
32'd18151: dataIn1 = 32'd739
; 
32'd18152: dataIn1 = 32'd745
; 
32'd18153: dataIn1 = 32'd758
; 
32'd18154: dataIn1 = 32'd781
; 
32'd18155: dataIn1 = 32'd791
; 
32'd18156: dataIn1 = 32'd798
; 
32'd18157: dataIn1 = 32'd266
; 
32'd18158: dataIn1 = 32'd270
; 
32'd18159: dataIn1 = 32'd281
; 
32'd18160: dataIn1 = 32'd293
; 
32'd18161: dataIn1 = 32'd311
; 
32'd18162: dataIn1 = 32'd312
; 
32'd18163: dataIn1 = 32'd313
; 
32'd18164: dataIn1 = 32'd330
; 
32'd18165: dataIn1 = 32'd334
; 
32'd18166: dataIn1 = 32'd354
; 
32'd18167: dataIn1 = 32'd382
; 
32'd18168: dataIn1 = 32'd385
; 
32'd18169: dataIn1 = 32'd389
; 
32'd18170: dataIn1 = 32'd426
; 
32'd18171: dataIn1 = 32'd433
; 
32'd18172: dataIn1 = 32'd444
; 
32'd18173: dataIn1 = 32'd452
; 
32'd18174: dataIn1 = 32'd455
; 
32'd18175: dataIn1 = 32'd464
; 
32'd18176: dataIn1 = 32'd477
; 
32'd18177: dataIn1 = 32'd489
; 
32'd18178: dataIn1 = 32'd509
; 
32'd18179: dataIn1 = 32'd519
; 
32'd18180: dataIn1 = 32'd525
; 
32'd18181: dataIn1 = 32'd527
; 
32'd18182: dataIn1 = 32'd531
; 
32'd18183: dataIn1 = 32'd546
; 
32'd18184: dataIn1 = 32'd561
; 
32'd18185: dataIn1 = 32'd567
; 
32'd18186: dataIn1 = 32'd580
; 
32'd18187: dataIn1 = 32'd589
; 
32'd18188: dataIn1 = 32'd596
; 
32'd18189: dataIn1 = 32'd597
; 
32'd18190: dataIn1 = 32'd611
; 
32'd18191: dataIn1 = 32'd619
; 
32'd18192: dataIn1 = 32'd642
; 
32'd18193: dataIn1 = 32'd665
; 
32'd18194: dataIn1 = 32'd704
; 
32'd18195: dataIn1 = 32'd714
; 
32'd18196: dataIn1 = 32'd725
; 
32'd18197: dataIn1 = 32'd735
; 
32'd18198: dataIn1 = 32'd739
; 
32'd18199: dataIn1 = 32'd750
; 
32'd18200: dataIn1 = 32'd752
; 
32'd18201: dataIn1 = 32'd753
; 
32'd18202: dataIn1 = 32'd758
; 
32'd18203: dataIn1 = 32'd763
; 
32'd18204: dataIn1 = 32'd777
; 
32'd18205: dataIn1 = 32'd780
; 
32'd18206: dataIn1 = 32'd283
; 
32'd18207: dataIn1 = 32'd296
; 
32'd18208: dataIn1 = 32'd327
; 
32'd18209: dataIn1 = 32'd332
; 
32'd18210: dataIn1 = 32'd349
; 
32'd18211: dataIn1 = 32'd364
; 
32'd18212: dataIn1 = 32'd396
; 
32'd18213: dataIn1 = 32'd419
; 
32'd18214: dataIn1 = 32'd426
; 
32'd18215: dataIn1 = 32'd429
; 
32'd18216: dataIn1 = 32'd438
; 
32'd18217: dataIn1 = 32'd482
; 
32'd18218: dataIn1 = 32'd484
; 
32'd18219: dataIn1 = 32'd491
; 
32'd18220: dataIn1 = 32'd508
; 
32'd18221: dataIn1 = 32'd521
; 
32'd18222: dataIn1 = 32'd540
; 
32'd18223: dataIn1 = 32'd548
; 
32'd18224: dataIn1 = 32'd587
; 
32'd18225: dataIn1 = 32'd604
; 
32'd18226: dataIn1 = 32'd618
; 
32'd18227: dataIn1 = 32'd628
; 
32'd18228: dataIn1 = 32'd672
; 
32'd18229: dataIn1 = 32'd681
; 
32'd18230: dataIn1 = 32'd709
; 
32'd18231: dataIn1 = 32'd726
; 
32'd18232: dataIn1 = 32'd732
; 
32'd18233: dataIn1 = 32'd741
; 
32'd18234: dataIn1 = 32'd755
; 
32'd18235: dataIn1 = 32'd781
; 
32'd18236: dataIn1 = 32'd263
; 
32'd18237: dataIn1 = 32'd284
; 
32'd18238: dataIn1 = 32'd310
; 
32'd18239: dataIn1 = 32'd321
; 
32'd18240: dataIn1 = 32'd325
; 
32'd18241: dataIn1 = 32'd330
; 
32'd18242: dataIn1 = 32'd333
; 
32'd18243: dataIn1 = 32'd344
; 
32'd18244: dataIn1 = 32'd353
; 
32'd18245: dataIn1 = 32'd375
; 
32'd18246: dataIn1 = 32'd382
; 
32'd18247: dataIn1 = 32'd393
; 
32'd18248: dataIn1 = 32'd424
; 
32'd18249: dataIn1 = 32'd455
; 
32'd18250: dataIn1 = 32'd462
; 
32'd18251: dataIn1 = 32'd470
; 
32'd18252: dataIn1 = 32'd478
; 
32'd18253: dataIn1 = 32'd490
; 
32'd18254: dataIn1 = 32'd506
; 
32'd18255: dataIn1 = 32'd516
; 
32'd18256: dataIn1 = 32'd522
; 
32'd18257: dataIn1 = 32'd526
; 
32'd18258: dataIn1 = 32'd541
; 
32'd18259: dataIn1 = 32'd546
; 
32'd18260: dataIn1 = 32'd548
; 
32'd18261: dataIn1 = 32'd554
; 
32'd18262: dataIn1 = 32'd557
; 
32'd18263: dataIn1 = 32'd572
; 
32'd18264: dataIn1 = 32'd573
; 
32'd18265: dataIn1 = 32'd599
; 
32'd18266: dataIn1 = 32'd639
; 
32'd18267: dataIn1 = 32'd644
; 
32'd18268: dataIn1 = 32'd647
; 
32'd18269: dataIn1 = 32'd655
; 
32'd18270: dataIn1 = 32'd661
; 
32'd18271: dataIn1 = 32'd665
; 
32'd18272: dataIn1 = 32'd672
; 
32'd18273: dataIn1 = 32'd685
; 
32'd18274: dataIn1 = 32'd736
; 
32'd18275: dataIn1 = 32'd786
; 
32'd18276: dataIn1 = 32'd799
; 
32'd18277: dataIn1 = 32'd276
; 
32'd18278: dataIn1 = 32'd283
; 
32'd18279: dataIn1 = 32'd293
; 
32'd18280: dataIn1 = 32'd304
; 
32'd18281: dataIn1 = 32'd309
; 
32'd18282: dataIn1 = 32'd324
; 
32'd18283: dataIn1 = 32'd329
; 
32'd18284: dataIn1 = 32'd341
; 
32'd18285: dataIn1 = 32'd346
; 
32'd18286: dataIn1 = 32'd367
; 
32'd18287: dataIn1 = 32'd462
; 
32'd18288: dataIn1 = 32'd485
; 
32'd18289: dataIn1 = 32'd552
; 
32'd18290: dataIn1 = 32'd583
; 
32'd18291: dataIn1 = 32'd587
; 
32'd18292: dataIn1 = 32'd608
; 
32'd18293: dataIn1 = 32'd630
; 
32'd18294: dataIn1 = 32'd639
; 
32'd18295: dataIn1 = 32'd649
; 
32'd18296: dataIn1 = 32'd650
; 
32'd18297: dataIn1 = 32'd657
; 
32'd18298: dataIn1 = 32'd675
; 
32'd18299: dataIn1 = 32'd678
; 
32'd18300: dataIn1 = 32'd703
; 
32'd18301: dataIn1 = 32'd704
; 
32'd18302: dataIn1 = 32'd708
; 
32'd18303: dataIn1 = 32'd709
; 
32'd18304: dataIn1 = 32'd719
; 
32'd18305: dataIn1 = 32'd721
; 
32'd18306: dataIn1 = 32'd722
; 
32'd18307: dataIn1 = 32'd723
; 
32'd18308: dataIn1 = 32'd725
; 
32'd18309: dataIn1 = 32'd760
; 
32'd18310: dataIn1 = 32'd762
; 
32'd18311: dataIn1 = 32'd770
; 
32'd18312: dataIn1 = 32'd776
; 
32'd18313: dataIn1 = 32'd796
; 
32'd18314: dataIn1 = 32'd800
; 
32'd18315: dataIn1 = 32'd273
; 
32'd18316: dataIn1 = 32'd291
; 
32'd18317: dataIn1 = 32'd295
; 
32'd18318: dataIn1 = 32'd297
; 
32'd18319: dataIn1 = 32'd332
; 
32'd18320: dataIn1 = 32'd345
; 
32'd18321: dataIn1 = 32'd369
; 
32'd18322: dataIn1 = 32'd404
; 
32'd18323: dataIn1 = 32'd422
; 
32'd18324: dataIn1 = 32'd426
; 
32'd18325: dataIn1 = 32'd441
; 
32'd18326: dataIn1 = 32'd471
; 
32'd18327: dataIn1 = 32'd486
; 
32'd18328: dataIn1 = 32'd489
; 
32'd18329: dataIn1 = 32'd519
; 
32'd18330: dataIn1 = 32'd525
; 
32'd18331: dataIn1 = 32'd552
; 
32'd18332: dataIn1 = 32'd558
; 
32'd18333: dataIn1 = 32'd559
; 
32'd18334: dataIn1 = 32'd560
; 
32'd18335: dataIn1 = 32'd564
; 
32'd18336: dataIn1 = 32'd566
; 
32'd18337: dataIn1 = 32'd578
; 
32'd18338: dataIn1 = 32'd601
; 
32'd18339: dataIn1 = 32'd602
; 
32'd18340: dataIn1 = 32'd603
; 
32'd18341: dataIn1 = 32'd606
; 
32'd18342: dataIn1 = 32'd616
; 
32'd18343: dataIn1 = 32'd617
; 
32'd18344: dataIn1 = 32'd639
; 
32'd18345: dataIn1 = 32'd673
; 
32'd18346: dataIn1 = 32'd693
; 
32'd18347: dataIn1 = 32'd701
; 
32'd18348: dataIn1 = 32'd702
; 
32'd18349: dataIn1 = 32'd704
; 
32'd18350: dataIn1 = 32'd713
; 
32'd18351: dataIn1 = 32'd747
; 
32'd18352: dataIn1 = 32'd752
; 
32'd18353: dataIn1 = 32'd753
; 
32'd18354: dataIn1 = 32'd770
; 
32'd18355: dataIn1 = 32'd771
; 
32'd18356: dataIn1 = 32'd774
; 
32'd18357: dataIn1 = 32'd797
; 
32'd18358: dataIn1 = 32'd798
; 
32'd18359: dataIn1 = 32'd262
; 
32'd18360: dataIn1 = 32'd269
; 
32'd18361: dataIn1 = 32'd274
; 
32'd18362: dataIn1 = 32'd284
; 
32'd18363: dataIn1 = 32'd295
; 
32'd18364: dataIn1 = 32'd298
; 
32'd18365: dataIn1 = 32'd300
; 
32'd18366: dataIn1 = 32'd301
; 
32'd18367: dataIn1 = 32'd309
; 
32'd18368: dataIn1 = 32'd321
; 
32'd18369: dataIn1 = 32'd325
; 
32'd18370: dataIn1 = 32'd328
; 
32'd18371: dataIn1 = 32'd341
; 
32'd18372: dataIn1 = 32'd345
; 
32'd18373: dataIn1 = 32'd366
; 
32'd18374: dataIn1 = 32'd385
; 
32'd18375: dataIn1 = 32'd400
; 
32'd18376: dataIn1 = 32'd402
; 
32'd18377: dataIn1 = 32'd413
; 
32'd18378: dataIn1 = 32'd423
; 
32'd18379: dataIn1 = 32'd463
; 
32'd18380: dataIn1 = 32'd466
; 
32'd18381: dataIn1 = 32'd476
; 
32'd18382: dataIn1 = 32'd507
; 
32'd18383: dataIn1 = 32'd531
; 
32'd18384: dataIn1 = 32'd563
; 
32'd18385: dataIn1 = 32'd570
; 
32'd18386: dataIn1 = 32'd624
; 
32'd18387: dataIn1 = 32'd625
; 
32'd18388: dataIn1 = 32'd663
; 
32'd18389: dataIn1 = 32'd671
; 
32'd18390: dataIn1 = 32'd688
; 
32'd18391: dataIn1 = 32'd696
; 
32'd18392: dataIn1 = 32'd698
; 
32'd18393: dataIn1 = 32'd713
; 
32'd18394: dataIn1 = 32'd734
; 
32'd18395: dataIn1 = 32'd737
; 
32'd18396: dataIn1 = 32'd748
; 
32'd18397: dataIn1 = 32'd770
; 
32'd18398: dataIn1 = 32'd778
; 
32'd18399: dataIn1 = 32'd783
; 
32'd18400: dataIn1 = 32'd273
; 
32'd18401: dataIn1 = 32'd279
; 
32'd18402: dataIn1 = 32'd309
; 
32'd18403: dataIn1 = 32'd319
; 
32'd18404: dataIn1 = 32'd360
; 
32'd18405: dataIn1 = 32'd361
; 
32'd18406: dataIn1 = 32'd402
; 
32'd18407: dataIn1 = 32'd405
; 
32'd18408: dataIn1 = 32'd439
; 
32'd18409: dataIn1 = 32'd453
; 
32'd18410: dataIn1 = 32'd457
; 
32'd18411: dataIn1 = 32'd469
; 
32'd18412: dataIn1 = 32'd473
; 
32'd18413: dataIn1 = 32'd476
; 
32'd18414: dataIn1 = 32'd482
; 
32'd18415: dataIn1 = 32'd489
; 
32'd18416: dataIn1 = 32'd502
; 
32'd18417: dataIn1 = 32'd505
; 
32'd18418: dataIn1 = 32'd538
; 
32'd18419: dataIn1 = 32'd554
; 
32'd18420: dataIn1 = 32'd570
; 
32'd18421: dataIn1 = 32'd577
; 
32'd18422: dataIn1 = 32'd600
; 
32'd18423: dataIn1 = 32'd635
; 
32'd18424: dataIn1 = 32'd643
; 
32'd18425: dataIn1 = 32'd662
; 
32'd18426: dataIn1 = 32'd695
; 
32'd18427: dataIn1 = 32'd707
; 
32'd18428: dataIn1 = 32'd719
; 
32'd18429: dataIn1 = 32'd723
; 
32'd18430: dataIn1 = 32'd774
; 
32'd18431: dataIn1 = 32'd798
; 
32'd18432: dataIn1 = 32'd285
; 
32'd18433: dataIn1 = 32'd288
; 
32'd18434: dataIn1 = 32'd308
; 
32'd18435: dataIn1 = 32'd310
; 
32'd18436: dataIn1 = 32'd312
; 
32'd18437: dataIn1 = 32'd335
; 
32'd18438: dataIn1 = 32'd339
; 
32'd18439: dataIn1 = 32'd340
; 
32'd18440: dataIn1 = 32'd341
; 
32'd18441: dataIn1 = 32'd346
; 
32'd18442: dataIn1 = 32'd363
; 
32'd18443: dataIn1 = 32'd365
; 
32'd18444: dataIn1 = 32'd379
; 
32'd18445: dataIn1 = 32'd399
; 
32'd18446: dataIn1 = 32'd418
; 
32'd18447: dataIn1 = 32'd426
; 
32'd18448: dataIn1 = 32'd462
; 
32'd18449: dataIn1 = 32'd465
; 
32'd18450: dataIn1 = 32'd476
; 
32'd18451: dataIn1 = 32'd477
; 
32'd18452: dataIn1 = 32'd483
; 
32'd18453: dataIn1 = 32'd486
; 
32'd18454: dataIn1 = 32'd497
; 
32'd18455: dataIn1 = 32'd516
; 
32'd18456: dataIn1 = 32'd572
; 
32'd18457: dataIn1 = 32'd589
; 
32'd18458: dataIn1 = 32'd602
; 
32'd18459: dataIn1 = 32'd617
; 
32'd18460: dataIn1 = 32'd627
; 
32'd18461: dataIn1 = 32'd642
; 
32'd18462: dataIn1 = 32'd654
; 
32'd18463: dataIn1 = 32'd672
; 
32'd18464: dataIn1 = 32'd726
; 
32'd18465: dataIn1 = 32'd759
; 
32'd18466: dataIn1 = 32'd776
; 
32'd18467: dataIn1 = 32'd791
; 
32'd18468: dataIn1 = 32'd792
; 
32'd18469: dataIn1 = 32'd800
; 
32'd18470: dataIn1 = 32'd262
; 
32'd18471: dataIn1 = 32'd269
; 
32'd18472: dataIn1 = 32'd290
; 
32'd18473: dataIn1 = 32'd297
; 
32'd18474: dataIn1 = 32'd298
; 
32'd18475: dataIn1 = 32'd309
; 
32'd18476: dataIn1 = 32'd310
; 
32'd18477: dataIn1 = 32'd327
; 
32'd18478: dataIn1 = 32'd346
; 
32'd18479: dataIn1 = 32'd356
; 
32'd18480: dataIn1 = 32'd359
; 
32'd18481: dataIn1 = 32'd362
; 
32'd18482: dataIn1 = 32'd365
; 
32'd18483: dataIn1 = 32'd370
; 
32'd18484: dataIn1 = 32'd375
; 
32'd18485: dataIn1 = 32'd388
; 
32'd18486: dataIn1 = 32'd426
; 
32'd18487: dataIn1 = 32'd427
; 
32'd18488: dataIn1 = 32'd430
; 
32'd18489: dataIn1 = 32'd435
; 
32'd18490: dataIn1 = 32'd442
; 
32'd18491: dataIn1 = 32'd446
; 
32'd18492: dataIn1 = 32'd459
; 
32'd18493: dataIn1 = 32'd464
; 
32'd18494: dataIn1 = 32'd472
; 
32'd18495: dataIn1 = 32'd479
; 
32'd18496: dataIn1 = 32'd481
; 
32'd18497: dataIn1 = 32'd495
; 
32'd18498: dataIn1 = 32'd504
; 
32'd18499: dataIn1 = 32'd513
; 
32'd18500: dataIn1 = 32'd626
; 
32'd18501: dataIn1 = 32'd655
; 
32'd18502: dataIn1 = 32'd705
; 
32'd18503: dataIn1 = 32'd717
; 
32'd18504: dataIn1 = 32'd730
; 
32'd18505: dataIn1 = 32'd738
; 
32'd18506: dataIn1 = 32'd746
; 
32'd18507: dataIn1 = 32'd753
; 
32'd18508: dataIn1 = 32'd762
; 
32'd18509: dataIn1 = 32'd272
; 
32'd18510: dataIn1 = 32'd289
; 
32'd18511: dataIn1 = 32'd357
; 
32'd18512: dataIn1 = 32'd366
; 
32'd18513: dataIn1 = 32'd421
; 
32'd18514: dataIn1 = 32'd435
; 
32'd18515: dataIn1 = 32'd455
; 
32'd18516: dataIn1 = 32'd469
; 
32'd18517: dataIn1 = 32'd472
; 
32'd18518: dataIn1 = 32'd479
; 
32'd18519: dataIn1 = 32'd505
; 
32'd18520: dataIn1 = 32'd567
; 
32'd18521: dataIn1 = 32'd587
; 
32'd18522: dataIn1 = 32'd626
; 
32'd18523: dataIn1 = 32'd635
; 
32'd18524: dataIn1 = 32'd648
; 
32'd18525: dataIn1 = 32'd681
; 
32'd18526: dataIn1 = 32'd684
; 
32'd18527: dataIn1 = 32'd710
; 
32'd18528: dataIn1 = 32'd736
; 
32'd18529: dataIn1 = 32'd738
; 
32'd18530: dataIn1 = 32'd751
; 
32'd18531: dataIn1 = 32'd761
; 
32'd18532: dataIn1 = 32'd782
; 
32'd18533: dataIn1 = 32'd789
; 
32'd18534: dataIn1 = 32'd283
; 
32'd18535: dataIn1 = 32'd297
; 
32'd18536: dataIn1 = 32'd304
; 
32'd18537: dataIn1 = 32'd314
; 
32'd18538: dataIn1 = 32'd316
; 
32'd18539: dataIn1 = 32'd359
; 
32'd18540: dataIn1 = 32'd378
; 
32'd18541: dataIn1 = 32'd394
; 
32'd18542: dataIn1 = 32'd408
; 
32'd18543: dataIn1 = 32'd466
; 
32'd18544: dataIn1 = 32'd480
; 
32'd18545: dataIn1 = 32'd482
; 
32'd18546: dataIn1 = 32'd484
; 
32'd18547: dataIn1 = 32'd509
; 
32'd18548: dataIn1 = 32'd514
; 
32'd18549: dataIn1 = 32'd517
; 
32'd18550: dataIn1 = 32'd519
; 
32'd18551: dataIn1 = 32'd521
; 
32'd18552: dataIn1 = 32'd537
; 
32'd18553: dataIn1 = 32'd555
; 
32'd18554: dataIn1 = 32'd569
; 
32'd18555: dataIn1 = 32'd617
; 
32'd18556: dataIn1 = 32'd642
; 
32'd18557: dataIn1 = 32'd644
; 
32'd18558: dataIn1 = 32'd658
; 
32'd18559: dataIn1 = 32'd696
; 
32'd18560: dataIn1 = 32'd708
; 
32'd18561: dataIn1 = 32'd729
; 
32'd18562: dataIn1 = 32'd736
; 
32'd18563: dataIn1 = 32'd757
; 
32'd18564: dataIn1 = 32'd772
; 
32'd18565: dataIn1 = 32'd780
; 
32'd18566: dataIn1 = 32'd787
; 
32'd18567: dataIn1 = 32'd275
; 
32'd18568: dataIn1 = 32'd291
; 
32'd18569: dataIn1 = 32'd293
; 
32'd18570: dataIn1 = 32'd296
; 
32'd18571: dataIn1 = 32'd334
; 
32'd18572: dataIn1 = 32'd362
; 
32'd18573: dataIn1 = 32'd372
; 
32'd18574: dataIn1 = 32'd386
; 
32'd18575: dataIn1 = 32'd388
; 
32'd18576: dataIn1 = 32'd423
; 
32'd18577: dataIn1 = 32'd447
; 
32'd18578: dataIn1 = 32'd450
; 
32'd18579: dataIn1 = 32'd497
; 
32'd18580: dataIn1 = 32'd506
; 
32'd18581: dataIn1 = 32'd517
; 
32'd18582: dataIn1 = 32'd545
; 
32'd18583: dataIn1 = 32'd560
; 
32'd18584: dataIn1 = 32'd563
; 
32'd18585: dataIn1 = 32'd567
; 
32'd18586: dataIn1 = 32'd570
; 
32'd18587: dataIn1 = 32'd580
; 
32'd18588: dataIn1 = 32'd582
; 
32'd18589: dataIn1 = 32'd583
; 
32'd18590: dataIn1 = 32'd589
; 
32'd18591: dataIn1 = 32'd605
; 
32'd18592: dataIn1 = 32'd606
; 
32'd18593: dataIn1 = 32'd625
; 
32'd18594: dataIn1 = 32'd627
; 
32'd18595: dataIn1 = 32'd663
; 
32'd18596: dataIn1 = 32'd667
; 
32'd18597: dataIn1 = 32'd675
; 
32'd18598: dataIn1 = 32'd681
; 
32'd18599: dataIn1 = 32'd695
; 
32'd18600: dataIn1 = 32'd717
; 
32'd18601: dataIn1 = 32'd723
; 
32'd18602: dataIn1 = 32'd736
; 
32'd18603: dataIn1 = 32'd751
; 
32'd18604: dataIn1 = 32'd753
; 
32'd18605: dataIn1 = 32'd757
; 
32'd18606: dataIn1 = 32'd759
; 
32'd18607: dataIn1 = 32'd778
; 
32'd18608: dataIn1 = 32'd783
; 
32'd18609: dataIn1 = 32'd793
; 
32'd18610: dataIn1 = 32'd268
; 
32'd18611: dataIn1 = 32'd279
; 
32'd18612: dataIn1 = 32'd283
; 
32'd18613: dataIn1 = 32'd295
; 
32'd18614: dataIn1 = 32'd306
; 
32'd18615: dataIn1 = 32'd307
; 
32'd18616: dataIn1 = 32'd319
; 
32'd18617: dataIn1 = 32'd327
; 
32'd18618: dataIn1 = 32'd354
; 
32'd18619: dataIn1 = 32'd357
; 
32'd18620: dataIn1 = 32'd382
; 
32'd18621: dataIn1 = 32'd389
; 
32'd18622: dataIn1 = 32'd428
; 
32'd18623: dataIn1 = 32'd478
; 
32'd18624: dataIn1 = 32'd497
; 
32'd18625: dataIn1 = 32'd498
; 
32'd18626: dataIn1 = 32'd509
; 
32'd18627: dataIn1 = 32'd523
; 
32'd18628: dataIn1 = 32'd557
; 
32'd18629: dataIn1 = 32'd564
; 
32'd18630: dataIn1 = 32'd573
; 
32'd18631: dataIn1 = 32'd575
; 
32'd18632: dataIn1 = 32'd593
; 
32'd18633: dataIn1 = 32'd603
; 
32'd18634: dataIn1 = 32'd617
; 
32'd18635: dataIn1 = 32'd620
; 
32'd18636: dataIn1 = 32'd622
; 
32'd18637: dataIn1 = 32'd635
; 
32'd18638: dataIn1 = 32'd639
; 
32'd18639: dataIn1 = 32'd655
; 
32'd18640: dataIn1 = 32'd664
; 
32'd18641: dataIn1 = 32'd705
; 
32'd18642: dataIn1 = 32'd712
; 
32'd18643: dataIn1 = 32'd733
; 
32'd18644: dataIn1 = 32'd746
; 
32'd18645: dataIn1 = 32'd747
; 
32'd18646: dataIn1 = 32'd761
; 
32'd18647: dataIn1 = 32'd795
; 
32'd18648: dataIn1 = 32'd266
; 
32'd18649: dataIn1 = 32'd286
; 
32'd18650: dataIn1 = 32'd319
; 
32'd18651: dataIn1 = 32'd330
; 
32'd18652: dataIn1 = 32'd332
; 
32'd18653: dataIn1 = 32'd379
; 
32'd18654: dataIn1 = 32'd400
; 
32'd18655: dataIn1 = 32'd439
; 
32'd18656: dataIn1 = 32'd440
; 
32'd18657: dataIn1 = 32'd442
; 
32'd18658: dataIn1 = 32'd470
; 
32'd18659: dataIn1 = 32'd480
; 
32'd18660: dataIn1 = 32'd483
; 
32'd18661: dataIn1 = 32'd498
; 
32'd18662: dataIn1 = 32'd518
; 
32'd18663: dataIn1 = 32'd519
; 
32'd18664: dataIn1 = 32'd535
; 
32'd18665: dataIn1 = 32'd548
; 
32'd18666: dataIn1 = 32'd550
; 
32'd18667: dataIn1 = 32'd557
; 
32'd18668: dataIn1 = 32'd558
; 
32'd18669: dataIn1 = 32'd578
; 
32'd18670: dataIn1 = 32'd610
; 
32'd18671: dataIn1 = 32'd626
; 
32'd18672: dataIn1 = 32'd643
; 
32'd18673: dataIn1 = 32'd680
; 
32'd18674: dataIn1 = 32'd684
; 
32'd18675: dataIn1 = 32'd717
; 
32'd18676: dataIn1 = 32'd738
; 
32'd18677: dataIn1 = 32'd742
; 
32'd18678: dataIn1 = 32'd760
; 
32'd18679: dataIn1 = 32'd768
; 
32'd18680: dataIn1 = 32'd770
; 
32'd18681: dataIn1 = 32'd771
; 
32'd18682: dataIn1 = 32'd786
; 
32'd18683: dataIn1 = 32'd367
; 
32'd18684: dataIn1 = 32'd371
; 
32'd18685: dataIn1 = 32'd373
; 
32'd18686: dataIn1 = 32'd424
; 
32'd18687: dataIn1 = 32'd482
; 
32'd18688: dataIn1 = 32'd513
; 
32'd18689: dataIn1 = 32'd531
; 
32'd18690: dataIn1 = 32'd577
; 
32'd18691: dataIn1 = 32'd590
; 
32'd18692: dataIn1 = 32'd603
; 
32'd18693: dataIn1 = 32'd608
; 
32'd18694: dataIn1 = 32'd623
; 
32'd18695: dataIn1 = 32'd634
; 
32'd18696: dataIn1 = 32'd635
; 
32'd18697: dataIn1 = 32'd674
; 
32'd18698: dataIn1 = 32'd678
; 
32'd18699: dataIn1 = 32'd682
; 
32'd18700: dataIn1 = 32'd696
; 
32'd18701: dataIn1 = 32'd712
; 
32'd18702: dataIn1 = 32'd731
; 
32'd18703: dataIn1 = 32'd744
; 
32'd18704: dataIn1 = 32'd759
; 
32'd18705: dataIn1 = 32'd769
; 
32'd18706: dataIn1 = 32'd790
; 
32'd18707: dataIn1 = 32'd792
; 
32'd18708: dataIn1 = 32'd272
; 
32'd18709: dataIn1 = 32'd279
; 
32'd18710: dataIn1 = 32'd291
; 
32'd18711: dataIn1 = 32'd313
; 
32'd18712: dataIn1 = 32'd325
; 
32'd18713: dataIn1 = 32'd331
; 
32'd18714: dataIn1 = 32'd338
; 
32'd18715: dataIn1 = 32'd430
; 
32'd18716: dataIn1 = 32'd448
; 
32'd18717: dataIn1 = 32'd471
; 
32'd18718: dataIn1 = 32'd483
; 
32'd18719: dataIn1 = 32'd498
; 
32'd18720: dataIn1 = 32'd504
; 
32'd18721: dataIn1 = 32'd514
; 
32'd18722: dataIn1 = 32'd516
; 
32'd18723: dataIn1 = 32'd519
; 
32'd18724: dataIn1 = 32'd523
; 
32'd18725: dataIn1 = 32'd602
; 
32'd18726: dataIn1 = 32'd618
; 
32'd18727: dataIn1 = 32'd621
; 
32'd18728: dataIn1 = 32'd622
; 
32'd18729: dataIn1 = 32'd627
; 
32'd18730: dataIn1 = 32'd641
; 
32'd18731: dataIn1 = 32'd644
; 
32'd18732: dataIn1 = 32'd654
; 
32'd18733: dataIn1 = 32'd659
; 
32'd18734: dataIn1 = 32'd672
; 
32'd18735: dataIn1 = 32'd683
; 
32'd18736: dataIn1 = 32'd688
; 
32'd18737: dataIn1 = 32'd708
; 
32'd18738: dataIn1 = 32'd732
; 
32'd18739: dataIn1 = 32'd756
; 
32'd18740: dataIn1 = 32'd786
; 
32'd18741: dataIn1 = 32'd794
; 
32'd18742: dataIn1 = 32'd269
; 
32'd18743: dataIn1 = 32'd291
; 
32'd18744: dataIn1 = 32'd295
; 
32'd18745: dataIn1 = 32'd322
; 
32'd18746: dataIn1 = 32'd323
; 
32'd18747: dataIn1 = 32'd367
; 
32'd18748: dataIn1 = 32'd376
; 
32'd18749: dataIn1 = 32'd400
; 
32'd18750: dataIn1 = 32'd432
; 
32'd18751: dataIn1 = 32'd433
; 
32'd18752: dataIn1 = 32'd446
; 
32'd18753: dataIn1 = 32'd453
; 
32'd18754: dataIn1 = 32'd471
; 
32'd18755: dataIn1 = 32'd499
; 
32'd18756: dataIn1 = 32'd511
; 
32'd18757: dataIn1 = 32'd524
; 
32'd18758: dataIn1 = 32'd576
; 
32'd18759: dataIn1 = 32'd595
; 
32'd18760: dataIn1 = 32'd600
; 
32'd18761: dataIn1 = 32'd601
; 
32'd18762: dataIn1 = 32'd643
; 
32'd18763: dataIn1 = 32'd649
; 
32'd18764: dataIn1 = 32'd661
; 
32'd18765: dataIn1 = 32'd683
; 
32'd18766: dataIn1 = 32'd687
; 
32'd18767: dataIn1 = 32'd743
; 
32'd18768: dataIn1 = 32'd747
; 
32'd18769: dataIn1 = 32'd755
; 
32'd18770: dataIn1 = 32'd761
; 
32'd18771: dataIn1 = 32'd765
; 
32'd18772: dataIn1 = 32'd769
; 
32'd18773: dataIn1 = 32'd795
; 
32'd18774: dataIn1 = 32'd797
; 
32'd18775: dataIn1 = 32'd799
; 
32'd18776: dataIn1 = 32'd326
; 
32'd18777: dataIn1 = 32'd342
; 
32'd18778: dataIn1 = 32'd350
; 
32'd18779: dataIn1 = 32'd356
; 
32'd18780: dataIn1 = 32'd359
; 
32'd18781: dataIn1 = 32'd362
; 
32'd18782: dataIn1 = 32'd372
; 
32'd18783: dataIn1 = 32'd383
; 
32'd18784: dataIn1 = 32'd406
; 
32'd18785: dataIn1 = 32'd441
; 
32'd18786: dataIn1 = 32'd477
; 
32'd18787: dataIn1 = 32'd490
; 
32'd18788: dataIn1 = 32'd539
; 
32'd18789: dataIn1 = 32'd586
; 
32'd18790: dataIn1 = 32'd623
; 
32'd18791: dataIn1 = 32'd631
; 
32'd18792: dataIn1 = 32'd632
; 
32'd18793: dataIn1 = 32'd668
; 
32'd18794: dataIn1 = 32'd673
; 
32'd18795: dataIn1 = 32'd722
; 
32'd18796: dataIn1 = 32'd725
; 
32'd18797: dataIn1 = 32'd754
; 
32'd18798: dataIn1 = 32'd762
; 
32'd18799: dataIn1 = 32'd764
; 
32'd18800: dataIn1 = 32'd778
; 
32'd18801: dataIn1 = 32'd279
; 
32'd18802: dataIn1 = 32'd283
; 
32'd18803: dataIn1 = 32'd289
; 
32'd18804: dataIn1 = 32'd292
; 
32'd18805: dataIn1 = 32'd294
; 
32'd18806: dataIn1 = 32'd303
; 
32'd18807: dataIn1 = 32'd305
; 
32'd18808: dataIn1 = 32'd333
; 
32'd18809: dataIn1 = 32'd342
; 
32'd18810: dataIn1 = 32'd346
; 
32'd18811: dataIn1 = 32'd367
; 
32'd18812: dataIn1 = 32'd376
; 
32'd18813: dataIn1 = 32'd409
; 
32'd18814: dataIn1 = 32'd434
; 
32'd18815: dataIn1 = 32'd475
; 
32'd18816: dataIn1 = 32'd491
; 
32'd18817: dataIn1 = 32'd493
; 
32'd18818: dataIn1 = 32'd496
; 
32'd18819: dataIn1 = 32'd520
; 
32'd18820: dataIn1 = 32'd529
; 
32'd18821: dataIn1 = 32'd558
; 
32'd18822: dataIn1 = 32'd580
; 
32'd18823: dataIn1 = 32'd610
; 
32'd18824: dataIn1 = 32'd638
; 
32'd18825: dataIn1 = 32'd659
; 
32'd18826: dataIn1 = 32'd669
; 
32'd18827: dataIn1 = 32'd675
; 
32'd18828: dataIn1 = 32'd685
; 
32'd18829: dataIn1 = 32'd706
; 
32'd18830: dataIn1 = 32'd712
; 
32'd18831: dataIn1 = 32'd745
; 
32'd18832: dataIn1 = 32'd768
; 
32'd18833: dataIn1 = 32'd778
; 
32'd18834: dataIn1 = 32'd280
; 
32'd18835: dataIn1 = 32'd287
; 
32'd18836: dataIn1 = 32'd335
; 
32'd18837: dataIn1 = 32'd336
; 
32'd18838: dataIn1 = 32'd337
; 
32'd18839: dataIn1 = 32'd346
; 
32'd18840: dataIn1 = 32'd370
; 
32'd18841: dataIn1 = 32'd374
; 
32'd18842: dataIn1 = 32'd382
; 
32'd18843: dataIn1 = 32'd396
; 
32'd18844: dataIn1 = 32'd420
; 
32'd18845: dataIn1 = 32'd424
; 
32'd18846: dataIn1 = 32'd425
; 
32'd18847: dataIn1 = 32'd432
; 
32'd18848: dataIn1 = 32'd455
; 
32'd18849: dataIn1 = 32'd460
; 
32'd18850: dataIn1 = 32'd468
; 
32'd18851: dataIn1 = 32'd473
; 
32'd18852: dataIn1 = 32'd488
; 
32'd18853: dataIn1 = 32'd489
; 
32'd18854: dataIn1 = 32'd532
; 
32'd18855: dataIn1 = 32'd542
; 
32'd18856: dataIn1 = 32'd551
; 
32'd18857: dataIn1 = 32'd559
; 
32'd18858: dataIn1 = 32'd577
; 
32'd18859: dataIn1 = 32'd585
; 
32'd18860: dataIn1 = 32'd636
; 
32'd18861: dataIn1 = 32'd690
; 
32'd18862: dataIn1 = 32'd695
; 
32'd18863: dataIn1 = 32'd716
; 
32'd18864: dataIn1 = 32'd717
; 
32'd18865: dataIn1 = 32'd730
; 
32'd18866: dataIn1 = 32'd740
; 
32'd18867: dataIn1 = 32'd746
; 
32'd18868: dataIn1 = 32'd767
; 
32'd18869: dataIn1 = 32'd768
; 
32'd18870: dataIn1 = 32'd789
; 
32'd18871: dataIn1 = 32'd284
; 
32'd18872: dataIn1 = 32'd285
; 
32'd18873: dataIn1 = 32'd296
; 
32'd18874: dataIn1 = 32'd332
; 
32'd18875: dataIn1 = 32'd356
; 
32'd18876: dataIn1 = 32'd361
; 
32'd18877: dataIn1 = 32'd393
; 
32'd18878: dataIn1 = 32'd395
; 
32'd18879: dataIn1 = 32'd447
; 
32'd18880: dataIn1 = 32'd455
; 
32'd18881: dataIn1 = 32'd460
; 
32'd18882: dataIn1 = 32'd463
; 
32'd18883: dataIn1 = 32'd476
; 
32'd18884: dataIn1 = 32'd483
; 
32'd18885: dataIn1 = 32'd491
; 
32'd18886: dataIn1 = 32'd495
; 
32'd18887: dataIn1 = 32'd498
; 
32'd18888: dataIn1 = 32'd522
; 
32'd18889: dataIn1 = 32'd523
; 
32'd18890: dataIn1 = 32'd533
; 
32'd18891: dataIn1 = 32'd535
; 
32'd18892: dataIn1 = 32'd565
; 
32'd18893: dataIn1 = 32'd572
; 
32'd18894: dataIn1 = 32'd608
; 
32'd18895: dataIn1 = 32'd651
; 
32'd18896: dataIn1 = 32'd654
; 
32'd18897: dataIn1 = 32'd658
; 
32'd18898: dataIn1 = 32'd663
; 
32'd18899: dataIn1 = 32'd674
; 
32'd18900: dataIn1 = 32'd691
; 
32'd18901: dataIn1 = 32'd699
; 
32'd18902: dataIn1 = 32'd713
; 
32'd18903: dataIn1 = 32'd748
; 
32'd18904: dataIn1 = 32'd749
; 
32'd18905: dataIn1 = 32'd788
; 
32'd18906: dataIn1 = 32'd798
; 
32'd18907: dataIn1 = 32'd290
; 
32'd18908: dataIn1 = 32'd318
; 
32'd18909: dataIn1 = 32'd327
; 
32'd18910: dataIn1 = 32'd333
; 
32'd18911: dataIn1 = 32'd344
; 
32'd18912: dataIn1 = 32'd355
; 
32'd18913: dataIn1 = 32'd382
; 
32'd18914: dataIn1 = 32'd393
; 
32'd18915: dataIn1 = 32'd402
; 
32'd18916: dataIn1 = 32'd410
; 
32'd18917: dataIn1 = 32'd415
; 
32'd18918: dataIn1 = 32'd424
; 
32'd18919: dataIn1 = 32'd457
; 
32'd18920: dataIn1 = 32'd516
; 
32'd18921: dataIn1 = 32'd548
; 
32'd18922: dataIn1 = 32'd553
; 
32'd18923: dataIn1 = 32'd582
; 
32'd18924: dataIn1 = 32'd588
; 
32'd18925: dataIn1 = 32'd592
; 
32'd18926: dataIn1 = 32'd603
; 
32'd18927: dataIn1 = 32'd614
; 
32'd18928: dataIn1 = 32'd616
; 
32'd18929: dataIn1 = 32'd632
; 
32'd18930: dataIn1 = 32'd643
; 
32'd18931: dataIn1 = 32'd661
; 
32'd18932: dataIn1 = 32'd665
; 
32'd18933: dataIn1 = 32'd666
; 
32'd18934: dataIn1 = 32'd689
; 
32'd18935: dataIn1 = 32'd691
; 
32'd18936: dataIn1 = 32'd694
; 
32'd18937: dataIn1 = 32'd697
; 
32'd18938: dataIn1 = 32'd701
; 
32'd18939: dataIn1 = 32'd737
; 
32'd18940: dataIn1 = 32'd747
; 
32'd18941: dataIn1 = 32'd749
; 
32'd18942: dataIn1 = 32'd773
; 
32'd18943: dataIn1 = 32'd796
; 
32'd18944: dataIn1 = 32'd296
; 
32'd18945: dataIn1 = 32'd321
; 
32'd18946: dataIn1 = 32'd336
; 
32'd18947: dataIn1 = 32'd338
; 
32'd18948: dataIn1 = 32'd343
; 
32'd18949: dataIn1 = 32'd389
; 
32'd18950: dataIn1 = 32'd396
; 
32'd18951: dataIn1 = 32'd435
; 
32'd18952: dataIn1 = 32'd437
; 
32'd18953: dataIn1 = 32'd444
; 
32'd18954: dataIn1 = 32'd445
; 
32'd18955: dataIn1 = 32'd460
; 
32'd18956: dataIn1 = 32'd470
; 
32'd18957: dataIn1 = 32'd502
; 
32'd18958: dataIn1 = 32'd535
; 
32'd18959: dataIn1 = 32'd548
; 
32'd18960: dataIn1 = 32'd560
; 
32'd18961: dataIn1 = 32'd590
; 
32'd18962: dataIn1 = 32'd592
; 
32'd18963: dataIn1 = 32'd602
; 
32'd18964: dataIn1 = 32'd613
; 
32'd18965: dataIn1 = 32'd669
; 
32'd18966: dataIn1 = 32'd704
; 
32'd18967: dataIn1 = 32'd705
; 
32'd18968: dataIn1 = 32'd714
; 
32'd18969: dataIn1 = 32'd720
; 
32'd18970: dataIn1 = 32'd732
; 
32'd18971: dataIn1 = 32'd752
; 
32'd18972: dataIn1 = 32'd769
; 
32'd18973: dataIn1 = 32'd781
; 
32'd18974: dataIn1 = 32'd786
; 
32'd18975: dataIn1 = 32'd792
; 
32'd18976: dataIn1 = 32'd286
; 
32'd18977: dataIn1 = 32'd289
; 
32'd18978: dataIn1 = 32'd290
; 
32'd18979: dataIn1 = 32'd300
; 
32'd18980: dataIn1 = 32'd304
; 
32'd18981: dataIn1 = 32'd322
; 
32'd18982: dataIn1 = 32'd366
; 
32'd18983: dataIn1 = 32'd384
; 
32'd18984: dataIn1 = 32'd387
; 
32'd18985: dataIn1 = 32'd388
; 
32'd18986: dataIn1 = 32'd390
; 
32'd18987: dataIn1 = 32'd398
; 
32'd18988: dataIn1 = 32'd404
; 
32'd18989: dataIn1 = 32'd407
; 
32'd18990: dataIn1 = 32'd437
; 
32'd18991: dataIn1 = 32'd494
; 
32'd18992: dataIn1 = 32'd496
; 
32'd18993: dataIn1 = 32'd515
; 
32'd18994: dataIn1 = 32'd535
; 
32'd18995: dataIn1 = 32'd536
; 
32'd18996: dataIn1 = 32'd561
; 
32'd18997: dataIn1 = 32'd591
; 
32'd18998: dataIn1 = 32'd609
; 
32'd18999: dataIn1 = 32'd620
; 
32'd19000: dataIn1 = 32'd656
; 
32'd19001: dataIn1 = 32'd664
; 
32'd19002: dataIn1 = 32'd666
; 
32'd19003: dataIn1 = 32'd683
; 
32'd19004: dataIn1 = 32'd720
; 
32'd19005: dataIn1 = 32'd722
; 
32'd19006: dataIn1 = 32'd733
; 
32'd19007: dataIn1 = 32'd737
; 
32'd19008: dataIn1 = 32'd743
; 
32'd19009: dataIn1 = 32'd778
; 
32'd19010: dataIn1 = 32'd792
; 
32'd19011: dataIn1 = 32'd795
; 
32'd19012: dataIn1 = 32'd797
; 
32'd19013: dataIn1 = 32'd284
; 
32'd19014: dataIn1 = 32'd287
; 
32'd19015: dataIn1 = 32'd293
; 
32'd19016: dataIn1 = 32'd300
; 
32'd19017: dataIn1 = 32'd304
; 
32'd19018: dataIn1 = 32'd323
; 
32'd19019: dataIn1 = 32'd340
; 
32'd19020: dataIn1 = 32'd342
; 
32'd19021: dataIn1 = 32'd348
; 
32'd19022: dataIn1 = 32'd383
; 
32'd19023: dataIn1 = 32'd409
; 
32'd19024: dataIn1 = 32'd410
; 
32'd19025: dataIn1 = 32'd419
; 
32'd19026: dataIn1 = 32'd423
; 
32'd19027: dataIn1 = 32'd445
; 
32'd19028: dataIn1 = 32'd459
; 
32'd19029: dataIn1 = 32'd482
; 
32'd19030: dataIn1 = 32'd491
; 
32'd19031: dataIn1 = 32'd525
; 
32'd19032: dataIn1 = 32'd552
; 
32'd19033: dataIn1 = 32'd560
; 
32'd19034: dataIn1 = 32'd576
; 
32'd19035: dataIn1 = 32'd628
; 
32'd19036: dataIn1 = 32'd649
; 
32'd19037: dataIn1 = 32'd650
; 
32'd19038: dataIn1 = 32'd651
; 
32'd19039: dataIn1 = 32'd671
; 
32'd19040: dataIn1 = 32'd707
; 
32'd19041: dataIn1 = 32'd723
; 
32'd19042: dataIn1 = 32'd730
; 
32'd19043: dataIn1 = 32'd741
; 
32'd19044: dataIn1 = 32'd749
; 
32'd19045: dataIn1 = 32'd779
; 
32'd19046: dataIn1 = 32'd797
; 
32'd19047: dataIn1 = 32'd278
; 
32'd19048: dataIn1 = 32'd284
; 
32'd19049: dataIn1 = 32'd286
; 
32'd19050: dataIn1 = 32'd292
; 
32'd19051: dataIn1 = 32'd295
; 
32'd19052: dataIn1 = 32'd307
; 
32'd19053: dataIn1 = 32'd308
; 
32'd19054: dataIn1 = 32'd310
; 
32'd19055: dataIn1 = 32'd315
; 
32'd19056: dataIn1 = 32'd336
; 
32'd19057: dataIn1 = 32'd375
; 
32'd19058: dataIn1 = 32'd380
; 
32'd19059: dataIn1 = 32'd388
; 
32'd19060: dataIn1 = 32'd391
; 
32'd19061: dataIn1 = 32'd402
; 
32'd19062: dataIn1 = 32'd410
; 
32'd19063: dataIn1 = 32'd413
; 
32'd19064: dataIn1 = 32'd435
; 
32'd19065: dataIn1 = 32'd448
; 
32'd19066: dataIn1 = 32'd450
; 
32'd19067: dataIn1 = 32'd454
; 
32'd19068: dataIn1 = 32'd464
; 
32'd19069: dataIn1 = 32'd495
; 
32'd19070: dataIn1 = 32'd522
; 
32'd19071: dataIn1 = 32'd543
; 
32'd19072: dataIn1 = 32'd544
; 
32'd19073: dataIn1 = 32'd546
; 
32'd19074: dataIn1 = 32'd549
; 
32'd19075: dataIn1 = 32'd576
; 
32'd19076: dataIn1 = 32'd577
; 
32'd19077: dataIn1 = 32'd636
; 
32'd19078: dataIn1 = 32'd671
; 
32'd19079: dataIn1 = 32'd690
; 
32'd19080: dataIn1 = 32'd717
; 
32'd19081: dataIn1 = 32'd720
; 
32'd19082: dataIn1 = 32'd725
; 
32'd19083: dataIn1 = 32'd746
; 
32'd19084: dataIn1 = 32'd753
; 
32'd19085: dataIn1 = 32'd760
; 
32'd19086: dataIn1 = 32'd764
; 
32'd19087: dataIn1 = 32'd791
; 
32'd19088: dataIn1 = 32'd793
; 
32'd19089: dataIn1 = 32'd798
; 
32'd19090: dataIn1 = 32'd279
; 
32'd19091: dataIn1 = 32'd293
; 
32'd19092: dataIn1 = 32'd295
; 
32'd19093: dataIn1 = 32'd296
; 
32'd19094: dataIn1 = 32'd308
; 
32'd19095: dataIn1 = 32'd318
; 
32'd19096: dataIn1 = 32'd321
; 
32'd19097: dataIn1 = 32'd340
; 
32'd19098: dataIn1 = 32'd361
; 
32'd19099: dataIn1 = 32'd370
; 
32'd19100: dataIn1 = 32'd383
; 
32'd19101: dataIn1 = 32'd398
; 
32'd19102: dataIn1 = 32'd408
; 
32'd19103: dataIn1 = 32'd411
; 
32'd19104: dataIn1 = 32'd420
; 
32'd19105: dataIn1 = 32'd437
; 
32'd19106: dataIn1 = 32'd467
; 
32'd19107: dataIn1 = 32'd471
; 
32'd19108: dataIn1 = 32'd489
; 
32'd19109: dataIn1 = 32'd518
; 
32'd19110: dataIn1 = 32'd533
; 
32'd19111: dataIn1 = 32'd536
; 
32'd19112: dataIn1 = 32'd537
; 
32'd19113: dataIn1 = 32'd565
; 
32'd19114: dataIn1 = 32'd585
; 
32'd19115: dataIn1 = 32'd606
; 
32'd19116: dataIn1 = 32'd614
; 
32'd19117: dataIn1 = 32'd669
; 
32'd19118: dataIn1 = 32'd682
; 
32'd19119: dataIn1 = 32'd687
; 
32'd19120: dataIn1 = 32'd714
; 
32'd19121: dataIn1 = 32'd736
; 
32'd19122: dataIn1 = 32'd738
; 
32'd19123: dataIn1 = 32'd748
; 
32'd19124: dataIn1 = 32'd753
; 
32'd19125: dataIn1 = 32'd779
; 
32'd19126: dataIn1 = 32'd285
; 
32'd19127: dataIn1 = 32'd302
; 
32'd19128: dataIn1 = 32'd307
; 
32'd19129: dataIn1 = 32'd308
; 
32'd19130: dataIn1 = 32'd311
; 
32'd19131: dataIn1 = 32'd316
; 
32'd19132: dataIn1 = 32'd340
; 
32'd19133: dataIn1 = 32'd347
; 
32'd19134: dataIn1 = 32'd353
; 
32'd19135: dataIn1 = 32'd354
; 
32'd19136: dataIn1 = 32'd363
; 
32'd19137: dataIn1 = 32'd366
; 
32'd19138: dataIn1 = 32'd374
; 
32'd19139: dataIn1 = 32'd376
; 
32'd19140: dataIn1 = 32'd402
; 
32'd19141: dataIn1 = 32'd448
; 
32'd19142: dataIn1 = 32'd490
; 
32'd19143: dataIn1 = 32'd504
; 
32'd19144: dataIn1 = 32'd522
; 
32'd19145: dataIn1 = 32'd584
; 
32'd19146: dataIn1 = 32'd595
; 
32'd19147: dataIn1 = 32'd618
; 
32'd19148: dataIn1 = 32'd644
; 
32'd19149: dataIn1 = 32'd649
; 
32'd19150: dataIn1 = 32'd653
; 
32'd19151: dataIn1 = 32'd674
; 
32'd19152: dataIn1 = 32'd679
; 
32'd19153: dataIn1 = 32'd684
; 
32'd19154: dataIn1 = 32'd685
; 
32'd19155: dataIn1 = 32'd285
; 
32'd19156: dataIn1 = 32'd286
; 
32'd19157: dataIn1 = 32'd304
; 
32'd19158: dataIn1 = 32'd309
; 
32'd19159: dataIn1 = 32'd349
; 
32'd19160: dataIn1 = 32'd359
; 
32'd19161: dataIn1 = 32'd365
; 
32'd19162: dataIn1 = 32'd382
; 
32'd19163: dataIn1 = 32'd403
; 
32'd19164: dataIn1 = 32'd408
; 
32'd19165: dataIn1 = 32'd412
; 
32'd19166: dataIn1 = 32'd432
; 
32'd19167: dataIn1 = 32'd461
; 
32'd19168: dataIn1 = 32'd473
; 
32'd19169: dataIn1 = 32'd497
; 
32'd19170: dataIn1 = 32'd522
; 
32'd19171: dataIn1 = 32'd523
; 
32'd19172: dataIn1 = 32'd539
; 
32'd19173: dataIn1 = 32'd552
; 
32'd19174: dataIn1 = 32'd559
; 
32'd19175: dataIn1 = 32'd560
; 
32'd19176: dataIn1 = 32'd624
; 
32'd19177: dataIn1 = 32'd641
; 
32'd19178: dataIn1 = 32'd646
; 
32'd19179: dataIn1 = 32'd647
; 
32'd19180: dataIn1 = 32'd692
; 
32'd19181: dataIn1 = 32'd755
; 
32'd19182: dataIn1 = 32'd761
; 
32'd19183: dataIn1 = 32'd782
; 
32'd19184: dataIn1 = 32'd793
; 
32'd19185: dataIn1 = 32'd799
; 
32'd19186: dataIn1 = 32'd287
; 
32'd19187: dataIn1 = 32'd301
; 
32'd19188: dataIn1 = 32'd351
; 
32'd19189: dataIn1 = 32'd365
; 
32'd19190: dataIn1 = 32'd369
; 
32'd19191: dataIn1 = 32'd371
; 
32'd19192: dataIn1 = 32'd394
; 
32'd19193: dataIn1 = 32'd402
; 
32'd19194: dataIn1 = 32'd414
; 
32'd19195: dataIn1 = 32'd424
; 
32'd19196: dataIn1 = 32'd466
; 
32'd19197: dataIn1 = 32'd467
; 
32'd19198: dataIn1 = 32'd476
; 
32'd19199: dataIn1 = 32'd504
; 
32'd19200: dataIn1 = 32'd514
; 
32'd19201: dataIn1 = 32'd526
; 
32'd19202: dataIn1 = 32'd543
; 
32'd19203: dataIn1 = 32'd554
; 
32'd19204: dataIn1 = 32'd560
; 
32'd19205: dataIn1 = 32'd569
; 
32'd19206: dataIn1 = 32'd570
; 
32'd19207: dataIn1 = 32'd587
; 
32'd19208: dataIn1 = 32'd622
; 
32'd19209: dataIn1 = 32'd640
; 
32'd19210: dataIn1 = 32'd644
; 
32'd19211: dataIn1 = 32'd677
; 
32'd19212: dataIn1 = 32'd684
; 
32'd19213: dataIn1 = 32'd691
; 
32'd19214: dataIn1 = 32'd703
; 
32'd19215: dataIn1 = 32'd777
; 
32'd19216: dataIn1 = 32'd793
; 
32'd19217: dataIn1 = 32'd800
; 
32'd19218: dataIn1 = 32'd283
; 
32'd19219: dataIn1 = 32'd286
; 
32'd19220: dataIn1 = 32'd294
; 
32'd19221: dataIn1 = 32'd304
; 
32'd19222: dataIn1 = 32'd311
; 
32'd19223: dataIn1 = 32'd321
; 
32'd19224: dataIn1 = 32'd332
; 
32'd19225: dataIn1 = 32'd349
; 
32'd19226: dataIn1 = 32'd376
; 
32'd19227: dataIn1 = 32'd383
; 
32'd19228: dataIn1 = 32'd400
; 
32'd19229: dataIn1 = 32'd408
; 
32'd19230: dataIn1 = 32'd410
; 
32'd19231: dataIn1 = 32'd411
; 
32'd19232: dataIn1 = 32'd413
; 
32'd19233: dataIn1 = 32'd427
; 
32'd19234: dataIn1 = 32'd468
; 
32'd19235: dataIn1 = 32'd512
; 
32'd19236: dataIn1 = 32'd525
; 
32'd19237: dataIn1 = 32'd528
; 
32'd19238: dataIn1 = 32'd533
; 
32'd19239: dataIn1 = 32'd538
; 
32'd19240: dataIn1 = 32'd558
; 
32'd19241: dataIn1 = 32'd560
; 
32'd19242: dataIn1 = 32'd576
; 
32'd19243: dataIn1 = 32'd623
; 
32'd19244: dataIn1 = 32'd656
; 
32'd19245: dataIn1 = 32'd682
; 
32'd19246: dataIn1 = 32'd689
; 
32'd19247: dataIn1 = 32'd699
; 
32'd19248: dataIn1 = 32'd718
; 
32'd19249: dataIn1 = 32'd726
; 
32'd19250: dataIn1 = 32'd738
; 
32'd19251: dataIn1 = 32'd750
; 
32'd19252: dataIn1 = 32'd758
; 
32'd19253: dataIn1 = 32'd794
; 
32'd19254: dataIn1 = 32'd296
; 
32'd19255: dataIn1 = 32'd312
; 
32'd19256: dataIn1 = 32'd315
; 
32'd19257: dataIn1 = 32'd330
; 
32'd19258: dataIn1 = 32'd349
; 
32'd19259: dataIn1 = 32'd358
; 
32'd19260: dataIn1 = 32'd375
; 
32'd19261: dataIn1 = 32'd398
; 
32'd19262: dataIn1 = 32'd403
; 
32'd19263: dataIn1 = 32'd441
; 
32'd19264: dataIn1 = 32'd463
; 
32'd19265: dataIn1 = 32'd483
; 
32'd19266: dataIn1 = 32'd498
; 
32'd19267: dataIn1 = 32'd499
; 
32'd19268: dataIn1 = 32'd550
; 
32'd19269: dataIn1 = 32'd570
; 
32'd19270: dataIn1 = 32'd574
; 
32'd19271: dataIn1 = 32'd596
; 
32'd19272: dataIn1 = 32'd629
; 
32'd19273: dataIn1 = 32'd639
; 
32'd19274: dataIn1 = 32'd658
; 
32'd19275: dataIn1 = 32'd667
; 
32'd19276: dataIn1 = 32'd673
; 
32'd19277: dataIn1 = 32'd719
; 
32'd19278: dataIn1 = 32'd727
; 
32'd19279: dataIn1 = 32'd735
; 
32'd19280: dataIn1 = 32'd743
; 
32'd19281: dataIn1 = 32'd748
; 
32'd19282: dataIn1 = 32'd753
; 
32'd19283: dataIn1 = 32'd771
; 
32'd19284: dataIn1 = 32'd787
; 
32'd19285: dataIn1 = 32'd795
; 
32'd19286: dataIn1 = 32'd310
; 
32'd19287: dataIn1 = 32'd316
; 
32'd19288: dataIn1 = 32'd332
; 
32'd19289: dataIn1 = 32'd341
; 
32'd19290: dataIn1 = 32'd376
; 
32'd19291: dataIn1 = 32'd377
; 
32'd19292: dataIn1 = 32'd379
; 
32'd19293: dataIn1 = 32'd384
; 
32'd19294: dataIn1 = 32'd394
; 
32'd19295: dataIn1 = 32'd397
; 
32'd19296: dataIn1 = 32'd404
; 
32'd19297: dataIn1 = 32'd407
; 
32'd19298: dataIn1 = 32'd427
; 
32'd19299: dataIn1 = 32'd456
; 
32'd19300: dataIn1 = 32'd464
; 
32'd19301: dataIn1 = 32'd473
; 
32'd19302: dataIn1 = 32'd475
; 
32'd19303: dataIn1 = 32'd528
; 
32'd19304: dataIn1 = 32'd594
; 
32'd19305: dataIn1 = 32'd602
; 
32'd19306: dataIn1 = 32'd613
; 
32'd19307: dataIn1 = 32'd630
; 
32'd19308: dataIn1 = 32'd640
; 
32'd19309: dataIn1 = 32'd642
; 
32'd19310: dataIn1 = 32'd645
; 
32'd19311: dataIn1 = 32'd672
; 
32'd19312: dataIn1 = 32'd717
; 
32'd19313: dataIn1 = 32'd721
; 
32'd19314: dataIn1 = 32'd777
; 
32'd19315: dataIn1 = 32'd300
; 
32'd19316: dataIn1 = 32'd309
; 
32'd19317: dataIn1 = 32'd314
; 
32'd19318: dataIn1 = 32'd323
; 
32'd19319: dataIn1 = 32'd388
; 
32'd19320: dataIn1 = 32'd394
; 
32'd19321: dataIn1 = 32'd410
; 
32'd19322: dataIn1 = 32'd423
; 
32'd19323: dataIn1 = 32'd424
; 
32'd19324: dataIn1 = 32'd450
; 
32'd19325: dataIn1 = 32'd496
; 
32'd19326: dataIn1 = 32'd515
; 
32'd19327: dataIn1 = 32'd517
; 
32'd19328: dataIn1 = 32'd519
; 
32'd19329: dataIn1 = 32'd520
; 
32'd19330: dataIn1 = 32'd524
; 
32'd19331: dataIn1 = 32'd528
; 
32'd19332: dataIn1 = 32'd538
; 
32'd19333: dataIn1 = 32'd546
; 
32'd19334: dataIn1 = 32'd562
; 
32'd19335: dataIn1 = 32'd572
; 
32'd19336: dataIn1 = 32'd593
; 
32'd19337: dataIn1 = 32'd610
; 
32'd19338: dataIn1 = 32'd706
; 
32'd19339: dataIn1 = 32'd718
; 
32'd19340: dataIn1 = 32'd748
; 
32'd19341: dataIn1 = 32'd753
; 
32'd19342: dataIn1 = 32'd755
; 
32'd19343: dataIn1 = 32'd759
; 
32'd19344: dataIn1 = 32'd761
; 
32'd19345: dataIn1 = 32'd796
; 
32'd19346: dataIn1 = 32'd299
; 
32'd19347: dataIn1 = 32'd300
; 
32'd19348: dataIn1 = 32'd303
; 
32'd19349: dataIn1 = 32'd336
; 
32'd19350: dataIn1 = 32'd355
; 
32'd19351: dataIn1 = 32'd377
; 
32'd19352: dataIn1 = 32'd382
; 
32'd19353: dataIn1 = 32'd394
; 
32'd19354: dataIn1 = 32'd397
; 
32'd19355: dataIn1 = 32'd408
; 
32'd19356: dataIn1 = 32'd421
; 
32'd19357: dataIn1 = 32'd422
; 
32'd19358: dataIn1 = 32'd434
; 
32'd19359: dataIn1 = 32'd439
; 
32'd19360: dataIn1 = 32'd447
; 
32'd19361: dataIn1 = 32'd475
; 
32'd19362: dataIn1 = 32'd500
; 
32'd19363: dataIn1 = 32'd507
; 
32'd19364: dataIn1 = 32'd572
; 
32'd19365: dataIn1 = 32'd579
; 
32'd19366: dataIn1 = 32'd607
; 
32'd19367: dataIn1 = 32'd642
; 
32'd19368: dataIn1 = 32'd665
; 
32'd19369: dataIn1 = 32'd669
; 
32'd19370: dataIn1 = 32'd678
; 
32'd19371: dataIn1 = 32'd697
; 
32'd19372: dataIn1 = 32'd709
; 
32'd19373: dataIn1 = 32'd714
; 
32'd19374: dataIn1 = 32'd715
; 
32'd19375: dataIn1 = 32'd728
; 
32'd19376: dataIn1 = 32'd766
; 
32'd19377: dataIn1 = 32'd296
; 
32'd19378: dataIn1 = 32'd320
; 
32'd19379: dataIn1 = 32'd327
; 
32'd19380: dataIn1 = 32'd336
; 
32'd19381: dataIn1 = 32'd349
; 
32'd19382: dataIn1 = 32'd359
; 
32'd19383: dataIn1 = 32'd364
; 
32'd19384: dataIn1 = 32'd394
; 
32'd19385: dataIn1 = 32'd419
; 
32'd19386: dataIn1 = 32'd480
; 
32'd19387: dataIn1 = 32'd482
; 
32'd19388: dataIn1 = 32'd490
; 
32'd19389: dataIn1 = 32'd560
; 
32'd19390: dataIn1 = 32'd570
; 
32'd19391: dataIn1 = 32'd575
; 
32'd19392: dataIn1 = 32'd599
; 
32'd19393: dataIn1 = 32'd605
; 
32'd19394: dataIn1 = 32'd611
; 
32'd19395: dataIn1 = 32'd615
; 
32'd19396: dataIn1 = 32'd640
; 
32'd19397: dataIn1 = 32'd661
; 
32'd19398: dataIn1 = 32'd676
; 
32'd19399: dataIn1 = 32'd683
; 
32'd19400: dataIn1 = 32'd711
; 
32'd19401: dataIn1 = 32'd744
; 
32'd19402: dataIn1 = 32'd751
; 
32'd19403: dataIn1 = 32'd334
; 
32'd19404: dataIn1 = 32'd335
; 
32'd19405: dataIn1 = 32'd341
; 
32'd19406: dataIn1 = 32'd351
; 
32'd19407: dataIn1 = 32'd365
; 
32'd19408: dataIn1 = 32'd406
; 
32'd19409: dataIn1 = 32'd440
; 
32'd19410: dataIn1 = 32'd463
; 
32'd19411: dataIn1 = 32'd495
; 
32'd19412: dataIn1 = 32'd501
; 
32'd19413: dataIn1 = 32'd513
; 
32'd19414: dataIn1 = 32'd515
; 
32'd19415: dataIn1 = 32'd546
; 
32'd19416: dataIn1 = 32'd561
; 
32'd19417: dataIn1 = 32'd569
; 
32'd19418: dataIn1 = 32'd574
; 
32'd19419: dataIn1 = 32'd600
; 
32'd19420: dataIn1 = 32'd625
; 
32'd19421: dataIn1 = 32'd637
; 
32'd19422: dataIn1 = 32'd660
; 
32'd19423: dataIn1 = 32'd669
; 
32'd19424: dataIn1 = 32'd714
; 
32'd19425: dataIn1 = 32'd763
; 
32'd19426: dataIn1 = 32'd769
; 
32'd19427: dataIn1 = 32'd784
; 
32'd19428: dataIn1 = 32'd786
; 
32'd19429: dataIn1 = 32'd787
; 
32'd19430: dataIn1 = 32'd295
; 
32'd19431: dataIn1 = 32'd297
; 
32'd19432: dataIn1 = 32'd346
; 
32'd19433: dataIn1 = 32'd352
; 
32'd19434: dataIn1 = 32'd359
; 
32'd19435: dataIn1 = 32'd366
; 
32'd19436: dataIn1 = 32'd369
; 
32'd19437: dataIn1 = 32'd422
; 
32'd19438: dataIn1 = 32'd455
; 
32'd19439: dataIn1 = 32'd468
; 
32'd19440: dataIn1 = 32'd477
; 
32'd19441: dataIn1 = 32'd486
; 
32'd19442: dataIn1 = 32'd511
; 
32'd19443: dataIn1 = 32'd515
; 
32'd19444: dataIn1 = 32'd540
; 
32'd19445: dataIn1 = 32'd544
; 
32'd19446: dataIn1 = 32'd564
; 
32'd19447: dataIn1 = 32'd576
; 
32'd19448: dataIn1 = 32'd579
; 
32'd19449: dataIn1 = 32'd598
; 
32'd19450: dataIn1 = 32'd623
; 
32'd19451: dataIn1 = 32'd641
; 
32'd19452: dataIn1 = 32'd657
; 
32'd19453: dataIn1 = 32'd666
; 
32'd19454: dataIn1 = 32'd719
; 
32'd19455: dataIn1 = 32'd724
; 
32'd19456: dataIn1 = 32'd754
; 
32'd19457: dataIn1 = 32'd765
; 
32'd19458: dataIn1 = 32'd766
; 
32'd19459: dataIn1 = 32'd798
; 
32'd19460: dataIn1 = 32'd305
; 
32'd19461: dataIn1 = 32'd353
; 
32'd19462: dataIn1 = 32'd357
; 
32'd19463: dataIn1 = 32'd370
; 
32'd19464: dataIn1 = 32'd380
; 
32'd19465: dataIn1 = 32'd397
; 
32'd19466: dataIn1 = 32'd400
; 
32'd19467: dataIn1 = 32'd403
; 
32'd19468: dataIn1 = 32'd443
; 
32'd19469: dataIn1 = 32'd476
; 
32'd19470: dataIn1 = 32'd482
; 
32'd19471: dataIn1 = 32'd492
; 
32'd19472: dataIn1 = 32'd512
; 
32'd19473: dataIn1 = 32'd530
; 
32'd19474: dataIn1 = 32'd535
; 
32'd19475: dataIn1 = 32'd536
; 
32'd19476: dataIn1 = 32'd592
; 
32'd19477: dataIn1 = 32'd644
; 
32'd19478: dataIn1 = 32'd647
; 
32'd19479: dataIn1 = 32'd652
; 
32'd19480: dataIn1 = 32'd698
; 
32'd19481: dataIn1 = 32'd705
; 
32'd19482: dataIn1 = 32'd718
; 
32'd19483: dataIn1 = 32'd723
; 
32'd19484: dataIn1 = 32'd767
; 
32'd19485: dataIn1 = 32'd774
; 
32'd19486: dataIn1 = 32'd791
; 
32'd19487: dataIn1 = 32'd295
; 
32'd19488: dataIn1 = 32'd302
; 
32'd19489: dataIn1 = 32'd329
; 
32'd19490: dataIn1 = 32'd355
; 
32'd19491: dataIn1 = 32'd356
; 
32'd19492: dataIn1 = 32'd362
; 
32'd19493: dataIn1 = 32'd368
; 
32'd19494: dataIn1 = 32'd372
; 
32'd19495: dataIn1 = 32'd398
; 
32'd19496: dataIn1 = 32'd401
; 
32'd19497: dataIn1 = 32'd412
; 
32'd19498: dataIn1 = 32'd431
; 
32'd19499: dataIn1 = 32'd434
; 
32'd19500: dataIn1 = 32'd442
; 
32'd19501: dataIn1 = 32'd448
; 
32'd19502: dataIn1 = 32'd506
; 
32'd19503: dataIn1 = 32'd538
; 
32'd19504: dataIn1 = 32'd550
; 
32'd19505: dataIn1 = 32'd558
; 
32'd19506: dataIn1 = 32'd561
; 
32'd19507: dataIn1 = 32'd563
; 
32'd19508: dataIn1 = 32'd584
; 
32'd19509: dataIn1 = 32'd587
; 
32'd19510: dataIn1 = 32'd620
; 
32'd19511: dataIn1 = 32'd627
; 
32'd19512: dataIn1 = 32'd634
; 
32'd19513: dataIn1 = 32'd646
; 
32'd19514: dataIn1 = 32'd667
; 
32'd19515: dataIn1 = 32'd675
; 
32'd19516: dataIn1 = 32'd697
; 
32'd19517: dataIn1 = 32'd722
; 
32'd19518: dataIn1 = 32'd732
; 
32'd19519: dataIn1 = 32'd794
; 
32'd19520: dataIn1 = 32'd304
; 
32'd19521: dataIn1 = 32'd310
; 
32'd19522: dataIn1 = 32'd313
; 
32'd19523: dataIn1 = 32'd353
; 
32'd19524: dataIn1 = 32'd396
; 
32'd19525: dataIn1 = 32'd410
; 
32'd19526: dataIn1 = 32'd464
; 
32'd19527: dataIn1 = 32'd470
; 
32'd19528: dataIn1 = 32'd506
; 
32'd19529: dataIn1 = 32'd545
; 
32'd19530: dataIn1 = 32'd546
; 
32'd19531: dataIn1 = 32'd562
; 
32'd19532: dataIn1 = 32'd594
; 
32'd19533: dataIn1 = 32'd600
; 
32'd19534: dataIn1 = 32'd631
; 
32'd19535: dataIn1 = 32'd646
; 
32'd19536: dataIn1 = 32'd656
; 
32'd19537: dataIn1 = 32'd696
; 
32'd19538: dataIn1 = 32'd721
; 
32'd19539: dataIn1 = 32'd755
; 
32'd19540: dataIn1 = 32'd769
; 
32'd19541: dataIn1 = 32'd770
; 
32'd19542: dataIn1 = 32'd776
; 
32'd19543: dataIn1 = 32'd787
; 
32'd19544: dataIn1 = 32'd791
; 
32'd19545: dataIn1 = 32'd795
; 
32'd19546: dataIn1 = 32'd356
; 
32'd19547: dataIn1 = 32'd397
; 
32'd19548: dataIn1 = 32'd417
; 
32'd19549: dataIn1 = 32'd421
; 
32'd19550: dataIn1 = 32'd468
; 
32'd19551: dataIn1 = 32'd469
; 
32'd19552: dataIn1 = 32'd472
; 
32'd19553: dataIn1 = 32'd482
; 
32'd19554: dataIn1 = 32'd490
; 
32'd19555: dataIn1 = 32'd525
; 
32'd19556: dataIn1 = 32'd541
; 
32'd19557: dataIn1 = 32'd608
; 
32'd19558: dataIn1 = 32'd610
; 
32'd19559: dataIn1 = 32'd612
; 
32'd19560: dataIn1 = 32'd623
; 
32'd19561: dataIn1 = 32'd625
; 
32'd19562: dataIn1 = 32'd632
; 
32'd19563: dataIn1 = 32'd653
; 
32'd19564: dataIn1 = 32'd660
; 
32'd19565: dataIn1 = 32'd716
; 
32'd19566: dataIn1 = 32'd720
; 
32'd19567: dataIn1 = 32'd726
; 
32'd19568: dataIn1 = 32'd737
; 
32'd19569: dataIn1 = 32'd742
; 
32'd19570: dataIn1 = 32'd792
; 
32'd19571: dataIn1 = 32'd794
; 
32'd19572: dataIn1 = 32'd301
; 
32'd19573: dataIn1 = 32'd319
; 
32'd19574: dataIn1 = 32'd343
; 
32'd19575: dataIn1 = 32'd344
; 
32'd19576: dataIn1 = 32'd366
; 
32'd19577: dataIn1 = 32'd370
; 
32'd19578: dataIn1 = 32'd379
; 
32'd19579: dataIn1 = 32'd380
; 
32'd19580: dataIn1 = 32'd386
; 
32'd19581: dataIn1 = 32'd432
; 
32'd19582: dataIn1 = 32'd439
; 
32'd19583: dataIn1 = 32'd466
; 
32'd19584: dataIn1 = 32'd482
; 
32'd19585: dataIn1 = 32'd491
; 
32'd19586: dataIn1 = 32'd495
; 
32'd19587: dataIn1 = 32'd499
; 
32'd19588: dataIn1 = 32'd534
; 
32'd19589: dataIn1 = 32'd542
; 
32'd19590: dataIn1 = 32'd592
; 
32'd19591: dataIn1 = 32'd605
; 
32'd19592: dataIn1 = 32'd624
; 
32'd19593: dataIn1 = 32'd629
; 
32'd19594: dataIn1 = 32'd638
; 
32'd19595: dataIn1 = 32'd649
; 
32'd19596: dataIn1 = 32'd682
; 
32'd19597: dataIn1 = 32'd685
; 
32'd19598: dataIn1 = 32'd686
; 
32'd19599: dataIn1 = 32'd693
; 
32'd19600: dataIn1 = 32'd695
; 
32'd19601: dataIn1 = 32'd746
; 
32'd19602: dataIn1 = 32'd758
; 
32'd19603: dataIn1 = 32'd766
; 
32'd19604: dataIn1 = 32'd767
; 
32'd19605: dataIn1 = 32'd772
; 
32'd19606: dataIn1 = 32'd305
; 
32'd19607: dataIn1 = 32'd327
; 
32'd19608: dataIn1 = 32'd334
; 
32'd19609: dataIn1 = 32'd340
; 
32'd19610: dataIn1 = 32'd341
; 
32'd19611: dataIn1 = 32'd402
; 
32'd19612: dataIn1 = 32'd406
; 
32'd19613: dataIn1 = 32'd419
; 
32'd19614: dataIn1 = 32'd491
; 
32'd19615: dataIn1 = 32'd509
; 
32'd19616: dataIn1 = 32'd534
; 
32'd19617: dataIn1 = 32'd557
; 
32'd19618: dataIn1 = 32'd603
; 
32'd19619: dataIn1 = 32'd609
; 
32'd19620: dataIn1 = 32'd614
; 
32'd19621: dataIn1 = 32'd621
; 
32'd19622: dataIn1 = 32'd682
; 
32'd19623: dataIn1 = 32'd686
; 
32'd19624: dataIn1 = 32'd691
; 
32'd19625: dataIn1 = 32'd694
; 
32'd19626: dataIn1 = 32'd751
; 
32'd19627: dataIn1 = 32'd778
; 
32'd19628: dataIn1 = 32'd779
; 
32'd19629: dataIn1 = 32'd306
; 
32'd19630: dataIn1 = 32'd316
; 
32'd19631: dataIn1 = 32'd319
; 
32'd19632: dataIn1 = 32'd384
; 
32'd19633: dataIn1 = 32'd425
; 
32'd19634: dataIn1 = 32'd446
; 
32'd19635: dataIn1 = 32'd457
; 
32'd19636: dataIn1 = 32'd468
; 
32'd19637: dataIn1 = 32'd487
; 
32'd19638: dataIn1 = 32'd493
; 
32'd19639: dataIn1 = 32'd513
; 
32'd19640: dataIn1 = 32'd556
; 
32'd19641: dataIn1 = 32'd580
; 
32'd19642: dataIn1 = 32'd601
; 
32'd19643: dataIn1 = 32'd680
; 
32'd19644: dataIn1 = 32'd736
; 
32'd19645: dataIn1 = 32'd768
; 
32'd19646: dataIn1 = 32'd792
; 
32'd19647: dataIn1 = 32'd312
; 
32'd19648: dataIn1 = 32'd315
; 
32'd19649: dataIn1 = 32'd337
; 
32'd19650: dataIn1 = 32'd380
; 
32'd19651: dataIn1 = 32'd392
; 
32'd19652: dataIn1 = 32'd399
; 
32'd19653: dataIn1 = 32'd402
; 
32'd19654: dataIn1 = 32'd406
; 
32'd19655: dataIn1 = 32'd410
; 
32'd19656: dataIn1 = 32'd425
; 
32'd19657: dataIn1 = 32'd503
; 
32'd19658: dataIn1 = 32'd526
; 
32'd19659: dataIn1 = 32'd547
; 
32'd19660: dataIn1 = 32'd560
; 
32'd19661: dataIn1 = 32'd571
; 
32'd19662: dataIn1 = 32'd576
; 
32'd19663: dataIn1 = 32'd596
; 
32'd19664: dataIn1 = 32'd609
; 
32'd19665: dataIn1 = 32'd626
; 
32'd19666: dataIn1 = 32'd652
; 
32'd19667: dataIn1 = 32'd703
; 
32'd19668: dataIn1 = 32'd706
; 
32'd19669: dataIn1 = 32'd708
; 
32'd19670: dataIn1 = 32'd731
; 
32'd19671: dataIn1 = 32'd736
; 
32'd19672: dataIn1 = 32'd741
; 
32'd19673: dataIn1 = 32'd325
; 
32'd19674: dataIn1 = 32'd327
; 
32'd19675: dataIn1 = 32'd334
; 
32'd19676: dataIn1 = 32'd416
; 
32'd19677: dataIn1 = 32'd449
; 
32'd19678: dataIn1 = 32'd472
; 
32'd19679: dataIn1 = 32'd484
; 
32'd19680: dataIn1 = 32'd491
; 
32'd19681: dataIn1 = 32'd530
; 
32'd19682: dataIn1 = 32'd532
; 
32'd19683: dataIn1 = 32'd571
; 
32'd19684: dataIn1 = 32'd584
; 
32'd19685: dataIn1 = 32'd622
; 
32'd19686: dataIn1 = 32'd646
; 
32'd19687: dataIn1 = 32'd648
; 
32'd19688: dataIn1 = 32'd651
; 
32'd19689: dataIn1 = 32'd655
; 
32'd19690: dataIn1 = 32'd656
; 
32'd19691: dataIn1 = 32'd668
; 
32'd19692: dataIn1 = 32'd707
; 
32'd19693: dataIn1 = 32'd720
; 
32'd19694: dataIn1 = 32'd739
; 
32'd19695: dataIn1 = 32'd777
; 
32'd19696: dataIn1 = 32'd783
; 
32'd19697: dataIn1 = 32'd795
; 
32'd19698: dataIn1 = 32'd800
; 
32'd19699: dataIn1 = 32'd311
; 
32'd19700: dataIn1 = 32'd315
; 
32'd19701: dataIn1 = 32'd316
; 
32'd19702: dataIn1 = 32'd339
; 
32'd19703: dataIn1 = 32'd343
; 
32'd19704: dataIn1 = 32'd349
; 
32'd19705: dataIn1 = 32'd362
; 
32'd19706: dataIn1 = 32'd378
; 
32'd19707: dataIn1 = 32'd386
; 
32'd19708: dataIn1 = 32'd387
; 
32'd19709: dataIn1 = 32'd406
; 
32'd19710: dataIn1 = 32'd421
; 
32'd19711: dataIn1 = 32'd443
; 
32'd19712: dataIn1 = 32'd448
; 
32'd19713: dataIn1 = 32'd449
; 
32'd19714: dataIn1 = 32'd461
; 
32'd19715: dataIn1 = 32'd468
; 
32'd19716: dataIn1 = 32'd511
; 
32'd19717: dataIn1 = 32'd521
; 
32'd19718: dataIn1 = 32'd523
; 
32'd19719: dataIn1 = 32'd549
; 
32'd19720: dataIn1 = 32'd559
; 
32'd19721: dataIn1 = 32'd561
; 
32'd19722: dataIn1 = 32'd568
; 
32'd19723: dataIn1 = 32'd591
; 
32'd19724: dataIn1 = 32'd592
; 
32'd19725: dataIn1 = 32'd661
; 
32'd19726: dataIn1 = 32'd662
; 
32'd19727: dataIn1 = 32'd673
; 
32'd19728: dataIn1 = 32'd688
; 
32'd19729: dataIn1 = 32'd693
; 
32'd19730: dataIn1 = 32'd696
; 
32'd19731: dataIn1 = 32'd711
; 
32'd19732: dataIn1 = 32'd720
; 
32'd19733: dataIn1 = 32'd756
; 
32'd19734: dataIn1 = 32'd758
; 
32'd19735: dataIn1 = 32'd765
; 
32'd19736: dataIn1 = 32'd787
; 
32'd19737: dataIn1 = 32'd790
; 
32'd19738: dataIn1 = 32'd337
; 
32'd19739: dataIn1 = 32'd344
; 
32'd19740: dataIn1 = 32'd360
; 
32'd19741: dataIn1 = 32'd365
; 
32'd19742: dataIn1 = 32'd380
; 
32'd19743: dataIn1 = 32'd416
; 
32'd19744: dataIn1 = 32'd446
; 
32'd19745: dataIn1 = 32'd454
; 
32'd19746: dataIn1 = 32'd471
; 
32'd19747: dataIn1 = 32'd487
; 
32'd19748: dataIn1 = 32'd501
; 
32'd19749: dataIn1 = 32'd506
; 
32'd19750: dataIn1 = 32'd516
; 
32'd19751: dataIn1 = 32'd528
; 
32'd19752: dataIn1 = 32'd535
; 
32'd19753: dataIn1 = 32'd537
; 
32'd19754: dataIn1 = 32'd560
; 
32'd19755: dataIn1 = 32'd626
; 
32'd19756: dataIn1 = 32'd656
; 
32'd19757: dataIn1 = 32'd666
; 
32'd19758: dataIn1 = 32'd674
; 
32'd19759: dataIn1 = 32'd690
; 
32'd19760: dataIn1 = 32'd709
; 
32'd19761: dataIn1 = 32'd746
; 
32'd19762: dataIn1 = 32'd787
; 
32'd19763: dataIn1 = 32'd304
; 
32'd19764: dataIn1 = 32'd316
; 
32'd19765: dataIn1 = 32'd321
; 
32'd19766: dataIn1 = 32'd327
; 
32'd19767: dataIn1 = 32'd342
; 
32'd19768: dataIn1 = 32'd353
; 
32'd19769: dataIn1 = 32'd369
; 
32'd19770: dataIn1 = 32'd388
; 
32'd19771: dataIn1 = 32'd389
; 
32'd19772: dataIn1 = 32'd433
; 
32'd19773: dataIn1 = 32'd440
; 
32'd19774: dataIn1 = 32'd450
; 
32'd19775: dataIn1 = 32'd466
; 
32'd19776: dataIn1 = 32'd474
; 
32'd19777: dataIn1 = 32'd476
; 
32'd19778: dataIn1 = 32'd531
; 
32'd19779: dataIn1 = 32'd554
; 
32'd19780: dataIn1 = 32'd598
; 
32'd19781: dataIn1 = 32'd602
; 
32'd19782: dataIn1 = 32'd621
; 
32'd19783: dataIn1 = 32'd655
; 
32'd19784: dataIn1 = 32'd664
; 
32'd19785: dataIn1 = 32'd687
; 
32'd19786: dataIn1 = 32'd693
; 
32'd19787: dataIn1 = 32'd705
; 
32'd19788: dataIn1 = 32'd750
; 
32'd19789: dataIn1 = 32'd760
; 
32'd19790: dataIn1 = 32'd769
; 
32'd19791: dataIn1 = 32'd770
; 
32'd19792: dataIn1 = 32'd791
; 
32'd19793: dataIn1 = 32'd797
; 
32'd19794: dataIn1 = 32'd320
; 
32'd19795: dataIn1 = 32'd422
; 
32'd19796: dataIn1 = 32'd438
; 
32'd19797: dataIn1 = 32'd447
; 
32'd19798: dataIn1 = 32'd474
; 
32'd19799: dataIn1 = 32'd492
; 
32'd19800: dataIn1 = 32'd508
; 
32'd19801: dataIn1 = 32'd516
; 
32'd19802: dataIn1 = 32'd545
; 
32'd19803: dataIn1 = 32'd555
; 
32'd19804: dataIn1 = 32'd575
; 
32'd19805: dataIn1 = 32'd582
; 
32'd19806: dataIn1 = 32'd584
; 
32'd19807: dataIn1 = 32'd611
; 
32'd19808: dataIn1 = 32'd614
; 
32'd19809: dataIn1 = 32'd636
; 
32'd19810: dataIn1 = 32'd644
; 
32'd19811: dataIn1 = 32'd656
; 
32'd19812: dataIn1 = 32'd661
; 
32'd19813: dataIn1 = 32'd670
; 
32'd19814: dataIn1 = 32'd674
; 
32'd19815: dataIn1 = 32'd695
; 
32'd19816: dataIn1 = 32'd700
; 
32'd19817: dataIn1 = 32'd723
; 
32'd19818: dataIn1 = 32'd727
; 
32'd19819: dataIn1 = 32'd737
; 
32'd19820: dataIn1 = 32'd763
; 
32'd19821: dataIn1 = 32'd777
; 
32'd19822: dataIn1 = 32'd318
; 
32'd19823: dataIn1 = 32'd338
; 
32'd19824: dataIn1 = 32'd351
; 
32'd19825: dataIn1 = 32'd353
; 
32'd19826: dataIn1 = 32'd361
; 
32'd19827: dataIn1 = 32'd369
; 
32'd19828: dataIn1 = 32'd375
; 
32'd19829: dataIn1 = 32'd384
; 
32'd19830: dataIn1 = 32'd398
; 
32'd19831: dataIn1 = 32'd405
; 
32'd19832: dataIn1 = 32'd431
; 
32'd19833: dataIn1 = 32'd497
; 
32'd19834: dataIn1 = 32'd498
; 
32'd19835: dataIn1 = 32'd516
; 
32'd19836: dataIn1 = 32'd548
; 
32'd19837: dataIn1 = 32'd551
; 
32'd19838: dataIn1 = 32'd564
; 
32'd19839: dataIn1 = 32'd577
; 
32'd19840: dataIn1 = 32'd579
; 
32'd19841: dataIn1 = 32'd580
; 
32'd19842: dataIn1 = 32'd593
; 
32'd19843: dataIn1 = 32'd614
; 
32'd19844: dataIn1 = 32'd667
; 
32'd19845: dataIn1 = 32'd675
; 
32'd19846: dataIn1 = 32'd704
; 
32'd19847: dataIn1 = 32'd716
; 
32'd19848: dataIn1 = 32'd719
; 
32'd19849: dataIn1 = 32'd741
; 
32'd19850: dataIn1 = 32'd760
; 
32'd19851: dataIn1 = 32'd764
; 
32'd19852: dataIn1 = 32'd769
; 
32'd19853: dataIn1 = 32'd320
; 
32'd19854: dataIn1 = 32'd327
; 
32'd19855: dataIn1 = 32'd328
; 
32'd19856: dataIn1 = 32'd337
; 
32'd19857: dataIn1 = 32'd343
; 
32'd19858: dataIn1 = 32'd373
; 
32'd19859: dataIn1 = 32'd375
; 
32'd19860: dataIn1 = 32'd384
; 
32'd19861: dataIn1 = 32'd395
; 
32'd19862: dataIn1 = 32'd419
; 
32'd19863: dataIn1 = 32'd427
; 
32'd19864: dataIn1 = 32'd430
; 
32'd19865: dataIn1 = 32'd432
; 
32'd19866: dataIn1 = 32'd441
; 
32'd19867: dataIn1 = 32'd455
; 
32'd19868: dataIn1 = 32'd470
; 
32'd19869: dataIn1 = 32'd494
; 
32'd19870: dataIn1 = 32'd495
; 
32'd19871: dataIn1 = 32'd539
; 
32'd19872: dataIn1 = 32'd546
; 
32'd19873: dataIn1 = 32'd560
; 
32'd19874: dataIn1 = 32'd561
; 
32'd19875: dataIn1 = 32'd627
; 
32'd19876: dataIn1 = 32'd637
; 
32'd19877: dataIn1 = 32'd645
; 
32'd19878: dataIn1 = 32'd659
; 
32'd19879: dataIn1 = 32'd661
; 
32'd19880: dataIn1 = 32'd675
; 
32'd19881: dataIn1 = 32'd684
; 
32'd19882: dataIn1 = 32'd685
; 
32'd19883: dataIn1 = 32'd727
; 
32'd19884: dataIn1 = 32'd729
; 
32'd19885: dataIn1 = 32'd746
; 
32'd19886: dataIn1 = 32'd775
; 
32'd19887: dataIn1 = 32'd776
; 
32'd19888: dataIn1 = 32'd782
; 
32'd19889: dataIn1 = 32'd800
; 
32'd19890: dataIn1 = 32'd316
; 
32'd19891: dataIn1 = 32'd325
; 
32'd19892: dataIn1 = 32'd336
; 
32'd19893: dataIn1 = 32'd345
; 
32'd19894: dataIn1 = 32'd366
; 
32'd19895: dataIn1 = 32'd370
; 
32'd19896: dataIn1 = 32'd382
; 
32'd19897: dataIn1 = 32'd397
; 
32'd19898: dataIn1 = 32'd439
; 
32'd19899: dataIn1 = 32'd463
; 
32'd19900: dataIn1 = 32'd476
; 
32'd19901: dataIn1 = 32'd492
; 
32'd19902: dataIn1 = 32'd520
; 
32'd19903: dataIn1 = 32'd534
; 
32'd19904: dataIn1 = 32'd542
; 
32'd19905: dataIn1 = 32'd549
; 
32'd19906: dataIn1 = 32'd566
; 
32'd19907: dataIn1 = 32'd591
; 
32'd19908: dataIn1 = 32'd608
; 
32'd19909: dataIn1 = 32'd614
; 
32'd19910: dataIn1 = 32'd621
; 
32'd19911: dataIn1 = 32'd623
; 
32'd19912: dataIn1 = 32'd655
; 
32'd19913: dataIn1 = 32'd672
; 
32'd19914: dataIn1 = 32'd674
; 
32'd19915: dataIn1 = 32'd712
; 
32'd19916: dataIn1 = 32'd762
; 
32'd19917: dataIn1 = 32'd783
; 
32'd19918: dataIn1 = 32'd785
; 
32'd19919: dataIn1 = 32'd320
; 
32'd19920: dataIn1 = 32'd345
; 
32'd19921: dataIn1 = 32'd394
; 
32'd19922: dataIn1 = 32'd415
; 
32'd19923: dataIn1 = 32'd421
; 
32'd19924: dataIn1 = 32'd440
; 
32'd19925: dataIn1 = 32'd460
; 
32'd19926: dataIn1 = 32'd482
; 
32'd19927: dataIn1 = 32'd491
; 
32'd19928: dataIn1 = 32'd568
; 
32'd19929: dataIn1 = 32'd574
; 
32'd19930: dataIn1 = 32'd601
; 
32'd19931: dataIn1 = 32'd664
; 
32'd19932: dataIn1 = 32'd668
; 
32'd19933: dataIn1 = 32'd672
; 
32'd19934: dataIn1 = 32'd683
; 
32'd19935: dataIn1 = 32'd728
; 
32'd19936: dataIn1 = 32'd733
; 
32'd19937: dataIn1 = 32'd737
; 
32'd19938: dataIn1 = 32'd741
; 
32'd19939: dataIn1 = 32'd744
; 
32'd19940: dataIn1 = 32'd799
; 
32'd19941: dataIn1 = 32'd328
; 
32'd19942: dataIn1 = 32'd338
; 
32'd19943: dataIn1 = 32'd345
; 
32'd19944: dataIn1 = 32'd347
; 
32'd19945: dataIn1 = 32'd360
; 
32'd19946: dataIn1 = 32'd370
; 
32'd19947: dataIn1 = 32'd388
; 
32'd19948: dataIn1 = 32'd418
; 
32'd19949: dataIn1 = 32'd441
; 
32'd19950: dataIn1 = 32'd442
; 
32'd19951: dataIn1 = 32'd461
; 
32'd19952: dataIn1 = 32'd468
; 
32'd19953: dataIn1 = 32'd469
; 
32'd19954: dataIn1 = 32'd485
; 
32'd19955: dataIn1 = 32'd517
; 
32'd19956: dataIn1 = 32'd519
; 
32'd19957: dataIn1 = 32'd525
; 
32'd19958: dataIn1 = 32'd534
; 
32'd19959: dataIn1 = 32'd541
; 
32'd19960: dataIn1 = 32'd559
; 
32'd19961: dataIn1 = 32'd571
; 
32'd19962: dataIn1 = 32'd577
; 
32'd19963: dataIn1 = 32'd594
; 
32'd19964: dataIn1 = 32'd673
; 
32'd19965: dataIn1 = 32'd687
; 
32'd19966: dataIn1 = 32'd691
; 
32'd19967: dataIn1 = 32'd714
; 
32'd19968: dataIn1 = 32'd756
; 
32'd19969: dataIn1 = 32'd794
; 
32'd19970: dataIn1 = 32'd314
; 
32'd19971: dataIn1 = 32'd337
; 
32'd19972: dataIn1 = 32'd354
; 
32'd19973: dataIn1 = 32'd356
; 
32'd19974: dataIn1 = 32'd359
; 
32'd19975: dataIn1 = 32'd383
; 
32'd19976: dataIn1 = 32'd386
; 
32'd19977: dataIn1 = 32'd422
; 
32'd19978: dataIn1 = 32'd440
; 
32'd19979: dataIn1 = 32'd500
; 
32'd19980: dataIn1 = 32'd507
; 
32'd19981: dataIn1 = 32'd509
; 
32'd19982: dataIn1 = 32'd521
; 
32'd19983: dataIn1 = 32'd526
; 
32'd19984: dataIn1 = 32'd528
; 
32'd19985: dataIn1 = 32'd536
; 
32'd19986: dataIn1 = 32'd546
; 
32'd19987: dataIn1 = 32'd579
; 
32'd19988: dataIn1 = 32'd596
; 
32'd19989: dataIn1 = 32'd599
; 
32'd19990: dataIn1 = 32'd611
; 
32'd19991: dataIn1 = 32'd630
; 
32'd19992: dataIn1 = 32'd631
; 
32'd19993: dataIn1 = 32'd636
; 
32'd19994: dataIn1 = 32'd642
; 
32'd19995: dataIn1 = 32'd671
; 
32'd19996: dataIn1 = 32'd677
; 
32'd19997: dataIn1 = 32'd681
; 
32'd19998: dataIn1 = 32'd700
; 
32'd19999: dataIn1 = 32'd708
; 
32'd20000: dataIn1 = 32'd718
; 
32'd20001: dataIn1 = 32'd733
; 
32'd20002: dataIn1 = 32'd743
; 
32'd20003: dataIn1 = 32'd759
; 
32'd20004: dataIn1 = 32'd774
; 
32'd20005: dataIn1 = 32'd783
; 
32'd20006: dataIn1 = 32'd317
; 
32'd20007: dataIn1 = 32'd326
; 
32'd20008: dataIn1 = 32'd330
; 
32'd20009: dataIn1 = 32'd348
; 
32'd20010: dataIn1 = 32'd374
; 
32'd20011: dataIn1 = 32'd375
; 
32'd20012: dataIn1 = 32'd408
; 
32'd20013: dataIn1 = 32'd409
; 
32'd20014: dataIn1 = 32'd413
; 
32'd20015: dataIn1 = 32'd420
; 
32'd20016: dataIn1 = 32'd430
; 
32'd20017: dataIn1 = 32'd431
; 
32'd20018: dataIn1 = 32'd446
; 
32'd20019: dataIn1 = 32'd480
; 
32'd20020: dataIn1 = 32'd496
; 
32'd20021: dataIn1 = 32'd500
; 
32'd20022: dataIn1 = 32'd526
; 
32'd20023: dataIn1 = 32'd535
; 
32'd20024: dataIn1 = 32'd536
; 
32'd20025: dataIn1 = 32'd550
; 
32'd20026: dataIn1 = 32'd555
; 
32'd20027: dataIn1 = 32'd558
; 
32'd20028: dataIn1 = 32'd567
; 
32'd20029: dataIn1 = 32'd577
; 
32'd20030: dataIn1 = 32'd596
; 
32'd20031: dataIn1 = 32'd632
; 
32'd20032: dataIn1 = 32'd645
; 
32'd20033: dataIn1 = 32'd647
; 
32'd20034: dataIn1 = 32'd649
; 
32'd20035: dataIn1 = 32'd675
; 
32'd20036: dataIn1 = 32'd682
; 
32'd20037: dataIn1 = 32'd705
; 
32'd20038: dataIn1 = 32'd714
; 
32'd20039: dataIn1 = 32'd766
; 
32'd20040: dataIn1 = 32'd312
; 
32'd20041: dataIn1 = 32'd330
; 
32'd20042: dataIn1 = 32'd340
; 
32'd20043: dataIn1 = 32'd343
; 
32'd20044: dataIn1 = 32'd353
; 
32'd20045: dataIn1 = 32'd375
; 
32'd20046: dataIn1 = 32'd382
; 
32'd20047: dataIn1 = 32'd448
; 
32'd20048: dataIn1 = 32'd458
; 
32'd20049: dataIn1 = 32'd474
; 
32'd20050: dataIn1 = 32'd475
; 
32'd20051: dataIn1 = 32'd503
; 
32'd20052: dataIn1 = 32'd542
; 
32'd20053: dataIn1 = 32'd548
; 
32'd20054: dataIn1 = 32'd572
; 
32'd20055: dataIn1 = 32'd591
; 
32'd20056: dataIn1 = 32'd618
; 
32'd20057: dataIn1 = 32'd622
; 
32'd20058: dataIn1 = 32'd645
; 
32'd20059: dataIn1 = 32'd649
; 
32'd20060: dataIn1 = 32'd658
; 
32'd20061: dataIn1 = 32'd668
; 
32'd20062: dataIn1 = 32'd674
; 
32'd20063: dataIn1 = 32'd677
; 
32'd20064: dataIn1 = 32'd683
; 
32'd20065: dataIn1 = 32'd690
; 
32'd20066: dataIn1 = 32'd692
; 
32'd20067: dataIn1 = 32'd722
; 
32'd20068: dataIn1 = 32'd739
; 
32'd20069: dataIn1 = 32'd750
; 
32'd20070: dataIn1 = 32'd758
; 
32'd20071: dataIn1 = 32'd779
; 
32'd20072: dataIn1 = 32'd781
; 
32'd20073: dataIn1 = 32'd791
; 
32'd20074: dataIn1 = 32'd343
; 
32'd20075: dataIn1 = 32'd368
; 
32'd20076: dataIn1 = 32'd383
; 
32'd20077: dataIn1 = 32'd388
; 
32'd20078: dataIn1 = 32'd425
; 
32'd20079: dataIn1 = 32'd442
; 
32'd20080: dataIn1 = 32'd464
; 
32'd20081: dataIn1 = 32'd479
; 
32'd20082: dataIn1 = 32'd483
; 
32'd20083: dataIn1 = 32'd501
; 
32'd20084: dataIn1 = 32'd531
; 
32'd20085: dataIn1 = 32'd534
; 
32'd20086: dataIn1 = 32'd545
; 
32'd20087: dataIn1 = 32'd550
; 
32'd20088: dataIn1 = 32'd576
; 
32'd20089: dataIn1 = 32'd615
; 
32'd20090: dataIn1 = 32'd625
; 
32'd20091: dataIn1 = 32'd629
; 
32'd20092: dataIn1 = 32'd643
; 
32'd20093: dataIn1 = 32'd654
; 
32'd20094: dataIn1 = 32'd668
; 
32'd20095: dataIn1 = 32'd713
; 
32'd20096: dataIn1 = 32'd731
; 
32'd20097: dataIn1 = 32'd734
; 
32'd20098: dataIn1 = 32'd742
; 
32'd20099: dataIn1 = 32'd752
; 
32'd20100: dataIn1 = 32'd753
; 
32'd20101: dataIn1 = 32'd756
; 
32'd20102: dataIn1 = 32'd758
; 
32'd20103: dataIn1 = 32'd772
; 
32'd20104: dataIn1 = 32'd332
; 
32'd20105: dataIn1 = 32'd349
; 
32'd20106: dataIn1 = 32'd351
; 
32'd20107: dataIn1 = 32'd393
; 
32'd20108: dataIn1 = 32'd412
; 
32'd20109: dataIn1 = 32'd418
; 
32'd20110: dataIn1 = 32'd430
; 
32'd20111: dataIn1 = 32'd458
; 
32'd20112: dataIn1 = 32'd461
; 
32'd20113: dataIn1 = 32'd484
; 
32'd20114: dataIn1 = 32'd504
; 
32'd20115: dataIn1 = 32'd505
; 
32'd20116: dataIn1 = 32'd519
; 
32'd20117: dataIn1 = 32'd537
; 
32'd20118: dataIn1 = 32'd543
; 
32'd20119: dataIn1 = 32'd571
; 
32'd20120: dataIn1 = 32'd591
; 
32'd20121: dataIn1 = 32'd605
; 
32'd20122: dataIn1 = 32'd623
; 
32'd20123: dataIn1 = 32'd639
; 
32'd20124: dataIn1 = 32'd649
; 
32'd20125: dataIn1 = 32'd681
; 
32'd20126: dataIn1 = 32'd694
; 
32'd20127: dataIn1 = 32'd704
; 
32'd20128: dataIn1 = 32'd707
; 
32'd20129: dataIn1 = 32'd718
; 
32'd20130: dataIn1 = 32'd736
; 
32'd20131: dataIn1 = 32'd741
; 
32'd20132: dataIn1 = 32'd766
; 
32'd20133: dataIn1 = 32'd314
; 
32'd20134: dataIn1 = 32'd333
; 
32'd20135: dataIn1 = 32'd338
; 
32'd20136: dataIn1 = 32'd370
; 
32'd20137: dataIn1 = 32'd440
; 
32'd20138: dataIn1 = 32'd456
; 
32'd20139: dataIn1 = 32'd461
; 
32'd20140: dataIn1 = 32'd469
; 
32'd20141: dataIn1 = 32'd498
; 
32'd20142: dataIn1 = 32'd499
; 
32'd20143: dataIn1 = 32'd575
; 
32'd20144: dataIn1 = 32'd604
; 
32'd20145: dataIn1 = 32'd628
; 
32'd20146: dataIn1 = 32'd667
; 
32'd20147: dataIn1 = 32'd669
; 
32'd20148: dataIn1 = 32'd672
; 
32'd20149: dataIn1 = 32'd693
; 
32'd20150: dataIn1 = 32'd711
; 
32'd20151: dataIn1 = 32'd774
; 
32'd20152: dataIn1 = 32'd778
; 
32'd20153: dataIn1 = 32'd791
; 
32'd20154: dataIn1 = 32'd792
; 
32'd20155: dataIn1 = 32'd323
; 
32'd20156: dataIn1 = 32'd329
; 
32'd20157: dataIn1 = 32'd349
; 
32'd20158: dataIn1 = 32'd364
; 
32'd20159: dataIn1 = 32'd392
; 
32'd20160: dataIn1 = 32'd416
; 
32'd20161: dataIn1 = 32'd458
; 
32'd20162: dataIn1 = 32'd464
; 
32'd20163: dataIn1 = 32'd471
; 
32'd20164: dataIn1 = 32'd473
; 
32'd20165: dataIn1 = 32'd490
; 
32'd20166: dataIn1 = 32'd498
; 
32'd20167: dataIn1 = 32'd502
; 
32'd20168: dataIn1 = 32'd530
; 
32'd20169: dataIn1 = 32'd564
; 
32'd20170: dataIn1 = 32'd579
; 
32'd20171: dataIn1 = 32'd586
; 
32'd20172: dataIn1 = 32'd604
; 
32'd20173: dataIn1 = 32'd626
; 
32'd20174: dataIn1 = 32'd635
; 
32'd20175: dataIn1 = 32'd648
; 
32'd20176: dataIn1 = 32'd657
; 
32'd20177: dataIn1 = 32'd673
; 
32'd20178: dataIn1 = 32'd692
; 
32'd20179: dataIn1 = 32'd706
; 
32'd20180: dataIn1 = 32'd709
; 
32'd20181: dataIn1 = 32'd736
; 
32'd20182: dataIn1 = 32'd740
; 
32'd20183: dataIn1 = 32'd750
; 
32'd20184: dataIn1 = 32'd773
; 
32'd20185: dataIn1 = 32'd783
; 
32'd20186: dataIn1 = 32'd339
; 
32'd20187: dataIn1 = 32'd345
; 
32'd20188: dataIn1 = 32'd358
; 
32'd20189: dataIn1 = 32'd388
; 
32'd20190: dataIn1 = 32'd406
; 
32'd20191: dataIn1 = 32'd408
; 
32'd20192: dataIn1 = 32'd431
; 
32'd20193: dataIn1 = 32'd442
; 
32'd20194: dataIn1 = 32'd446
; 
32'd20195: dataIn1 = 32'd452
; 
32'd20196: dataIn1 = 32'd459
; 
32'd20197: dataIn1 = 32'd469
; 
32'd20198: dataIn1 = 32'd487
; 
32'd20199: dataIn1 = 32'd492
; 
32'd20200: dataIn1 = 32'd514
; 
32'd20201: dataIn1 = 32'd582
; 
32'd20202: dataIn1 = 32'd602
; 
32'd20203: dataIn1 = 32'd615
; 
32'd20204: dataIn1 = 32'd618
; 
32'd20205: dataIn1 = 32'd624
; 
32'd20206: dataIn1 = 32'd629
; 
32'd20207: dataIn1 = 32'd656
; 
32'd20208: dataIn1 = 32'd678
; 
32'd20209: dataIn1 = 32'd682
; 
32'd20210: dataIn1 = 32'd683
; 
32'd20211: dataIn1 = 32'd696
; 
32'd20212: dataIn1 = 32'd708
; 
32'd20213: dataIn1 = 32'd720
; 
32'd20214: dataIn1 = 32'd728
; 
32'd20215: dataIn1 = 32'd736
; 
32'd20216: dataIn1 = 32'd748
; 
32'd20217: dataIn1 = 32'd749
; 
32'd20218: dataIn1 = 32'd754
; 
32'd20219: dataIn1 = 32'd779
; 
32'd20220: dataIn1 = 32'd786
; 
32'd20221: dataIn1 = 32'd789
; 
32'd20222: dataIn1 = 32'd792
; 
32'd20223: dataIn1 = 32'd319
; 
32'd20224: dataIn1 = 32'd350
; 
32'd20225: dataIn1 = 32'd352
; 
32'd20226: dataIn1 = 32'd357
; 
32'd20227: dataIn1 = 32'd367
; 
32'd20228: dataIn1 = 32'd420
; 
32'd20229: dataIn1 = 32'd429
; 
32'd20230: dataIn1 = 32'd446
; 
32'd20231: dataIn1 = 32'd451
; 
32'd20232: dataIn1 = 32'd454
; 
32'd20233: dataIn1 = 32'd473
; 
32'd20234: dataIn1 = 32'd496
; 
32'd20235: dataIn1 = 32'd500
; 
32'd20236: dataIn1 = 32'd514
; 
32'd20237: dataIn1 = 32'd515
; 
32'd20238: dataIn1 = 32'd528
; 
32'd20239: dataIn1 = 32'd550
; 
32'd20240: dataIn1 = 32'd555
; 
32'd20241: dataIn1 = 32'd565
; 
32'd20242: dataIn1 = 32'd571
; 
32'd20243: dataIn1 = 32'd582
; 
32'd20244: dataIn1 = 32'd592
; 
32'd20245: dataIn1 = 32'd609
; 
32'd20246: dataIn1 = 32'd616
; 
32'd20247: dataIn1 = 32'd622
; 
32'd20248: dataIn1 = 32'd629
; 
32'd20249: dataIn1 = 32'd635
; 
32'd20250: dataIn1 = 32'd637
; 
32'd20251: dataIn1 = 32'd666
; 
32'd20252: dataIn1 = 32'd675
; 
32'd20253: dataIn1 = 32'd682
; 
32'd20254: dataIn1 = 32'd709
; 
32'd20255: dataIn1 = 32'd724
; 
32'd20256: dataIn1 = 32'd738
; 
32'd20257: dataIn1 = 32'd760
; 
32'd20258: dataIn1 = 32'd772
; 
32'd20259: dataIn1 = 32'd336
; 
32'd20260: dataIn1 = 32'd367
; 
32'd20261: dataIn1 = 32'd380
; 
32'd20262: dataIn1 = 32'd383
; 
32'd20263: dataIn1 = 32'd402
; 
32'd20264: dataIn1 = 32'd418
; 
32'd20265: dataIn1 = 32'd437
; 
32'd20266: dataIn1 = 32'd438
; 
32'd20267: dataIn1 = 32'd446
; 
32'd20268: dataIn1 = 32'd450
; 
32'd20269: dataIn1 = 32'd472
; 
32'd20270: dataIn1 = 32'd503
; 
32'd20271: dataIn1 = 32'd543
; 
32'd20272: dataIn1 = 32'd577
; 
32'd20273: dataIn1 = 32'd677
; 
32'd20274: dataIn1 = 32'd688
; 
32'd20275: dataIn1 = 32'd716
; 
32'd20276: dataIn1 = 32'd727
; 
32'd20277: dataIn1 = 32'd752
; 
32'd20278: dataIn1 = 32'd770
; 
32'd20279: dataIn1 = 32'd783
; 
32'd20280: dataIn1 = 32'd794
; 
32'd20281: dataIn1 = 32'd796
; 
32'd20282: dataIn1 = 32'd319
; 
32'd20283: dataIn1 = 32'd326
; 
32'd20284: dataIn1 = 32'd400
; 
32'd20285: dataIn1 = 32'd432
; 
32'd20286: dataIn1 = 32'd438
; 
32'd20287: dataIn1 = 32'd489
; 
32'd20288: dataIn1 = 32'd493
; 
32'd20289: dataIn1 = 32'd502
; 
32'd20290: dataIn1 = 32'd522
; 
32'd20291: dataIn1 = 32'd572
; 
32'd20292: dataIn1 = 32'd575
; 
32'd20293: dataIn1 = 32'd581
; 
32'd20294: dataIn1 = 32'd582
; 
32'd20295: dataIn1 = 32'd592
; 
32'd20296: dataIn1 = 32'd616
; 
32'd20297: dataIn1 = 32'd638
; 
32'd20298: dataIn1 = 32'd651
; 
32'd20299: dataIn1 = 32'd696
; 
32'd20300: dataIn1 = 32'd782
; 
32'd20301: dataIn1 = 32'd783
; 
32'd20302: dataIn1 = 32'd784
; 
32'd20303: dataIn1 = 32'd786
; 
32'd20304: dataIn1 = 32'd795
; 
32'd20305: dataIn1 = 32'd326
; 
32'd20306: dataIn1 = 32'd328
; 
32'd20307: dataIn1 = 32'd333
; 
32'd20308: dataIn1 = 32'd362
; 
32'd20309: dataIn1 = 32'd375
; 
32'd20310: dataIn1 = 32'd389
; 
32'd20311: dataIn1 = 32'd407
; 
32'd20312: dataIn1 = 32'd412
; 
32'd20313: dataIn1 = 32'd420
; 
32'd20314: dataIn1 = 32'd427
; 
32'd20315: dataIn1 = 32'd481
; 
32'd20316: dataIn1 = 32'd506
; 
32'd20317: dataIn1 = 32'd508
; 
32'd20318: dataIn1 = 32'd525
; 
32'd20319: dataIn1 = 32'd570
; 
32'd20320: dataIn1 = 32'd578
; 
32'd20321: dataIn1 = 32'd610
; 
32'd20322: dataIn1 = 32'd617
; 
32'd20323: dataIn1 = 32'd716
; 
32'd20324: dataIn1 = 32'd718
; 
32'd20325: dataIn1 = 32'd726
; 
32'd20326: dataIn1 = 32'd769
; 
32'd20327: dataIn1 = 32'd399
; 
32'd20328: dataIn1 = 32'd402
; 
32'd20329: dataIn1 = 32'd403
; 
32'd20330: dataIn1 = 32'd409
; 
32'd20331: dataIn1 = 32'd420
; 
32'd20332: dataIn1 = 32'd432
; 
32'd20333: dataIn1 = 32'd448
; 
32'd20334: dataIn1 = 32'd471
; 
32'd20335: dataIn1 = 32'd509
; 
32'd20336: dataIn1 = 32'd512
; 
32'd20337: dataIn1 = 32'd516
; 
32'd20338: dataIn1 = 32'd553
; 
32'd20339: dataIn1 = 32'd557
; 
32'd20340: dataIn1 = 32'd564
; 
32'd20341: dataIn1 = 32'd582
; 
32'd20342: dataIn1 = 32'd592
; 
32'd20343: dataIn1 = 32'd598
; 
32'd20344: dataIn1 = 32'd620
; 
32'd20345: dataIn1 = 32'd630
; 
32'd20346: dataIn1 = 32'd644
; 
32'd20347: dataIn1 = 32'd668
; 
32'd20348: dataIn1 = 32'd670
; 
32'd20349: dataIn1 = 32'd700
; 
32'd20350: dataIn1 = 32'd743
; 
32'd20351: dataIn1 = 32'd746
; 
32'd20352: dataIn1 = 32'd754
; 
32'd20353: dataIn1 = 32'd782
; 
32'd20354: dataIn1 = 32'd786
; 
32'd20355: dataIn1 = 32'd791
; 
32'd20356: dataIn1 = 32'd798
; 
32'd20357: dataIn1 = 32'd323
; 
32'd20358: dataIn1 = 32'd340
; 
32'd20359: dataIn1 = 32'd380
; 
32'd20360: dataIn1 = 32'd388
; 
32'd20361: dataIn1 = 32'd401
; 
32'd20362: dataIn1 = 32'd423
; 
32'd20363: dataIn1 = 32'd437
; 
32'd20364: dataIn1 = 32'd460
; 
32'd20365: dataIn1 = 32'd475
; 
32'd20366: dataIn1 = 32'd481
; 
32'd20367: dataIn1 = 32'd485
; 
32'd20368: dataIn1 = 32'd487
; 
32'd20369: dataIn1 = 32'd492
; 
32'd20370: dataIn1 = 32'd496
; 
32'd20371: dataIn1 = 32'd550
; 
32'd20372: dataIn1 = 32'd555
; 
32'd20373: dataIn1 = 32'd557
; 
32'd20374: dataIn1 = 32'd605
; 
32'd20375: dataIn1 = 32'd606
; 
32'd20376: dataIn1 = 32'd646
; 
32'd20377: dataIn1 = 32'd647
; 
32'd20378: dataIn1 = 32'd653
; 
32'd20379: dataIn1 = 32'd664
; 
32'd20380: dataIn1 = 32'd676
; 
32'd20381: dataIn1 = 32'd692
; 
32'd20382: dataIn1 = 32'd755
; 
32'd20383: dataIn1 = 32'd756
; 
32'd20384: dataIn1 = 32'd773
; 
32'd20385: dataIn1 = 32'd774
; 
32'd20386: dataIn1 = 32'd778
; 
32'd20387: dataIn1 = 32'd784
; 
32'd20388: dataIn1 = 32'd799
; 
32'd20389: dataIn1 = 32'd331
; 
32'd20390: dataIn1 = 32'd332
; 
32'd20391: dataIn1 = 32'd391
; 
32'd20392: dataIn1 = 32'd414
; 
32'd20393: dataIn1 = 32'd439
; 
32'd20394: dataIn1 = 32'd477
; 
32'd20395: dataIn1 = 32'd480
; 
32'd20396: dataIn1 = 32'd486
; 
32'd20397: dataIn1 = 32'd487
; 
32'd20398: dataIn1 = 32'd517
; 
32'd20399: dataIn1 = 32'd520
; 
32'd20400: dataIn1 = 32'd526
; 
32'd20401: dataIn1 = 32'd534
; 
32'd20402: dataIn1 = 32'd555
; 
32'd20403: dataIn1 = 32'd559
; 
32'd20404: dataIn1 = 32'd564
; 
32'd20405: dataIn1 = 32'd571
; 
32'd20406: dataIn1 = 32'd589
; 
32'd20407: dataIn1 = 32'd611
; 
32'd20408: dataIn1 = 32'd620
; 
32'd20409: dataIn1 = 32'd643
; 
32'd20410: dataIn1 = 32'd654
; 
32'd20411: dataIn1 = 32'd687
; 
32'd20412: dataIn1 = 32'd701
; 
32'd20413: dataIn1 = 32'd709
; 
32'd20414: dataIn1 = 32'd739
; 
32'd20415: dataIn1 = 32'd755
; 
32'd20416: dataIn1 = 32'd757
; 
32'd20417: dataIn1 = 32'd794
; 
32'd20418: dataIn1 = 32'd333
; 
32'd20419: dataIn1 = 32'd362
; 
32'd20420: dataIn1 = 32'd381
; 
32'd20421: dataIn1 = 32'd491
; 
32'd20422: dataIn1 = 32'd497
; 
32'd20423: dataIn1 = 32'd498
; 
32'd20424: dataIn1 = 32'd514
; 
32'd20425: dataIn1 = 32'd524
; 
32'd20426: dataIn1 = 32'd553
; 
32'd20427: dataIn1 = 32'd561
; 
32'd20428: dataIn1 = 32'd587
; 
32'd20429: dataIn1 = 32'd600
; 
32'd20430: dataIn1 = 32'd616
; 
32'd20431: dataIn1 = 32'd634
; 
32'd20432: dataIn1 = 32'd653
; 
32'd20433: dataIn1 = 32'd673
; 
32'd20434: dataIn1 = 32'd704
; 
32'd20435: dataIn1 = 32'd723
; 
32'd20436: dataIn1 = 32'd732
; 
32'd20437: dataIn1 = 32'd741
; 
32'd20438: dataIn1 = 32'd746
; 
32'd20439: dataIn1 = 32'd767
; 
32'd20440: dataIn1 = 32'd774
; 
32'd20441: dataIn1 = 32'd778
; 
32'd20442: dataIn1 = 32'd795
; 
32'd20443: dataIn1 = 32'd352
; 
32'd20444: dataIn1 = 32'd366
; 
32'd20445: dataIn1 = 32'd368
; 
32'd20446: dataIn1 = 32'd369
; 
32'd20447: dataIn1 = 32'd414
; 
32'd20448: dataIn1 = 32'd427
; 
32'd20449: dataIn1 = 32'd508
; 
32'd20450: dataIn1 = 32'd510
; 
32'd20451: dataIn1 = 32'd523
; 
32'd20452: dataIn1 = 32'd525
; 
32'd20453: dataIn1 = 32'd526
; 
32'd20454: dataIn1 = 32'd557
; 
32'd20455: dataIn1 = 32'd569
; 
32'd20456: dataIn1 = 32'd594
; 
32'd20457: dataIn1 = 32'd599
; 
32'd20458: dataIn1 = 32'd611
; 
32'd20459: dataIn1 = 32'd613
; 
32'd20460: dataIn1 = 32'd639
; 
32'd20461: dataIn1 = 32'd646
; 
32'd20462: dataIn1 = 32'd677
; 
32'd20463: dataIn1 = 32'd685
; 
32'd20464: dataIn1 = 32'd698
; 
32'd20465: dataIn1 = 32'd709
; 
32'd20466: dataIn1 = 32'd710
; 
32'd20467: dataIn1 = 32'd720
; 
32'd20468: dataIn1 = 32'd750
; 
32'd20469: dataIn1 = 32'd767
; 
32'd20470: dataIn1 = 32'd330
; 
32'd20471: dataIn1 = 32'd365
; 
32'd20472: dataIn1 = 32'd416
; 
32'd20473: dataIn1 = 32'd433
; 
32'd20474: dataIn1 = 32'd463
; 
32'd20475: dataIn1 = 32'd466
; 
32'd20476: dataIn1 = 32'd499
; 
32'd20477: dataIn1 = 32'd506
; 
32'd20478: dataIn1 = 32'd536
; 
32'd20479: dataIn1 = 32'd539
; 
32'd20480: dataIn1 = 32'd554
; 
32'd20481: dataIn1 = 32'd567
; 
32'd20482: dataIn1 = 32'd629
; 
32'd20483: dataIn1 = 32'd645
; 
32'd20484: dataIn1 = 32'd653
; 
32'd20485: dataIn1 = 32'd654
; 
32'd20486: dataIn1 = 32'd692
; 
32'd20487: dataIn1 = 32'd712
; 
32'd20488: dataIn1 = 32'd719
; 
32'd20489: dataIn1 = 32'd721
; 
32'd20490: dataIn1 = 32'd748
; 
32'd20491: dataIn1 = 32'd332
; 
32'd20492: dataIn1 = 32'd341
; 
32'd20493: dataIn1 = 32'd375
; 
32'd20494: dataIn1 = 32'd384
; 
32'd20495: dataIn1 = 32'd403
; 
32'd20496: dataIn1 = 32'd426
; 
32'd20497: dataIn1 = 32'd428
; 
32'd20498: dataIn1 = 32'd462
; 
32'd20499: dataIn1 = 32'd472
; 
32'd20500: dataIn1 = 32'd481
; 
32'd20501: dataIn1 = 32'd491
; 
32'd20502: dataIn1 = 32'd501
; 
32'd20503: dataIn1 = 32'd549
; 
32'd20504: dataIn1 = 32'd554
; 
32'd20505: dataIn1 = 32'd564
; 
32'd20506: dataIn1 = 32'd572
; 
32'd20507: dataIn1 = 32'd592
; 
32'd20508: dataIn1 = 32'd597
; 
32'd20509: dataIn1 = 32'd604
; 
32'd20510: dataIn1 = 32'd613
; 
32'd20511: dataIn1 = 32'd619
; 
32'd20512: dataIn1 = 32'd633
; 
32'd20513: dataIn1 = 32'd643
; 
32'd20514: dataIn1 = 32'd663
; 
32'd20515: dataIn1 = 32'd674
; 
32'd20516: dataIn1 = 32'd676
; 
32'd20517: dataIn1 = 32'd707
; 
32'd20518: dataIn1 = 32'd711
; 
32'd20519: dataIn1 = 32'd713
; 
32'd20520: dataIn1 = 32'd730
; 
32'd20521: dataIn1 = 32'd732
; 
32'd20522: dataIn1 = 32'd761
; 
32'd20523: dataIn1 = 32'd766
; 
32'd20524: dataIn1 = 32'd767
; 
32'd20525: dataIn1 = 32'd783
; 
32'd20526: dataIn1 = 32'd793
; 
32'd20527: dataIn1 = 32'd338
; 
32'd20528: dataIn1 = 32'd345
; 
32'd20529: dataIn1 = 32'd377
; 
32'd20530: dataIn1 = 32'd391
; 
32'd20531: dataIn1 = 32'd396
; 
32'd20532: dataIn1 = 32'd415
; 
32'd20533: dataIn1 = 32'd418
; 
32'd20534: dataIn1 = 32'd423
; 
32'd20535: dataIn1 = 32'd426
; 
32'd20536: dataIn1 = 32'd427
; 
32'd20537: dataIn1 = 32'd428
; 
32'd20538: dataIn1 = 32'd432
; 
32'd20539: dataIn1 = 32'd450
; 
32'd20540: dataIn1 = 32'd454
; 
32'd20541: dataIn1 = 32'd554
; 
32'd20542: dataIn1 = 32'd575
; 
32'd20543: dataIn1 = 32'd594
; 
32'd20544: dataIn1 = 32'd598
; 
32'd20545: dataIn1 = 32'd602
; 
32'd20546: dataIn1 = 32'd613
; 
32'd20547: dataIn1 = 32'd625
; 
32'd20548: dataIn1 = 32'd628
; 
32'd20549: dataIn1 = 32'd644
; 
32'd20550: dataIn1 = 32'd647
; 
32'd20551: dataIn1 = 32'd651
; 
32'd20552: dataIn1 = 32'd691
; 
32'd20553: dataIn1 = 32'd695
; 
32'd20554: dataIn1 = 32'd700
; 
32'd20555: dataIn1 = 32'd702
; 
32'd20556: dataIn1 = 32'd713
; 
32'd20557: dataIn1 = 32'd717
; 
32'd20558: dataIn1 = 32'd719
; 
32'd20559: dataIn1 = 32'd748
; 
32'd20560: dataIn1 = 32'd762
; 
32'd20561: dataIn1 = 32'd768
; 
32'd20562: dataIn1 = 32'd330
; 
32'd20563: dataIn1 = 32'd352
; 
32'd20564: dataIn1 = 32'd376
; 
32'd20565: dataIn1 = 32'd387
; 
32'd20566: dataIn1 = 32'd397
; 
32'd20567: dataIn1 = 32'd400
; 
32'd20568: dataIn1 = 32'd414
; 
32'd20569: dataIn1 = 32'd438
; 
32'd20570: dataIn1 = 32'd468
; 
32'd20571: dataIn1 = 32'd493
; 
32'd20572: dataIn1 = 32'd507
; 
32'd20573: dataIn1 = 32'd528
; 
32'd20574: dataIn1 = 32'd550
; 
32'd20575: dataIn1 = 32'd589
; 
32'd20576: dataIn1 = 32'd627
; 
32'd20577: dataIn1 = 32'd657
; 
32'd20578: dataIn1 = 32'd666
; 
32'd20579: dataIn1 = 32'd686
; 
32'd20580: dataIn1 = 32'd690
; 
32'd20581: dataIn1 = 32'd707
; 
32'd20582: dataIn1 = 32'd708
; 
32'd20583: dataIn1 = 32'd709
; 
32'd20584: dataIn1 = 32'd757
; 
32'd20585: dataIn1 = 32'd763
; 
32'd20586: dataIn1 = 32'd797
; 
32'd20587: dataIn1 = 32'd339
; 
32'd20588: dataIn1 = 32'd341
; 
32'd20589: dataIn1 = 32'd419
; 
32'd20590: dataIn1 = 32'd454
; 
32'd20591: dataIn1 = 32'd456
; 
32'd20592: dataIn1 = 32'd462
; 
32'd20593: dataIn1 = 32'd470
; 
32'd20594: dataIn1 = 32'd505
; 
32'd20595: dataIn1 = 32'd508
; 
32'd20596: dataIn1 = 32'd517
; 
32'd20597: dataIn1 = 32'd518
; 
32'd20598: dataIn1 = 32'd531
; 
32'd20599: dataIn1 = 32'd554
; 
32'd20600: dataIn1 = 32'd592
; 
32'd20601: dataIn1 = 32'd613
; 
32'd20602: dataIn1 = 32'd629
; 
32'd20603: dataIn1 = 32'd634
; 
32'd20604: dataIn1 = 32'd637
; 
32'd20605: dataIn1 = 32'd655
; 
32'd20606: dataIn1 = 32'd660
; 
32'd20607: dataIn1 = 32'd684
; 
32'd20608: dataIn1 = 32'd685
; 
32'd20609: dataIn1 = 32'd687
; 
32'd20610: dataIn1 = 32'd707
; 
32'd20611: dataIn1 = 32'd738
; 
32'd20612: dataIn1 = 32'd770
; 
32'd20613: dataIn1 = 32'd787
; 
32'd20614: dataIn1 = 32'd797
; 
32'd20615: dataIn1 = 32'd338
; 
32'd20616: dataIn1 = 32'd343
; 
32'd20617: dataIn1 = 32'd364
; 
32'd20618: dataIn1 = 32'd378
; 
32'd20619: dataIn1 = 32'd381
; 
32'd20620: dataIn1 = 32'd409
; 
32'd20621: dataIn1 = 32'd411
; 
32'd20622: dataIn1 = 32'd426
; 
32'd20623: dataIn1 = 32'd435
; 
32'd20624: dataIn1 = 32'd436
; 
32'd20625: dataIn1 = 32'd444
; 
32'd20626: dataIn1 = 32'd468
; 
32'd20627: dataIn1 = 32'd471
; 
32'd20628: dataIn1 = 32'd475
; 
32'd20629: dataIn1 = 32'd484
; 
32'd20630: dataIn1 = 32'd532
; 
32'd20631: dataIn1 = 32'd576
; 
32'd20632: dataIn1 = 32'd620
; 
32'd20633: dataIn1 = 32'd634
; 
32'd20634: dataIn1 = 32'd639
; 
32'd20635: dataIn1 = 32'd660
; 
32'd20636: dataIn1 = 32'd669
; 
32'd20637: dataIn1 = 32'd682
; 
32'd20638: dataIn1 = 32'd686
; 
32'd20639: dataIn1 = 32'd688
; 
32'd20640: dataIn1 = 32'd710
; 
32'd20641: dataIn1 = 32'd713
; 
32'd20642: dataIn1 = 32'd718
; 
32'd20643: dataIn1 = 32'd762
; 
32'd20644: dataIn1 = 32'd770
; 
32'd20645: dataIn1 = 32'd788
; 
32'd20646: dataIn1 = 32'd789
; 
32'd20647: dataIn1 = 32'd793
; 
32'd20648: dataIn1 = 32'd800
; 
32'd20649: dataIn1 = 32'd342
; 
32'd20650: dataIn1 = 32'd349
; 
32'd20651: dataIn1 = 32'd367
; 
32'd20652: dataIn1 = 32'd389
; 
32'd20653: dataIn1 = 32'd397
; 
32'd20654: dataIn1 = 32'd412
; 
32'd20655: dataIn1 = 32'd426
; 
32'd20656: dataIn1 = 32'd470
; 
32'd20657: dataIn1 = 32'd500
; 
32'd20658: dataIn1 = 32'd518
; 
32'd20659: dataIn1 = 32'd554
; 
32'd20660: dataIn1 = 32'd582
; 
32'd20661: dataIn1 = 32'd601
; 
32'd20662: dataIn1 = 32'd618
; 
32'd20663: dataIn1 = 32'd619
; 
32'd20664: dataIn1 = 32'd637
; 
32'd20665: dataIn1 = 32'd660
; 
32'd20666: dataIn1 = 32'd664
; 
32'd20667: dataIn1 = 32'd681
; 
32'd20668: dataIn1 = 32'd694
; 
32'd20669: dataIn1 = 32'd716
; 
32'd20670: dataIn1 = 32'd745
; 
32'd20671: dataIn1 = 32'd746
; 
32'd20672: dataIn1 = 32'd763
; 
32'd20673: dataIn1 = 32'd779
; 
32'd20674: dataIn1 = 32'd338
; 
32'd20675: dataIn1 = 32'd394
; 
32'd20676: dataIn1 = 32'd396
; 
32'd20677: dataIn1 = 32'd405
; 
32'd20678: dataIn1 = 32'd419
; 
32'd20679: dataIn1 = 32'd430
; 
32'd20680: dataIn1 = 32'd456
; 
32'd20681: dataIn1 = 32'd511
; 
32'd20682: dataIn1 = 32'd534
; 
32'd20683: dataIn1 = 32'd554
; 
32'd20684: dataIn1 = 32'd568
; 
32'd20685: dataIn1 = 32'd569
; 
32'd20686: dataIn1 = 32'd594
; 
32'd20687: dataIn1 = 32'd622
; 
32'd20688: dataIn1 = 32'd656
; 
32'd20689: dataIn1 = 32'd672
; 
32'd20690: dataIn1 = 32'd698
; 
32'd20691: dataIn1 = 32'd704
; 
32'd20692: dataIn1 = 32'd706
; 
32'd20693: dataIn1 = 32'd709
; 
32'd20694: dataIn1 = 32'd743
; 
32'd20695: dataIn1 = 32'd746
; 
32'd20696: dataIn1 = 32'd752
; 
32'd20697: dataIn1 = 32'd786
; 
32'd20698: dataIn1 = 32'd789
; 
32'd20699: dataIn1 = 32'd344
; 
32'd20700: dataIn1 = 32'd359
; 
32'd20701: dataIn1 = 32'd373
; 
32'd20702: dataIn1 = 32'd376
; 
32'd20703: dataIn1 = 32'd377
; 
32'd20704: dataIn1 = 32'd399
; 
32'd20705: dataIn1 = 32'd406
; 
32'd20706: dataIn1 = 32'd420
; 
32'd20707: dataIn1 = 32'd441
; 
32'd20708: dataIn1 = 32'd448
; 
32'd20709: dataIn1 = 32'd496
; 
32'd20710: dataIn1 = 32'd500
; 
32'd20711: dataIn1 = 32'd503
; 
32'd20712: dataIn1 = 32'd518
; 
32'd20713: dataIn1 = 32'd532
; 
32'd20714: dataIn1 = 32'd549
; 
32'd20715: dataIn1 = 32'd564
; 
32'd20716: dataIn1 = 32'd572
; 
32'd20717: dataIn1 = 32'd593
; 
32'd20718: dataIn1 = 32'd598
; 
32'd20719: dataIn1 = 32'd632
; 
32'd20720: dataIn1 = 32'd676
; 
32'd20721: dataIn1 = 32'd682
; 
32'd20722: dataIn1 = 32'd690
; 
32'd20723: dataIn1 = 32'd694
; 
32'd20724: dataIn1 = 32'd710
; 
32'd20725: dataIn1 = 32'd711
; 
32'd20726: dataIn1 = 32'd728
; 
32'd20727: dataIn1 = 32'd729
; 
32'd20728: dataIn1 = 32'd765
; 
32'd20729: dataIn1 = 32'd796
; 
32'd20730: dataIn1 = 32'd365
; 
32'd20731: dataIn1 = 32'd386
; 
32'd20732: dataIn1 = 32'd390
; 
32'd20733: dataIn1 = 32'd394
; 
32'd20734: dataIn1 = 32'd442
; 
32'd20735: dataIn1 = 32'd448
; 
32'd20736: dataIn1 = 32'd478
; 
32'd20737: dataIn1 = 32'd502
; 
32'd20738: dataIn1 = 32'd527
; 
32'd20739: dataIn1 = 32'd534
; 
32'd20740: dataIn1 = 32'd545
; 
32'd20741: dataIn1 = 32'd554
; 
32'd20742: dataIn1 = 32'd556
; 
32'd20743: dataIn1 = 32'd583
; 
32'd20744: dataIn1 = 32'd595
; 
32'd20745: dataIn1 = 32'd643
; 
32'd20746: dataIn1 = 32'd654
; 
32'd20747: dataIn1 = 32'd667
; 
32'd20748: dataIn1 = 32'd672
; 
32'd20749: dataIn1 = 32'd690
; 
32'd20750: dataIn1 = 32'd702
; 
32'd20751: dataIn1 = 32'd706
; 
32'd20752: dataIn1 = 32'd721
; 
32'd20753: dataIn1 = 32'd751
; 
32'd20754: dataIn1 = 32'd782
; 
32'd20755: dataIn1 = 32'd343
; 
32'd20756: dataIn1 = 32'd378
; 
32'd20757: dataIn1 = 32'd391
; 
32'd20758: dataIn1 = 32'd399
; 
32'd20759: dataIn1 = 32'd407
; 
32'd20760: dataIn1 = 32'd422
; 
32'd20761: dataIn1 = 32'd424
; 
32'd20762: dataIn1 = 32'd450
; 
32'd20763: dataIn1 = 32'd520
; 
32'd20764: dataIn1 = 32'd530
; 
32'd20765: dataIn1 = 32'd563
; 
32'd20766: dataIn1 = 32'd568
; 
32'd20767: dataIn1 = 32'd608
; 
32'd20768: dataIn1 = 32'd623
; 
32'd20769: dataIn1 = 32'd665
; 
32'd20770: dataIn1 = 32'd676
; 
32'd20771: dataIn1 = 32'd684
; 
32'd20772: dataIn1 = 32'd756
; 
32'd20773: dataIn1 = 32'd781
; 
32'd20774: dataIn1 = 32'd798
; 
32'd20775: dataIn1 = 32'd356
; 
32'd20776: dataIn1 = 32'd367
; 
32'd20777: dataIn1 = 32'd389
; 
32'd20778: dataIn1 = 32'd400
; 
32'd20779: dataIn1 = 32'd418
; 
32'd20780: dataIn1 = 32'd444
; 
32'd20781: dataIn1 = 32'd466
; 
32'd20782: dataIn1 = 32'd473
; 
32'd20783: dataIn1 = 32'd486
; 
32'd20784: dataIn1 = 32'd507
; 
32'd20785: dataIn1 = 32'd518
; 
32'd20786: dataIn1 = 32'd523
; 
32'd20787: dataIn1 = 32'd586
; 
32'd20788: dataIn1 = 32'd613
; 
32'd20789: dataIn1 = 32'd616
; 
32'd20790: dataIn1 = 32'd626
; 
32'd20791: dataIn1 = 32'd633
; 
32'd20792: dataIn1 = 32'd635
; 
32'd20793: dataIn1 = 32'd637
; 
32'd20794: dataIn1 = 32'd638
; 
32'd20795: dataIn1 = 32'd677
; 
32'd20796: dataIn1 = 32'd678
; 
32'd20797: dataIn1 = 32'd698
; 
32'd20798: dataIn1 = 32'd704
; 
32'd20799: dataIn1 = 32'd799
; 
32'd20800: dataIn1 = 32'd800
; 
32'd20801: dataIn1 = 32'd338
; 
32'd20802: dataIn1 = 32'd340
; 
32'd20803: dataIn1 = 32'd376
; 
32'd20804: dataIn1 = 32'd430
; 
32'd20805: dataIn1 = 32'd442
; 
32'd20806: dataIn1 = 32'd451
; 
32'd20807: dataIn1 = 32'd462
; 
32'd20808: dataIn1 = 32'd483
; 
32'd20809: dataIn1 = 32'd576
; 
32'd20810: dataIn1 = 32'd602
; 
32'd20811: dataIn1 = 32'd603
; 
32'd20812: dataIn1 = 32'd614
; 
32'd20813: dataIn1 = 32'd618
; 
32'd20814: dataIn1 = 32'd619
; 
32'd20815: dataIn1 = 32'd641
; 
32'd20816: dataIn1 = 32'd647
; 
32'd20817: dataIn1 = 32'd654
; 
32'd20818: dataIn1 = 32'd663
; 
32'd20819: dataIn1 = 32'd682
; 
32'd20820: dataIn1 = 32'd684
; 
32'd20821: dataIn1 = 32'd691
; 
32'd20822: dataIn1 = 32'd721
; 
32'd20823: dataIn1 = 32'd772
; 
32'd20824: dataIn1 = 32'd791
; 
32'd20825: dataIn1 = 32'd342
; 
32'd20826: dataIn1 = 32'd382
; 
32'd20827: dataIn1 = 32'd396
; 
32'd20828: dataIn1 = 32'd414
; 
32'd20829: dataIn1 = 32'd418
; 
32'd20830: dataIn1 = 32'd422
; 
32'd20831: dataIn1 = 32'd433
; 
32'd20832: dataIn1 = 32'd497
; 
32'd20833: dataIn1 = 32'd532
; 
32'd20834: dataIn1 = 32'd559
; 
32'd20835: dataIn1 = 32'd602
; 
32'd20836: dataIn1 = 32'd615
; 
32'd20837: dataIn1 = 32'd625
; 
32'd20838: dataIn1 = 32'd631
; 
32'd20839: dataIn1 = 32'd646
; 
32'd20840: dataIn1 = 32'd665
; 
32'd20841: dataIn1 = 32'd681
; 
32'd20842: dataIn1 = 32'd688
; 
32'd20843: dataIn1 = 32'd692
; 
32'd20844: dataIn1 = 32'd694
; 
32'd20845: dataIn1 = 32'd707
; 
32'd20846: dataIn1 = 32'd716
; 
32'd20847: dataIn1 = 32'd735
; 
32'd20848: dataIn1 = 32'd770
; 
32'd20849: dataIn1 = 32'd799
; 
32'd20850: dataIn1 = 32'd345
; 
32'd20851: dataIn1 = 32'd353
; 
32'd20852: dataIn1 = 32'd373
; 
32'd20853: dataIn1 = 32'd380
; 
32'd20854: dataIn1 = 32'd419
; 
32'd20855: dataIn1 = 32'd492
; 
32'd20856: dataIn1 = 32'd494
; 
32'd20857: dataIn1 = 32'd504
; 
32'd20858: dataIn1 = 32'd509
; 
32'd20859: dataIn1 = 32'd538
; 
32'd20860: dataIn1 = 32'd545
; 
32'd20861: dataIn1 = 32'd554
; 
32'd20862: dataIn1 = 32'd562
; 
32'd20863: dataIn1 = 32'd575
; 
32'd20864: dataIn1 = 32'd577
; 
32'd20865: dataIn1 = 32'd622
; 
32'd20866: dataIn1 = 32'd623
; 
32'd20867: dataIn1 = 32'd633
; 
32'd20868: dataIn1 = 32'd634
; 
32'd20869: dataIn1 = 32'd655
; 
32'd20870: dataIn1 = 32'd660
; 
32'd20871: dataIn1 = 32'd683
; 
32'd20872: dataIn1 = 32'd687
; 
32'd20873: dataIn1 = 32'd745
; 
32'd20874: dataIn1 = 32'd746
; 
32'd20875: dataIn1 = 32'd766
; 
32'd20876: dataIn1 = 32'd782
; 
32'd20877: dataIn1 = 32'd791
; 
32'd20878: dataIn1 = 32'd345
; 
32'd20879: dataIn1 = 32'd371
; 
32'd20880: dataIn1 = 32'd394
; 
32'd20881: dataIn1 = 32'd396
; 
32'd20882: dataIn1 = 32'd400
; 
32'd20883: dataIn1 = 32'd420
; 
32'd20884: dataIn1 = 32'd453
; 
32'd20885: dataIn1 = 32'd468
; 
32'd20886: dataIn1 = 32'd471
; 
32'd20887: dataIn1 = 32'd474
; 
32'd20888: dataIn1 = 32'd523
; 
32'd20889: dataIn1 = 32'd556
; 
32'd20890: dataIn1 = 32'd562
; 
32'd20891: dataIn1 = 32'd586
; 
32'd20892: dataIn1 = 32'd602
; 
32'd20893: dataIn1 = 32'd612
; 
32'd20894: dataIn1 = 32'd617
; 
32'd20895: dataIn1 = 32'd643
; 
32'd20896: dataIn1 = 32'd654
; 
32'd20897: dataIn1 = 32'd661
; 
32'd20898: dataIn1 = 32'd662
; 
32'd20899: dataIn1 = 32'd674
; 
32'd20900: dataIn1 = 32'd713
; 
32'd20901: dataIn1 = 32'd744
; 
32'd20902: dataIn1 = 32'd771
; 
32'd20903: dataIn1 = 32'd780
; 
32'd20904: dataIn1 = 32'd782
; 
32'd20905: dataIn1 = 32'd785
; 
32'd20906: dataIn1 = 32'd794
; 
32'd20907: dataIn1 = 32'd796
; 
32'd20908: dataIn1 = 32'd350
; 
32'd20909: dataIn1 = 32'd410
; 
32'd20910: dataIn1 = 32'd413
; 
32'd20911: dataIn1 = 32'd422
; 
32'd20912: dataIn1 = 32'd429
; 
32'd20913: dataIn1 = 32'd431
; 
32'd20914: dataIn1 = 32'd444
; 
32'd20915: dataIn1 = 32'd448
; 
32'd20916: dataIn1 = 32'd473
; 
32'd20917: dataIn1 = 32'd476
; 
32'd20918: dataIn1 = 32'd483
; 
32'd20919: dataIn1 = 32'd484
; 
32'd20920: dataIn1 = 32'd490
; 
32'd20921: dataIn1 = 32'd491
; 
32'd20922: dataIn1 = 32'd551
; 
32'd20923: dataIn1 = 32'd630
; 
32'd20924: dataIn1 = 32'd664
; 
32'd20925: dataIn1 = 32'd665
; 
32'd20926: dataIn1 = 32'd666
; 
32'd20927: dataIn1 = 32'd715
; 
32'd20928: dataIn1 = 32'd749
; 
32'd20929: dataIn1 = 32'd756
; 
32'd20930: dataIn1 = 32'd763
; 
32'd20931: dataIn1 = 32'd787
; 
32'd20932: dataIn1 = 32'd798
; 
32'd20933: dataIn1 = 32'd362
; 
32'd20934: dataIn1 = 32'd365
; 
32'd20935: dataIn1 = 32'd366
; 
32'd20936: dataIn1 = 32'd373
; 
32'd20937: dataIn1 = 32'd375
; 
32'd20938: dataIn1 = 32'd467
; 
32'd20939: dataIn1 = 32'd469
; 
32'd20940: dataIn1 = 32'd478
; 
32'd20941: dataIn1 = 32'd483
; 
32'd20942: dataIn1 = 32'd501
; 
32'd20943: dataIn1 = 32'd548
; 
32'd20944: dataIn1 = 32'd572
; 
32'd20945: dataIn1 = 32'd577
; 
32'd20946: dataIn1 = 32'd579
; 
32'd20947: dataIn1 = 32'd602
; 
32'd20948: dataIn1 = 32'd629
; 
32'd20949: dataIn1 = 32'd635
; 
32'd20950: dataIn1 = 32'd640
; 
32'd20951: dataIn1 = 32'd643
; 
32'd20952: dataIn1 = 32'd698
; 
32'd20953: dataIn1 = 32'd723
; 
32'd20954: dataIn1 = 32'd759
; 
32'd20955: dataIn1 = 32'd785
; 
32'd20956: dataIn1 = 32'd344
; 
32'd20957: dataIn1 = 32'd371
; 
32'd20958: dataIn1 = 32'd374
; 
32'd20959: dataIn1 = 32'd377
; 
32'd20960: dataIn1 = 32'd384
; 
32'd20961: dataIn1 = 32'd439
; 
32'd20962: dataIn1 = 32'd444
; 
32'd20963: dataIn1 = 32'd501
; 
32'd20964: dataIn1 = 32'd505
; 
32'd20965: dataIn1 = 32'd517
; 
32'd20966: dataIn1 = 32'd526
; 
32'd20967: dataIn1 = 32'd582
; 
32'd20968: dataIn1 = 32'd610
; 
32'd20969: dataIn1 = 32'd626
; 
32'd20970: dataIn1 = 32'd643
; 
32'd20971: dataIn1 = 32'd649
; 
32'd20972: dataIn1 = 32'd660
; 
32'd20973: dataIn1 = 32'd661
; 
32'd20974: dataIn1 = 32'd700
; 
32'd20975: dataIn1 = 32'd701
; 
32'd20976: dataIn1 = 32'd720
; 
32'd20977: dataIn1 = 32'd725
; 
32'd20978: dataIn1 = 32'd747
; 
32'd20979: dataIn1 = 32'd751
; 
32'd20980: dataIn1 = 32'd770
; 
32'd20981: dataIn1 = 32'd797
; 
32'd20982: dataIn1 = 32'd362
; 
32'd20983: dataIn1 = 32'd378
; 
32'd20984: dataIn1 = 32'd380
; 
32'd20985: dataIn1 = 32'd383
; 
32'd20986: dataIn1 = 32'd390
; 
32'd20987: dataIn1 = 32'd428
; 
32'd20988: dataIn1 = 32'd515
; 
32'd20989: dataIn1 = 32'd543
; 
32'd20990: dataIn1 = 32'd557
; 
32'd20991: dataIn1 = 32'd561
; 
32'd20992: dataIn1 = 32'd567
; 
32'd20993: dataIn1 = 32'd586
; 
32'd20994: dataIn1 = 32'd609
; 
32'd20995: dataIn1 = 32'd635
; 
32'd20996: dataIn1 = 32'd670
; 
32'd20997: dataIn1 = 32'd673
; 
32'd20998: dataIn1 = 32'd676
; 
32'd20999: dataIn1 = 32'd750
; 
32'd21000: dataIn1 = 32'd780
; 
32'd21001: dataIn1 = 32'd784
; 
32'd21002: dataIn1 = 32'd346
; 
32'd21003: dataIn1 = 32'd348
; 
32'd21004: dataIn1 = 32'd375
; 
32'd21005: dataIn1 = 32'd377
; 
32'd21006: dataIn1 = 32'd388
; 
32'd21007: dataIn1 = 32'd398
; 
32'd21008: dataIn1 = 32'd400
; 
32'd21009: dataIn1 = 32'd448
; 
32'd21010: dataIn1 = 32'd472
; 
32'd21011: dataIn1 = 32'd488
; 
32'd21012: dataIn1 = 32'd511
; 
32'd21013: dataIn1 = 32'd513
; 
32'd21014: dataIn1 = 32'd521
; 
32'd21015: dataIn1 = 32'd539
; 
32'd21016: dataIn1 = 32'd558
; 
32'd21017: dataIn1 = 32'd566
; 
32'd21018: dataIn1 = 32'd573
; 
32'd21019: dataIn1 = 32'd595
; 
32'd21020: dataIn1 = 32'd605
; 
32'd21021: dataIn1 = 32'd613
; 
32'd21022: dataIn1 = 32'd634
; 
32'd21023: dataIn1 = 32'd647
; 
32'd21024: dataIn1 = 32'd656
; 
32'd21025: dataIn1 = 32'd665
; 
32'd21026: dataIn1 = 32'd670
; 
32'd21027: dataIn1 = 32'd683
; 
32'd21028: dataIn1 = 32'd704
; 
32'd21029: dataIn1 = 32'd712
; 
32'd21030: dataIn1 = 32'd716
; 
32'd21031: dataIn1 = 32'd720
; 
32'd21032: dataIn1 = 32'd728
; 
32'd21033: dataIn1 = 32'd744
; 
32'd21034: dataIn1 = 32'd357
; 
32'd21035: dataIn1 = 32'd371
; 
32'd21036: dataIn1 = 32'd374
; 
32'd21037: dataIn1 = 32'd379
; 
32'd21038: dataIn1 = 32'd380
; 
32'd21039: dataIn1 = 32'd395
; 
32'd21040: dataIn1 = 32'd401
; 
32'd21041: dataIn1 = 32'd410
; 
32'd21042: dataIn1 = 32'd421
; 
32'd21043: dataIn1 = 32'd423
; 
32'd21044: dataIn1 = 32'd424
; 
32'd21045: dataIn1 = 32'd433
; 
32'd21046: dataIn1 = 32'd454
; 
32'd21047: dataIn1 = 32'd470
; 
32'd21048: dataIn1 = 32'd477
; 
32'd21049: dataIn1 = 32'd503
; 
32'd21050: dataIn1 = 32'd505
; 
32'd21051: dataIn1 = 32'd536
; 
32'd21052: dataIn1 = 32'd576
; 
32'd21053: dataIn1 = 32'd584
; 
32'd21054: dataIn1 = 32'd606
; 
32'd21055: dataIn1 = 32'd611
; 
32'd21056: dataIn1 = 32'd648
; 
32'd21057: dataIn1 = 32'd656
; 
32'd21058: dataIn1 = 32'd701
; 
32'd21059: dataIn1 = 32'd704
; 
32'd21060: dataIn1 = 32'd707
; 
32'd21061: dataIn1 = 32'd723
; 
32'd21062: dataIn1 = 32'd727
; 
32'd21063: dataIn1 = 32'd728
; 
32'd21064: dataIn1 = 32'd744
; 
32'd21065: dataIn1 = 32'd765
; 
32'd21066: dataIn1 = 32'd775
; 
32'd21067: dataIn1 = 32'd779
; 
32'd21068: dataIn1 = 32'd793
; 
32'd21069: dataIn1 = 32'd796
; 
32'd21070: dataIn1 = 32'd364
; 
32'd21071: dataIn1 = 32'd373
; 
32'd21072: dataIn1 = 32'd394
; 
32'd21073: dataIn1 = 32'd404
; 
32'd21074: dataIn1 = 32'd415
; 
32'd21075: dataIn1 = 32'd423
; 
32'd21076: dataIn1 = 32'd429
; 
32'd21077: dataIn1 = 32'd437
; 
32'd21078: dataIn1 = 32'd453
; 
32'd21079: dataIn1 = 32'd460
; 
32'd21080: dataIn1 = 32'd515
; 
32'd21081: dataIn1 = 32'd538
; 
32'd21082: dataIn1 = 32'd580
; 
32'd21083: dataIn1 = 32'd581
; 
32'd21084: dataIn1 = 32'd583
; 
32'd21085: dataIn1 = 32'd596
; 
32'd21086: dataIn1 = 32'd606
; 
32'd21087: dataIn1 = 32'd646
; 
32'd21088: dataIn1 = 32'd655
; 
32'd21089: dataIn1 = 32'd670
; 
32'd21090: dataIn1 = 32'd688
; 
32'd21091: dataIn1 = 32'd706
; 
32'd21092: dataIn1 = 32'd720
; 
32'd21093: dataIn1 = 32'd767
; 
32'd21094: dataIn1 = 32'd779
; 
32'd21095: dataIn1 = 32'd798
; 
32'd21096: dataIn1 = 32'd402
; 
32'd21097: dataIn1 = 32'd404
; 
32'd21098: dataIn1 = 32'd416
; 
32'd21099: dataIn1 = 32'd417
; 
32'd21100: dataIn1 = 32'd427
; 
32'd21101: dataIn1 = 32'd440
; 
32'd21102: dataIn1 = 32'd482
; 
32'd21103: dataIn1 = 32'd493
; 
32'd21104: dataIn1 = 32'd515
; 
32'd21105: dataIn1 = 32'd540
; 
32'd21106: dataIn1 = 32'd554
; 
32'd21107: dataIn1 = 32'd559
; 
32'd21108: dataIn1 = 32'd564
; 
32'd21109: dataIn1 = 32'd568
; 
32'd21110: dataIn1 = 32'd590
; 
32'd21111: dataIn1 = 32'd605
; 
32'd21112: dataIn1 = 32'd609
; 
32'd21113: dataIn1 = 32'd647
; 
32'd21114: dataIn1 = 32'd669
; 
32'd21115: dataIn1 = 32'd683
; 
32'd21116: dataIn1 = 32'd689
; 
32'd21117: dataIn1 = 32'd701
; 
32'd21118: dataIn1 = 32'd710
; 
32'd21119: dataIn1 = 32'd723
; 
32'd21120: dataIn1 = 32'd728
; 
32'd21121: dataIn1 = 32'd748
; 
32'd21122: dataIn1 = 32'd799
; 
32'd21123: dataIn1 = 32'd357
; 
32'd21124: dataIn1 = 32'd374
; 
32'd21125: dataIn1 = 32'd403
; 
32'd21126: dataIn1 = 32'd416
; 
32'd21127: dataIn1 = 32'd425
; 
32'd21128: dataIn1 = 32'd429
; 
32'd21129: dataIn1 = 32'd435
; 
32'd21130: dataIn1 = 32'd444
; 
32'd21131: dataIn1 = 32'd450
; 
32'd21132: dataIn1 = 32'd466
; 
32'd21133: dataIn1 = 32'd478
; 
32'd21134: dataIn1 = 32'd491
; 
32'd21135: dataIn1 = 32'd511
; 
32'd21136: dataIn1 = 32'd527
; 
32'd21137: dataIn1 = 32'd542
; 
32'd21138: dataIn1 = 32'd552
; 
32'd21139: dataIn1 = 32'd561
; 
32'd21140: dataIn1 = 32'd581
; 
32'd21141: dataIn1 = 32'd596
; 
32'd21142: dataIn1 = 32'd631
; 
32'd21143: dataIn1 = 32'd686
; 
32'd21144: dataIn1 = 32'd719
; 
32'd21145: dataIn1 = 32'd721
; 
32'd21146: dataIn1 = 32'd726
; 
32'd21147: dataIn1 = 32'd767
; 
32'd21148: dataIn1 = 32'd781
; 
32'd21149: dataIn1 = 32'd796
; 
32'd21150: dataIn1 = 32'd361
; 
32'd21151: dataIn1 = 32'd382
; 
32'd21152: dataIn1 = 32'd399
; 
32'd21153: dataIn1 = 32'd401
; 
32'd21154: dataIn1 = 32'd419
; 
32'd21155: dataIn1 = 32'd429
; 
32'd21156: dataIn1 = 32'd446
; 
32'd21157: dataIn1 = 32'd508
; 
32'd21158: dataIn1 = 32'd516
; 
32'd21159: dataIn1 = 32'd545
; 
32'd21160: dataIn1 = 32'd548
; 
32'd21161: dataIn1 = 32'd559
; 
32'd21162: dataIn1 = 32'd580
; 
32'd21163: dataIn1 = 32'd615
; 
32'd21164: dataIn1 = 32'd617
; 
32'd21165: dataIn1 = 32'd620
; 
32'd21166: dataIn1 = 32'd638
; 
32'd21167: dataIn1 = 32'd668
; 
32'd21168: dataIn1 = 32'd672
; 
32'd21169: dataIn1 = 32'd708
; 
32'd21170: dataIn1 = 32'd730
; 
32'd21171: dataIn1 = 32'd758
; 
32'd21172: dataIn1 = 32'd353
; 
32'd21173: dataIn1 = 32'd369
; 
32'd21174: dataIn1 = 32'd379
; 
32'd21175: dataIn1 = 32'd399
; 
32'd21176: dataIn1 = 32'd414
; 
32'd21177: dataIn1 = 32'd427
; 
32'd21178: dataIn1 = 32'd442
; 
32'd21179: dataIn1 = 32'd465
; 
32'd21180: dataIn1 = 32'd485
; 
32'd21181: dataIn1 = 32'd499
; 
32'd21182: dataIn1 = 32'd523
; 
32'd21183: dataIn1 = 32'd568
; 
32'd21184: dataIn1 = 32'd575
; 
32'd21185: dataIn1 = 32'd585
; 
32'd21186: dataIn1 = 32'd607
; 
32'd21187: dataIn1 = 32'd615
; 
32'd21188: dataIn1 = 32'd672
; 
32'd21189: dataIn1 = 32'd702
; 
32'd21190: dataIn1 = 32'd707
; 
32'd21191: dataIn1 = 32'd715
; 
32'd21192: dataIn1 = 32'd780
; 
32'd21193: dataIn1 = 32'd354
; 
32'd21194: dataIn1 = 32'd393
; 
32'd21195: dataIn1 = 32'd457
; 
32'd21196: dataIn1 = 32'd477
; 
32'd21197: dataIn1 = 32'd510
; 
32'd21198: dataIn1 = 32'd521
; 
32'd21199: dataIn1 = 32'd532
; 
32'd21200: dataIn1 = 32'd537
; 
32'd21201: dataIn1 = 32'd557
; 
32'd21202: dataIn1 = 32'd563
; 
32'd21203: dataIn1 = 32'd588
; 
32'd21204: dataIn1 = 32'd598
; 
32'd21205: dataIn1 = 32'd610
; 
32'd21206: dataIn1 = 32'd615
; 
32'd21207: dataIn1 = 32'd644
; 
32'd21208: dataIn1 = 32'd674
; 
32'd21209: dataIn1 = 32'd688
; 
32'd21210: dataIn1 = 32'd800
; 
32'd21211: dataIn1 = 32'd356
; 
32'd21212: dataIn1 = 32'd367
; 
32'd21213: dataIn1 = 32'd417
; 
32'd21214: dataIn1 = 32'd425
; 
32'd21215: dataIn1 = 32'd437
; 
32'd21216: dataIn1 = 32'd442
; 
32'd21217: dataIn1 = 32'd456
; 
32'd21218: dataIn1 = 32'd464
; 
32'd21219: dataIn1 = 32'd489
; 
32'd21220: dataIn1 = 32'd491
; 
32'd21221: dataIn1 = 32'd493
; 
32'd21222: dataIn1 = 32'd513
; 
32'd21223: dataIn1 = 32'd546
; 
32'd21224: dataIn1 = 32'd552
; 
32'd21225: dataIn1 = 32'd561
; 
32'd21226: dataIn1 = 32'd567
; 
32'd21227: dataIn1 = 32'd606
; 
32'd21228: dataIn1 = 32'd612
; 
32'd21229: dataIn1 = 32'd615
; 
32'd21230: dataIn1 = 32'd624
; 
32'd21231: dataIn1 = 32'd653
; 
32'd21232: dataIn1 = 32'd669
; 
32'd21233: dataIn1 = 32'd672
; 
32'd21234: dataIn1 = 32'd694
; 
32'd21235: dataIn1 = 32'd712
; 
32'd21236: dataIn1 = 32'd728
; 
32'd21237: dataIn1 = 32'd760
; 
32'd21238: dataIn1 = 32'd766
; 
32'd21239: dataIn1 = 32'd771
; 
32'd21240: dataIn1 = 32'd779
; 
32'd21241: dataIn1 = 32'd784
; 
32'd21242: dataIn1 = 32'd355
; 
32'd21243: dataIn1 = 32'd372
; 
32'd21244: dataIn1 = 32'd424
; 
32'd21245: dataIn1 = 32'd431
; 
32'd21246: dataIn1 = 32'd448
; 
32'd21247: dataIn1 = 32'd474
; 
32'd21248: dataIn1 = 32'd512
; 
32'd21249: dataIn1 = 32'd523
; 
32'd21250: dataIn1 = 32'd546
; 
32'd21251: dataIn1 = 32'd568
; 
32'd21252: dataIn1 = 32'd603
; 
32'd21253: dataIn1 = 32'd611
; 
32'd21254: dataIn1 = 32'd616
; 
32'd21255: dataIn1 = 32'd619
; 
32'd21256: dataIn1 = 32'd626
; 
32'd21257: dataIn1 = 32'd657
; 
32'd21258: dataIn1 = 32'd659
; 
32'd21259: dataIn1 = 32'd698
; 
32'd21260: dataIn1 = 32'd699
; 
32'd21261: dataIn1 = 32'd710
; 
32'd21262: dataIn1 = 32'd731
; 
32'd21263: dataIn1 = 32'd756
; 
32'd21264: dataIn1 = 32'd770
; 
32'd21265: dataIn1 = 32'd368
; 
32'd21266: dataIn1 = 32'd370
; 
32'd21267: dataIn1 = 32'd389
; 
32'd21268: dataIn1 = 32'd391
; 
32'd21269: dataIn1 = 32'd410
; 
32'd21270: dataIn1 = 32'd413
; 
32'd21271: dataIn1 = 32'd419
; 
32'd21272: dataIn1 = 32'd423
; 
32'd21273: dataIn1 = 32'd425
; 
32'd21274: dataIn1 = 32'd441
; 
32'd21275: dataIn1 = 32'd460
; 
32'd21276: dataIn1 = 32'd513
; 
32'd21277: dataIn1 = 32'd515
; 
32'd21278: dataIn1 = 32'd518
; 
32'd21279: dataIn1 = 32'd520
; 
32'd21280: dataIn1 = 32'd523
; 
32'd21281: dataIn1 = 32'd538
; 
32'd21282: dataIn1 = 32'd543
; 
32'd21283: dataIn1 = 32'd564
; 
32'd21284: dataIn1 = 32'd609
; 
32'd21285: dataIn1 = 32'd619
; 
32'd21286: dataIn1 = 32'd647
; 
32'd21287: dataIn1 = 32'd657
; 
32'd21288: dataIn1 = 32'd679
; 
32'd21289: dataIn1 = 32'd687
; 
32'd21290: dataIn1 = 32'd696
; 
32'd21291: dataIn1 = 32'd699
; 
32'd21292: dataIn1 = 32'd700
; 
32'd21293: dataIn1 = 32'd703
; 
32'd21294: dataIn1 = 32'd727
; 
32'd21295: dataIn1 = 32'd737
; 
32'd21296: dataIn1 = 32'd741
; 
32'd21297: dataIn1 = 32'd782
; 
32'd21298: dataIn1 = 32'd375
; 
32'd21299: dataIn1 = 32'd387
; 
32'd21300: dataIn1 = 32'd403
; 
32'd21301: dataIn1 = 32'd407
; 
32'd21302: dataIn1 = 32'd418
; 
32'd21303: dataIn1 = 32'd431
; 
32'd21304: dataIn1 = 32'd460
; 
32'd21305: dataIn1 = 32'd474
; 
32'd21306: dataIn1 = 32'd479
; 
32'd21307: dataIn1 = 32'd511
; 
32'd21308: dataIn1 = 32'd531
; 
32'd21309: dataIn1 = 32'd545
; 
32'd21310: dataIn1 = 32'd548
; 
32'd21311: dataIn1 = 32'd549
; 
32'd21312: dataIn1 = 32'd577
; 
32'd21313: dataIn1 = 32'd580
; 
32'd21314: dataIn1 = 32'd596
; 
32'd21315: dataIn1 = 32'd656
; 
32'd21316: dataIn1 = 32'd668
; 
32'd21317: dataIn1 = 32'd669
; 
32'd21318: dataIn1 = 32'd672
; 
32'd21319: dataIn1 = 32'd721
; 
32'd21320: dataIn1 = 32'd742
; 
32'd21321: dataIn1 = 32'd764
; 
32'd21322: dataIn1 = 32'd776
; 
32'd21323: dataIn1 = 32'd792
; 
32'd21324: dataIn1 = 32'd366
; 
32'd21325: dataIn1 = 32'd378
; 
32'd21326: dataIn1 = 32'd384
; 
32'd21327: dataIn1 = 32'd387
; 
32'd21328: dataIn1 = 32'd434
; 
32'd21329: dataIn1 = 32'd441
; 
32'd21330: dataIn1 = 32'd443
; 
32'd21331: dataIn1 = 32'd446
; 
32'd21332: dataIn1 = 32'd452
; 
32'd21333: dataIn1 = 32'd456
; 
32'd21334: dataIn1 = 32'd464
; 
32'd21335: dataIn1 = 32'd465
; 
32'd21336: dataIn1 = 32'd471
; 
32'd21337: dataIn1 = 32'd489
; 
32'd21338: dataIn1 = 32'd503
; 
32'd21339: dataIn1 = 32'd525
; 
32'd21340: dataIn1 = 32'd530
; 
32'd21341: dataIn1 = 32'd536
; 
32'd21342: dataIn1 = 32'd589
; 
32'd21343: dataIn1 = 32'd645
; 
32'd21344: dataIn1 = 32'd648
; 
32'd21345: dataIn1 = 32'd666
; 
32'd21346: dataIn1 = 32'd678
; 
32'd21347: dataIn1 = 32'd698
; 
32'd21348: dataIn1 = 32'd705
; 
32'd21349: dataIn1 = 32'd708
; 
32'd21350: dataIn1 = 32'd426
; 
32'd21351: dataIn1 = 32'd436
; 
32'd21352: dataIn1 = 32'd437
; 
32'd21353: dataIn1 = 32'd450
; 
32'd21354: dataIn1 = 32'd476
; 
32'd21355: dataIn1 = 32'd489
; 
32'd21356: dataIn1 = 32'd497
; 
32'd21357: dataIn1 = 32'd499
; 
32'd21358: dataIn1 = 32'd503
; 
32'd21359: dataIn1 = 32'd512
; 
32'd21360: dataIn1 = 32'd521
; 
32'd21361: dataIn1 = 32'd527
; 
32'd21362: dataIn1 = 32'd546
; 
32'd21363: dataIn1 = 32'd556
; 
32'd21364: dataIn1 = 32'd567
; 
32'd21365: dataIn1 = 32'd580
; 
32'd21366: dataIn1 = 32'd594
; 
32'd21367: dataIn1 = 32'd608
; 
32'd21368: dataIn1 = 32'd642
; 
32'd21369: dataIn1 = 32'd654
; 
32'd21370: dataIn1 = 32'd658
; 
32'd21371: dataIn1 = 32'd661
; 
32'd21372: dataIn1 = 32'd680
; 
32'd21373: dataIn1 = 32'd700
; 
32'd21374: dataIn1 = 32'd711
; 
32'd21375: dataIn1 = 32'd716
; 
32'd21376: dataIn1 = 32'd733
; 
32'd21377: dataIn1 = 32'd777
; 
32'd21378: dataIn1 = 32'd396
; 
32'd21379: dataIn1 = 32'd410
; 
32'd21380: dataIn1 = 32'd411
; 
32'd21381: dataIn1 = 32'd422
; 
32'd21382: dataIn1 = 32'd439
; 
32'd21383: dataIn1 = 32'd452
; 
32'd21384: dataIn1 = 32'd453
; 
32'd21385: dataIn1 = 32'd486
; 
32'd21386: dataIn1 = 32'd490
; 
32'd21387: dataIn1 = 32'd499
; 
32'd21388: dataIn1 = 32'd533
; 
32'd21389: dataIn1 = 32'd546
; 
32'd21390: dataIn1 = 32'd553
; 
32'd21391: dataIn1 = 32'd565
; 
32'd21392: dataIn1 = 32'd584
; 
32'd21393: dataIn1 = 32'd591
; 
32'd21394: dataIn1 = 32'd617
; 
32'd21395: dataIn1 = 32'd619
; 
32'd21396: dataIn1 = 32'd633
; 
32'd21397: dataIn1 = 32'd638
; 
32'd21398: dataIn1 = 32'd671
; 
32'd21399: dataIn1 = 32'd688
; 
32'd21400: dataIn1 = 32'd689
; 
32'd21401: dataIn1 = 32'd691
; 
32'd21402: dataIn1 = 32'd713
; 
32'd21403: dataIn1 = 32'd715
; 
32'd21404: dataIn1 = 32'd718
; 
32'd21405: dataIn1 = 32'd734
; 
32'd21406: dataIn1 = 32'd764
; 
32'd21407: dataIn1 = 32'd411
; 
32'd21408: dataIn1 = 32'd432
; 
32'd21409: dataIn1 = 32'd446
; 
32'd21410: dataIn1 = 32'd464
; 
32'd21411: dataIn1 = 32'd524
; 
32'd21412: dataIn1 = 32'd531
; 
32'd21413: dataIn1 = 32'd596
; 
32'd21414: dataIn1 = 32'd615
; 
32'd21415: dataIn1 = 32'd620
; 
32'd21416: dataIn1 = 32'd644
; 
32'd21417: dataIn1 = 32'd652
; 
32'd21418: dataIn1 = 32'd674
; 
32'd21419: dataIn1 = 32'd685
; 
32'd21420: dataIn1 = 32'd687
; 
32'd21421: dataIn1 = 32'd711
; 
32'd21422: dataIn1 = 32'd794
; 
32'd21423: dataIn1 = 32'd796
; 
32'd21424: dataIn1 = 32'd366
; 
32'd21425: dataIn1 = 32'd396
; 
32'd21426: dataIn1 = 32'd437
; 
32'd21427: dataIn1 = 32'd456
; 
32'd21428: dataIn1 = 32'd520
; 
32'd21429: dataIn1 = 32'd548
; 
32'd21430: dataIn1 = 32'd556
; 
32'd21431: dataIn1 = 32'd569
; 
32'd21432: dataIn1 = 32'd590
; 
32'd21433: dataIn1 = 32'd592
; 
32'd21434: dataIn1 = 32'd655
; 
32'd21435: dataIn1 = 32'd657
; 
32'd21436: dataIn1 = 32'd662
; 
32'd21437: dataIn1 = 32'd680
; 
32'd21438: dataIn1 = 32'd684
; 
32'd21439: dataIn1 = 32'd695
; 
32'd21440: dataIn1 = 32'd719
; 
32'd21441: dataIn1 = 32'd724
; 
32'd21442: dataIn1 = 32'd730
; 
32'd21443: dataIn1 = 32'd732
; 
32'd21444: dataIn1 = 32'd743
; 
32'd21445: dataIn1 = 32'd792
; 
32'd21446: dataIn1 = 32'd383
; 
32'd21447: dataIn1 = 32'd389
; 
32'd21448: dataIn1 = 32'd394
; 
32'd21449: dataIn1 = 32'd396
; 
32'd21450: dataIn1 = 32'd403
; 
32'd21451: dataIn1 = 32'd435
; 
32'd21452: dataIn1 = 32'd468
; 
32'd21453: dataIn1 = 32'd529
; 
32'd21454: dataIn1 = 32'd534
; 
32'd21455: dataIn1 = 32'd577
; 
32'd21456: dataIn1 = 32'd599
; 
32'd21457: dataIn1 = 32'd610
; 
32'd21458: dataIn1 = 32'd623
; 
32'd21459: dataIn1 = 32'd626
; 
32'd21460: dataIn1 = 32'd648
; 
32'd21461: dataIn1 = 32'd689
; 
32'd21462: dataIn1 = 32'd696
; 
32'd21463: dataIn1 = 32'd712
; 
32'd21464: dataIn1 = 32'd724
; 
32'd21465: dataIn1 = 32'd759
; 
32'd21466: dataIn1 = 32'd776
; 
32'd21467: dataIn1 = 32'd372
; 
32'd21468: dataIn1 = 32'd379
; 
32'd21469: dataIn1 = 32'd390
; 
32'd21470: dataIn1 = 32'd398
; 
32'd21471: dataIn1 = 32'd399
; 
32'd21472: dataIn1 = 32'd404
; 
32'd21473: dataIn1 = 32'd412
; 
32'd21474: dataIn1 = 32'd430
; 
32'd21475: dataIn1 = 32'd452
; 
32'd21476: dataIn1 = 32'd463
; 
32'd21477: dataIn1 = 32'd473
; 
32'd21478: dataIn1 = 32'd475
; 
32'd21479: dataIn1 = 32'd485
; 
32'd21480: dataIn1 = 32'd502
; 
32'd21481: dataIn1 = 32'd503
; 
32'd21482: dataIn1 = 32'd507
; 
32'd21483: dataIn1 = 32'd508
; 
32'd21484: dataIn1 = 32'd510
; 
32'd21485: dataIn1 = 32'd520
; 
32'd21486: dataIn1 = 32'd521
; 
32'd21487: dataIn1 = 32'd525
; 
32'd21488: dataIn1 = 32'd547
; 
32'd21489: dataIn1 = 32'd657
; 
32'd21490: dataIn1 = 32'd690
; 
32'd21491: dataIn1 = 32'd718
; 
32'd21492: dataIn1 = 32'd720
; 
32'd21493: dataIn1 = 32'd730
; 
32'd21494: dataIn1 = 32'd731
; 
32'd21495: dataIn1 = 32'd742
; 
32'd21496: dataIn1 = 32'd750
; 
32'd21497: dataIn1 = 32'd753
; 
32'd21498: dataIn1 = 32'd791
; 
32'd21499: dataIn1 = 32'd793
; 
32'd21500: dataIn1 = 32'd382
; 
32'd21501: dataIn1 = 32'd388
; 
32'd21502: dataIn1 = 32'd389
; 
32'd21503: dataIn1 = 32'd402
; 
32'd21504: dataIn1 = 32'd409
; 
32'd21505: dataIn1 = 32'd438
; 
32'd21506: dataIn1 = 32'd469
; 
32'd21507: dataIn1 = 32'd475
; 
32'd21508: dataIn1 = 32'd478
; 
32'd21509: dataIn1 = 32'd511
; 
32'd21510: dataIn1 = 32'd553
; 
32'd21511: dataIn1 = 32'd620
; 
32'd21512: dataIn1 = 32'd623
; 
32'd21513: dataIn1 = 32'd655
; 
32'd21514: dataIn1 = 32'd661
; 
32'd21515: dataIn1 = 32'd666
; 
32'd21516: dataIn1 = 32'd677
; 
32'd21517: dataIn1 = 32'd694
; 
32'd21518: dataIn1 = 32'd702
; 
32'd21519: dataIn1 = 32'd703
; 
32'd21520: dataIn1 = 32'd723
; 
32'd21521: dataIn1 = 32'd757
; 
32'd21522: dataIn1 = 32'd764
; 
32'd21523: dataIn1 = 32'd787
; 
32'd21524: dataIn1 = 32'd791
; 
32'd21525: dataIn1 = 32'd418
; 
32'd21526: dataIn1 = 32'd419
; 
32'd21527: dataIn1 = 32'd423
; 
32'd21528: dataIn1 = 32'd433
; 
32'd21529: dataIn1 = 32'd506
; 
32'd21530: dataIn1 = 32'd512
; 
32'd21531: dataIn1 = 32'd528
; 
32'd21532: dataIn1 = 32'd541
; 
32'd21533: dataIn1 = 32'd544
; 
32'd21534: dataIn1 = 32'd551
; 
32'd21535: dataIn1 = 32'd578
; 
32'd21536: dataIn1 = 32'd634
; 
32'd21537: dataIn1 = 32'd652
; 
32'd21538: dataIn1 = 32'd653
; 
32'd21539: dataIn1 = 32'd655
; 
32'd21540: dataIn1 = 32'd694
; 
32'd21541: dataIn1 = 32'd718
; 
32'd21542: dataIn1 = 32'd767
; 
32'd21543: dataIn1 = 32'd775
; 
32'd21544: dataIn1 = 32'd380
; 
32'd21545: dataIn1 = 32'd382
; 
32'd21546: dataIn1 = 32'd385
; 
32'd21547: dataIn1 = 32'd389
; 
32'd21548: dataIn1 = 32'd397
; 
32'd21549: dataIn1 = 32'd401
; 
32'd21550: dataIn1 = 32'd414
; 
32'd21551: dataIn1 = 32'd439
; 
32'd21552: dataIn1 = 32'd456
; 
32'd21553: dataIn1 = 32'd506
; 
32'd21554: dataIn1 = 32'd508
; 
32'd21555: dataIn1 = 32'd511
; 
32'd21556: dataIn1 = 32'd531
; 
32'd21557: dataIn1 = 32'd560
; 
32'd21558: dataIn1 = 32'd582
; 
32'd21559: dataIn1 = 32'd583
; 
32'd21560: dataIn1 = 32'd594
; 
32'd21561: dataIn1 = 32'd610
; 
32'd21562: dataIn1 = 32'd627
; 
32'd21563: dataIn1 = 32'd631
; 
32'd21564: dataIn1 = 32'd647
; 
32'd21565: dataIn1 = 32'd648
; 
32'd21566: dataIn1 = 32'd718
; 
32'd21567: dataIn1 = 32'd738
; 
32'd21568: dataIn1 = 32'd749
; 
32'd21569: dataIn1 = 32'd762
; 
32'd21570: dataIn1 = 32'd769
; 
32'd21571: dataIn1 = 32'd372
; 
32'd21572: dataIn1 = 32'd410
; 
32'd21573: dataIn1 = 32'd420
; 
32'd21574: dataIn1 = 32'd423
; 
32'd21575: dataIn1 = 32'd518
; 
32'd21576: dataIn1 = 32'd520
; 
32'd21577: dataIn1 = 32'd531
; 
32'd21578: dataIn1 = 32'd578
; 
32'd21579: dataIn1 = 32'd636
; 
32'd21580: dataIn1 = 32'd650
; 
32'd21581: dataIn1 = 32'd663
; 
32'd21582: dataIn1 = 32'd679
; 
32'd21583: dataIn1 = 32'd682
; 
32'd21584: dataIn1 = 32'd705
; 
32'd21585: dataIn1 = 32'd734
; 
32'd21586: dataIn1 = 32'd758
; 
32'd21587: dataIn1 = 32'd787
; 
32'd21588: dataIn1 = 32'd791
; 
32'd21589: dataIn1 = 32'd373
; 
32'd21590: dataIn1 = 32'd391
; 
32'd21591: dataIn1 = 32'd401
; 
32'd21592: dataIn1 = 32'd425
; 
32'd21593: dataIn1 = 32'd426
; 
32'd21594: dataIn1 = 32'd429
; 
32'd21595: dataIn1 = 32'd448
; 
32'd21596: dataIn1 = 32'd450
; 
32'd21597: dataIn1 = 32'd462
; 
32'd21598: dataIn1 = 32'd467
; 
32'd21599: dataIn1 = 32'd498
; 
32'd21600: dataIn1 = 32'd499
; 
32'd21601: dataIn1 = 32'd509
; 
32'd21602: dataIn1 = 32'd550
; 
32'd21603: dataIn1 = 32'd567
; 
32'd21604: dataIn1 = 32'd606
; 
32'd21605: dataIn1 = 32'd607
; 
32'd21606: dataIn1 = 32'd609
; 
32'd21607: dataIn1 = 32'd614
; 
32'd21608: dataIn1 = 32'd624
; 
32'd21609: dataIn1 = 32'd627
; 
32'd21610: dataIn1 = 32'd655
; 
32'd21611: dataIn1 = 32'd716
; 
32'd21612: dataIn1 = 32'd741
; 
32'd21613: dataIn1 = 32'd761
; 
32'd21614: dataIn1 = 32'd375
; 
32'd21615: dataIn1 = 32'd391
; 
32'd21616: dataIn1 = 32'd396
; 
32'd21617: dataIn1 = 32'd405
; 
32'd21618: dataIn1 = 32'd447
; 
32'd21619: dataIn1 = 32'd456
; 
32'd21620: dataIn1 = 32'd459
; 
32'd21621: dataIn1 = 32'd489
; 
32'd21622: dataIn1 = 32'd504
; 
32'd21623: dataIn1 = 32'd528
; 
32'd21624: dataIn1 = 32'd540
; 
32'd21625: dataIn1 = 32'd571
; 
32'd21626: dataIn1 = 32'd578
; 
32'd21627: dataIn1 = 32'd588
; 
32'd21628: dataIn1 = 32'd600
; 
32'd21629: dataIn1 = 32'd630
; 
32'd21630: dataIn1 = 32'd633
; 
32'd21631: dataIn1 = 32'd634
; 
32'd21632: dataIn1 = 32'd674
; 
32'd21633: dataIn1 = 32'd683
; 
32'd21634: dataIn1 = 32'd685
; 
32'd21635: dataIn1 = 32'd706
; 
32'd21636: dataIn1 = 32'd733
; 
32'd21637: dataIn1 = 32'd734
; 
32'd21638: dataIn1 = 32'd750
; 
32'd21639: dataIn1 = 32'd757
; 
32'd21640: dataIn1 = 32'd763
; 
32'd21641: dataIn1 = 32'd787
; 
32'd21642: dataIn1 = 32'd389
; 
32'd21643: dataIn1 = 32'd422
; 
32'd21644: dataIn1 = 32'd432
; 
32'd21645: dataIn1 = 32'd437
; 
32'd21646: dataIn1 = 32'd444
; 
32'd21647: dataIn1 = 32'd445
; 
32'd21648: dataIn1 = 32'd507
; 
32'd21649: dataIn1 = 32'd526
; 
32'd21650: dataIn1 = 32'd532
; 
32'd21651: dataIn1 = 32'd544
; 
32'd21652: dataIn1 = 32'd590
; 
32'd21653: dataIn1 = 32'd629
; 
32'd21654: dataIn1 = 32'd635
; 
32'd21655: dataIn1 = 32'd644
; 
32'd21656: dataIn1 = 32'd653
; 
32'd21657: dataIn1 = 32'd655
; 
32'd21658: dataIn1 = 32'd682
; 
32'd21659: dataIn1 = 32'd690
; 
32'd21660: dataIn1 = 32'd710
; 
32'd21661: dataIn1 = 32'd716
; 
32'd21662: dataIn1 = 32'd736
; 
32'd21663: dataIn1 = 32'd748
; 
32'd21664: dataIn1 = 32'd760
; 
32'd21665: dataIn1 = 32'd769
; 
32'd21666: dataIn1 = 32'd798
; 
32'd21667: dataIn1 = 32'd397
; 
32'd21668: dataIn1 = 32'd402
; 
32'd21669: dataIn1 = 32'd413
; 
32'd21670: dataIn1 = 32'd433
; 
32'd21671: dataIn1 = 32'd437
; 
32'd21672: dataIn1 = 32'd458
; 
32'd21673: dataIn1 = 32'd493
; 
32'd21674: dataIn1 = 32'd496
; 
32'd21675: dataIn1 = 32'd499
; 
32'd21676: dataIn1 = 32'd504
; 
32'd21677: dataIn1 = 32'd539
; 
32'd21678: dataIn1 = 32'd549
; 
32'd21679: dataIn1 = 32'd566
; 
32'd21680: dataIn1 = 32'd621
; 
32'd21681: dataIn1 = 32'd624
; 
32'd21682: dataIn1 = 32'd680
; 
32'd21683: dataIn1 = 32'd683
; 
32'd21684: dataIn1 = 32'd742
; 
32'd21685: dataIn1 = 32'd762
; 
32'd21686: dataIn1 = 32'd771
; 
32'd21687: dataIn1 = 32'd788
; 
32'd21688: dataIn1 = 32'd791
; 
32'd21689: dataIn1 = 32'd799
; 
32'd21690: dataIn1 = 32'd376
; 
32'd21691: dataIn1 = 32'd409
; 
32'd21692: dataIn1 = 32'd421
; 
32'd21693: dataIn1 = 32'd426
; 
32'd21694: dataIn1 = 32'd432
; 
32'd21695: dataIn1 = 32'd465
; 
32'd21696: dataIn1 = 32'd478
; 
32'd21697: dataIn1 = 32'd483
; 
32'd21698: dataIn1 = 32'd490
; 
32'd21699: dataIn1 = 32'd494
; 
32'd21700: dataIn1 = 32'd496
; 
32'd21701: dataIn1 = 32'd501
; 
32'd21702: dataIn1 = 32'd512
; 
32'd21703: dataIn1 = 32'd521
; 
32'd21704: dataIn1 = 32'd536
; 
32'd21705: dataIn1 = 32'd542
; 
32'd21706: dataIn1 = 32'd562
; 
32'd21707: dataIn1 = 32'd583
; 
32'd21708: dataIn1 = 32'd607
; 
32'd21709: dataIn1 = 32'd624
; 
32'd21710: dataIn1 = 32'd635
; 
32'd21711: dataIn1 = 32'd640
; 
32'd21712: dataIn1 = 32'd652
; 
32'd21713: dataIn1 = 32'd667
; 
32'd21714: dataIn1 = 32'd678
; 
32'd21715: dataIn1 = 32'd684
; 
32'd21716: dataIn1 = 32'd746
; 
32'd21717: dataIn1 = 32'd749
; 
32'd21718: dataIn1 = 32'd771
; 
32'd21719: dataIn1 = 32'd792
; 
32'd21720: dataIn1 = 32'd377
; 
32'd21721: dataIn1 = 32'd399
; 
32'd21722: dataIn1 = 32'd401
; 
32'd21723: dataIn1 = 32'd405
; 
32'd21724: dataIn1 = 32'd443
; 
32'd21725: dataIn1 = 32'd478
; 
32'd21726: dataIn1 = 32'd483
; 
32'd21727: dataIn1 = 32'd497
; 
32'd21728: dataIn1 = 32'd522
; 
32'd21729: dataIn1 = 32'd537
; 
32'd21730: dataIn1 = 32'd562
; 
32'd21731: dataIn1 = 32'd567
; 
32'd21732: dataIn1 = 32'd583
; 
32'd21733: dataIn1 = 32'd626
; 
32'd21734: dataIn1 = 32'd644
; 
32'd21735: dataIn1 = 32'd677
; 
32'd21736: dataIn1 = 32'd686
; 
32'd21737: dataIn1 = 32'd687
; 
32'd21738: dataIn1 = 32'd689
; 
32'd21739: dataIn1 = 32'd708
; 
32'd21740: dataIn1 = 32'd717
; 
32'd21741: dataIn1 = 32'd736
; 
32'd21742: dataIn1 = 32'd743
; 
32'd21743: dataIn1 = 32'd768
; 
32'd21744: dataIn1 = 32'd782
; 
32'd21745: dataIn1 = 32'd379
; 
32'd21746: dataIn1 = 32'd384
; 
32'd21747: dataIn1 = 32'd424
; 
32'd21748: dataIn1 = 32'd436
; 
32'd21749: dataIn1 = 32'd446
; 
32'd21750: dataIn1 = 32'd453
; 
32'd21751: dataIn1 = 32'd459
; 
32'd21752: dataIn1 = 32'd503
; 
32'd21753: dataIn1 = 32'd507
; 
32'd21754: dataIn1 = 32'd512
; 
32'd21755: dataIn1 = 32'd523
; 
32'd21756: dataIn1 = 32'd538
; 
32'd21757: dataIn1 = 32'd539
; 
32'd21758: dataIn1 = 32'd541
; 
32'd21759: dataIn1 = 32'd562
; 
32'd21760: dataIn1 = 32'd580
; 
32'd21761: dataIn1 = 32'd602
; 
32'd21762: dataIn1 = 32'd614
; 
32'd21763: dataIn1 = 32'd620
; 
32'd21764: dataIn1 = 32'd639
; 
32'd21765: dataIn1 = 32'd643
; 
32'd21766: dataIn1 = 32'd653
; 
32'd21767: dataIn1 = 32'd674
; 
32'd21768: dataIn1 = 32'd698
; 
32'd21769: dataIn1 = 32'd701
; 
32'd21770: dataIn1 = 32'd706
; 
32'd21771: dataIn1 = 32'd735
; 
32'd21772: dataIn1 = 32'd764
; 
32'd21773: dataIn1 = 32'd797
; 
32'd21774: dataIn1 = 32'd377
; 
32'd21775: dataIn1 = 32'd383
; 
32'd21776: dataIn1 = 32'd413
; 
32'd21777: dataIn1 = 32'd428
; 
32'd21778: dataIn1 = 32'd442
; 
32'd21779: dataIn1 = 32'd450
; 
32'd21780: dataIn1 = 32'd464
; 
32'd21781: dataIn1 = 32'd489
; 
32'd21782: dataIn1 = 32'd508
; 
32'd21783: dataIn1 = 32'd510
; 
32'd21784: dataIn1 = 32'd520
; 
32'd21785: dataIn1 = 32'd527
; 
32'd21786: dataIn1 = 32'd538
; 
32'd21787: dataIn1 = 32'd550
; 
32'd21788: dataIn1 = 32'd556
; 
32'd21789: dataIn1 = 32'd570
; 
32'd21790: dataIn1 = 32'd580
; 
32'd21791: dataIn1 = 32'd603
; 
32'd21792: dataIn1 = 32'd614
; 
32'd21793: dataIn1 = 32'd623
; 
32'd21794: dataIn1 = 32'd651
; 
32'd21795: dataIn1 = 32'd674
; 
32'd21796: dataIn1 = 32'd708
; 
32'd21797: dataIn1 = 32'd720
; 
32'd21798: dataIn1 = 32'd740
; 
32'd21799: dataIn1 = 32'd751
; 
32'd21800: dataIn1 = 32'd755
; 
32'd21801: dataIn1 = 32'd757
; 
32'd21802: dataIn1 = 32'd758
; 
32'd21803: dataIn1 = 32'd766
; 
32'd21804: dataIn1 = 32'd790
; 
32'd21805: dataIn1 = 32'd797
; 
32'd21806: dataIn1 = 32'd387
; 
32'd21807: dataIn1 = 32'd388
; 
32'd21808: dataIn1 = 32'd393
; 
32'd21809: dataIn1 = 32'd398
; 
32'd21810: dataIn1 = 32'd440
; 
32'd21811: dataIn1 = 32'd441
; 
32'd21812: dataIn1 = 32'd443
; 
32'd21813: dataIn1 = 32'd458
; 
32'd21814: dataIn1 = 32'd459
; 
32'd21815: dataIn1 = 32'd488
; 
32'd21816: dataIn1 = 32'd525
; 
32'd21817: dataIn1 = 32'd547
; 
32'd21818: dataIn1 = 32'd553
; 
32'd21819: dataIn1 = 32'd558
; 
32'd21820: dataIn1 = 32'd583
; 
32'd21821: dataIn1 = 32'd591
; 
32'd21822: dataIn1 = 32'd593
; 
32'd21823: dataIn1 = 32'd600
; 
32'd21824: dataIn1 = 32'd630
; 
32'd21825: dataIn1 = 32'd681
; 
32'd21826: dataIn1 = 32'd696
; 
32'd21827: dataIn1 = 32'd705
; 
32'd21828: dataIn1 = 32'd740
; 
32'd21829: dataIn1 = 32'd742
; 
32'd21830: dataIn1 = 32'd749
; 
32'd21831: dataIn1 = 32'd756
; 
32'd21832: dataIn1 = 32'd764
; 
32'd21833: dataIn1 = 32'd783
; 
32'd21834: dataIn1 = 32'd798
; 
32'd21835: dataIn1 = 32'd385
; 
32'd21836: dataIn1 = 32'd392
; 
32'd21837: dataIn1 = 32'd419
; 
32'd21838: dataIn1 = 32'd445
; 
32'd21839: dataIn1 = 32'd451
; 
32'd21840: dataIn1 = 32'd485
; 
32'd21841: dataIn1 = 32'd517
; 
32'd21842: dataIn1 = 32'd519
; 
32'd21843: dataIn1 = 32'd563
; 
32'd21844: dataIn1 = 32'd573
; 
32'd21845: dataIn1 = 32'd593
; 
32'd21846: dataIn1 = 32'd601
; 
32'd21847: dataIn1 = 32'd632
; 
32'd21848: dataIn1 = 32'd678
; 
32'd21849: dataIn1 = 32'd688
; 
32'd21850: dataIn1 = 32'd696
; 
32'd21851: dataIn1 = 32'd710
; 
32'd21852: dataIn1 = 32'd714
; 
32'd21853: dataIn1 = 32'd733
; 
32'd21854: dataIn1 = 32'd741
; 
32'd21855: dataIn1 = 32'd743
; 
32'd21856: dataIn1 = 32'd758
; 
32'd21857: dataIn1 = 32'd788
; 
32'd21858: dataIn1 = 32'd385
; 
32'd21859: dataIn1 = 32'd414
; 
32'd21860: dataIn1 = 32'd430
; 
32'd21861: dataIn1 = 32'd466
; 
32'd21862: dataIn1 = 32'd469
; 
32'd21863: dataIn1 = 32'd494
; 
32'd21864: dataIn1 = 32'd506
; 
32'd21865: dataIn1 = 32'd556
; 
32'd21866: dataIn1 = 32'd562
; 
32'd21867: dataIn1 = 32'd566
; 
32'd21868: dataIn1 = 32'd625
; 
32'd21869: dataIn1 = 32'd670
; 
32'd21870: dataIn1 = 32'd681
; 
32'd21871: dataIn1 = 32'd685
; 
32'd21872: dataIn1 = 32'd731
; 
32'd21873: dataIn1 = 32'd740
; 
32'd21874: dataIn1 = 32'd763
; 
32'd21875: dataIn1 = 32'd779
; 
32'd21876: dataIn1 = 32'd382
; 
32'd21877: dataIn1 = 32'd417
; 
32'd21878: dataIn1 = 32'd426
; 
32'd21879: dataIn1 = 32'd444
; 
32'd21880: dataIn1 = 32'd461
; 
32'd21881: dataIn1 = 32'd466
; 
32'd21882: dataIn1 = 32'd473
; 
32'd21883: dataIn1 = 32'd485
; 
32'd21884: dataIn1 = 32'd490
; 
32'd21885: dataIn1 = 32'd500
; 
32'd21886: dataIn1 = 32'd503
; 
32'd21887: dataIn1 = 32'd525
; 
32'd21888: dataIn1 = 32'd548
; 
32'd21889: dataIn1 = 32'd584
; 
32'd21890: dataIn1 = 32'd591
; 
32'd21891: dataIn1 = 32'd601
; 
32'd21892: dataIn1 = 32'd623
; 
32'd21893: dataIn1 = 32'd661
; 
32'd21894: dataIn1 = 32'd699
; 
32'd21895: dataIn1 = 32'd708
; 
32'd21896: dataIn1 = 32'd726
; 
32'd21897: dataIn1 = 32'd739
; 
32'd21898: dataIn1 = 32'd785
; 
32'd21899: dataIn1 = 32'd383
; 
32'd21900: dataIn1 = 32'd408
; 
32'd21901: dataIn1 = 32'd410
; 
32'd21902: dataIn1 = 32'd424
; 
32'd21903: dataIn1 = 32'd433
; 
32'd21904: dataIn1 = 32'd434
; 
32'd21905: dataIn1 = 32'd435
; 
32'd21906: dataIn1 = 32'd441
; 
32'd21907: dataIn1 = 32'd443
; 
32'd21908: dataIn1 = 32'd446
; 
32'd21909: dataIn1 = 32'd486
; 
32'd21910: dataIn1 = 32'd487
; 
32'd21911: dataIn1 = 32'd526
; 
32'd21912: dataIn1 = 32'd550
; 
32'd21913: dataIn1 = 32'd551
; 
32'd21914: dataIn1 = 32'd578
; 
32'd21915: dataIn1 = 32'd604
; 
32'd21916: dataIn1 = 32'd621
; 
32'd21917: dataIn1 = 32'd658
; 
32'd21918: dataIn1 = 32'd720
; 
32'd21919: dataIn1 = 32'd726
; 
32'd21920: dataIn1 = 32'd743
; 
32'd21921: dataIn1 = 32'd748
; 
32'd21922: dataIn1 = 32'd753
; 
32'd21923: dataIn1 = 32'd782
; 
32'd21924: dataIn1 = 32'd783
; 
32'd21925: dataIn1 = 32'd789
; 
32'd21926: dataIn1 = 32'd390
; 
32'd21927: dataIn1 = 32'd402
; 
32'd21928: dataIn1 = 32'd418
; 
32'd21929: dataIn1 = 32'd436
; 
32'd21930: dataIn1 = 32'd441
; 
32'd21931: dataIn1 = 32'd453
; 
32'd21932: dataIn1 = 32'd465
; 
32'd21933: dataIn1 = 32'd472
; 
32'd21934: dataIn1 = 32'd479
; 
32'd21935: dataIn1 = 32'd502
; 
32'd21936: dataIn1 = 32'd523
; 
32'd21937: dataIn1 = 32'd546
; 
32'd21938: dataIn1 = 32'd564
; 
32'd21939: dataIn1 = 32'd565
; 
32'd21940: dataIn1 = 32'd576
; 
32'd21941: dataIn1 = 32'd604
; 
32'd21942: dataIn1 = 32'd606
; 
32'd21943: dataIn1 = 32'd643
; 
32'd21944: dataIn1 = 32'd644
; 
32'd21945: dataIn1 = 32'd649
; 
32'd21946: dataIn1 = 32'd674
; 
32'd21947: dataIn1 = 32'd678
; 
32'd21948: dataIn1 = 32'd730
; 
32'd21949: dataIn1 = 32'd745
; 
32'd21950: dataIn1 = 32'd765
; 
32'd21951: dataIn1 = 32'd782
; 
32'd21952: dataIn1 = 32'd785
; 
32'd21953: dataIn1 = 32'd384
; 
32'd21954: dataIn1 = 32'd388
; 
32'd21955: dataIn1 = 32'd391
; 
32'd21956: dataIn1 = 32'd412
; 
32'd21957: dataIn1 = 32'd418
; 
32'd21958: dataIn1 = 32'd429
; 
32'd21959: dataIn1 = 32'd459
; 
32'd21960: dataIn1 = 32'd467
; 
32'd21961: dataIn1 = 32'd469
; 
32'd21962: dataIn1 = 32'd476
; 
32'd21963: dataIn1 = 32'd479
; 
32'd21964: dataIn1 = 32'd543
; 
32'd21965: dataIn1 = 32'd565
; 
32'd21966: dataIn1 = 32'd585
; 
32'd21967: dataIn1 = 32'd598
; 
32'd21968: dataIn1 = 32'd602
; 
32'd21969: dataIn1 = 32'd620
; 
32'd21970: dataIn1 = 32'd622
; 
32'd21971: dataIn1 = 32'd626
; 
32'd21972: dataIn1 = 32'd650
; 
32'd21973: dataIn1 = 32'd668
; 
32'd21974: dataIn1 = 32'd673
; 
32'd21975: dataIn1 = 32'd677
; 
32'd21976: dataIn1 = 32'd683
; 
32'd21977: dataIn1 = 32'd684
; 
32'd21978: dataIn1 = 32'd687
; 
32'd21979: dataIn1 = 32'd700
; 
32'd21980: dataIn1 = 32'd723
; 
32'd21981: dataIn1 = 32'd725
; 
32'd21982: dataIn1 = 32'd748
; 
32'd21983: dataIn1 = 32'd752
; 
32'd21984: dataIn1 = 32'd754
; 
32'd21985: dataIn1 = 32'd755
; 
32'd21986: dataIn1 = 32'd759
; 
32'd21987: dataIn1 = 32'd782
; 
32'd21988: dataIn1 = 32'd797
; 
32'd21989: dataIn1 = 32'd395
; 
32'd21990: dataIn1 = 32'd407
; 
32'd21991: dataIn1 = 32'd419
; 
32'd21992: dataIn1 = 32'd427
; 
32'd21993: dataIn1 = 32'd443
; 
32'd21994: dataIn1 = 32'd449
; 
32'd21995: dataIn1 = 32'd450
; 
32'd21996: dataIn1 = 32'd459
; 
32'd21997: dataIn1 = 32'd481
; 
32'd21998: dataIn1 = 32'd488
; 
32'd21999: dataIn1 = 32'd503
; 
32'd22000: dataIn1 = 32'd515
; 
32'd22001: dataIn1 = 32'd535
; 
32'd22002: dataIn1 = 32'd538
; 
32'd22003: dataIn1 = 32'd553
; 
32'd22004: dataIn1 = 32'd590
; 
32'd22005: dataIn1 = 32'd652
; 
32'd22006: dataIn1 = 32'd654
; 
32'd22007: dataIn1 = 32'd667
; 
32'd22008: dataIn1 = 32'd687
; 
32'd22009: dataIn1 = 32'd698
; 
32'd22010: dataIn1 = 32'd715
; 
32'd22011: dataIn1 = 32'd726
; 
32'd22012: dataIn1 = 32'd768
; 
32'd22013: dataIn1 = 32'd773
; 
32'd22014: dataIn1 = 32'd390
; 
32'd22015: dataIn1 = 32'd395
; 
32'd22016: dataIn1 = 32'd458
; 
32'd22017: dataIn1 = 32'd523
; 
32'd22018: dataIn1 = 32'd539
; 
32'd22019: dataIn1 = 32'd540
; 
32'd22020: dataIn1 = 32'd555
; 
32'd22021: dataIn1 = 32'd573
; 
32'd22022: dataIn1 = 32'd584
; 
32'd22023: dataIn1 = 32'd586
; 
32'd22024: dataIn1 = 32'd589
; 
32'd22025: dataIn1 = 32'd593
; 
32'd22026: dataIn1 = 32'd616
; 
32'd22027: dataIn1 = 32'd619
; 
32'd22028: dataIn1 = 32'd639
; 
32'd22029: dataIn1 = 32'd665
; 
32'd22030: dataIn1 = 32'd666
; 
32'd22031: dataIn1 = 32'd684
; 
32'd22032: dataIn1 = 32'd725
; 
32'd22033: dataIn1 = 32'd731
; 
32'd22034: dataIn1 = 32'd748
; 
32'd22035: dataIn1 = 32'd760
; 
32'd22036: dataIn1 = 32'd422
; 
32'd22037: dataIn1 = 32'd454
; 
32'd22038: dataIn1 = 32'd468
; 
32'd22039: dataIn1 = 32'd484
; 
32'd22040: dataIn1 = 32'd501
; 
32'd22041: dataIn1 = 32'd507
; 
32'd22042: dataIn1 = 32'd519
; 
32'd22043: dataIn1 = 32'd524
; 
32'd22044: dataIn1 = 32'd537
; 
32'd22045: dataIn1 = 32'd552
; 
32'd22046: dataIn1 = 32'd556
; 
32'd22047: dataIn1 = 32'd577
; 
32'd22048: dataIn1 = 32'd593
; 
32'd22049: dataIn1 = 32'd606
; 
32'd22050: dataIn1 = 32'd619
; 
32'd22051: dataIn1 = 32'd624
; 
32'd22052: dataIn1 = 32'd651
; 
32'd22053: dataIn1 = 32'd653
; 
32'd22054: dataIn1 = 32'd667
; 
32'd22055: dataIn1 = 32'd668
; 
32'd22056: dataIn1 = 32'd679
; 
32'd22057: dataIn1 = 32'd680
; 
32'd22058: dataIn1 = 32'd688
; 
32'd22059: dataIn1 = 32'd700
; 
32'd22060: dataIn1 = 32'd712
; 
32'd22061: dataIn1 = 32'd719
; 
32'd22062: dataIn1 = 32'd742
; 
32'd22063: dataIn1 = 32'd745
; 
32'd22064: dataIn1 = 32'd772
; 
32'd22065: dataIn1 = 32'd800
; 
32'd22066: dataIn1 = 32'd425
; 
32'd22067: dataIn1 = 32'd427
; 
32'd22068: dataIn1 = 32'd458
; 
32'd22069: dataIn1 = 32'd470
; 
32'd22070: dataIn1 = 32'd507
; 
32'd22071: dataIn1 = 32'd535
; 
32'd22072: dataIn1 = 32'd546
; 
32'd22073: dataIn1 = 32'd560
; 
32'd22074: dataIn1 = 32'd609
; 
32'd22075: dataIn1 = 32'd612
; 
32'd22076: dataIn1 = 32'd614
; 
32'd22077: dataIn1 = 32'd629
; 
32'd22078: dataIn1 = 32'd648
; 
32'd22079: dataIn1 = 32'd651
; 
32'd22080: dataIn1 = 32'd665
; 
32'd22081: dataIn1 = 32'd680
; 
32'd22082: dataIn1 = 32'd689
; 
32'd22083: dataIn1 = 32'd724
; 
32'd22084: dataIn1 = 32'd739
; 
32'd22085: dataIn1 = 32'd740
; 
32'd22086: dataIn1 = 32'd758
; 
32'd22087: dataIn1 = 32'd767
; 
32'd22088: dataIn1 = 32'd772
; 
32'd22089: dataIn1 = 32'd777
; 
32'd22090: dataIn1 = 32'd787
; 
32'd22091: dataIn1 = 32'd409
; 
32'd22092: dataIn1 = 32'd412
; 
32'd22093: dataIn1 = 32'd438
; 
32'd22094: dataIn1 = 32'd467
; 
32'd22095: dataIn1 = 32'd470
; 
32'd22096: dataIn1 = 32'd485
; 
32'd22097: dataIn1 = 32'd530
; 
32'd22098: dataIn1 = 32'd549
; 
32'd22099: dataIn1 = 32'd564
; 
32'd22100: dataIn1 = 32'd569
; 
32'd22101: dataIn1 = 32'd606
; 
32'd22102: dataIn1 = 32'd611
; 
32'd22103: dataIn1 = 32'd627
; 
32'd22104: dataIn1 = 32'd629
; 
32'd22105: dataIn1 = 32'd718
; 
32'd22106: dataIn1 = 32'd722
; 
32'd22107: dataIn1 = 32'd723
; 
32'd22108: dataIn1 = 32'd729
; 
32'd22109: dataIn1 = 32'd744
; 
32'd22110: dataIn1 = 32'd749
; 
32'd22111: dataIn1 = 32'd787
; 
32'd22112: dataIn1 = 32'd796
; 
32'd22113: dataIn1 = 32'd408
; 
32'd22114: dataIn1 = 32'd422
; 
32'd22115: dataIn1 = 32'd424
; 
32'd22116: dataIn1 = 32'd426
; 
32'd22117: dataIn1 = 32'd434
; 
32'd22118: dataIn1 = 32'd436
; 
32'd22119: dataIn1 = 32'd481
; 
32'd22120: dataIn1 = 32'd542
; 
32'd22121: dataIn1 = 32'd564
; 
32'd22122: dataIn1 = 32'd569
; 
32'd22123: dataIn1 = 32'd590
; 
32'd22124: dataIn1 = 32'd599
; 
32'd22125: dataIn1 = 32'd615
; 
32'd22126: dataIn1 = 32'd623
; 
32'd22127: dataIn1 = 32'd656
; 
32'd22128: dataIn1 = 32'd677
; 
32'd22129: dataIn1 = 32'd692
; 
32'd22130: dataIn1 = 32'd712
; 
32'd22131: dataIn1 = 32'd729
; 
32'd22132: dataIn1 = 32'd736
; 
32'd22133: dataIn1 = 32'd752
; 
32'd22134: dataIn1 = 32'd761
; 
32'd22135: dataIn1 = 32'd788
; 
32'd22136: dataIn1 = 32'd799
; 
32'd22137: dataIn1 = 32'd405
; 
32'd22138: dataIn1 = 32'd437
; 
32'd22139: dataIn1 = 32'd464
; 
32'd22140: dataIn1 = 32'd472
; 
32'd22141: dataIn1 = 32'd479
; 
32'd22142: dataIn1 = 32'd513
; 
32'd22143: dataIn1 = 32'd517
; 
32'd22144: dataIn1 = 32'd518
; 
32'd22145: dataIn1 = 32'd526
; 
32'd22146: dataIn1 = 32'd531
; 
32'd22147: dataIn1 = 32'd533
; 
32'd22148: dataIn1 = 32'd586
; 
32'd22149: dataIn1 = 32'd595
; 
32'd22150: dataIn1 = 32'd608
; 
32'd22151: dataIn1 = 32'd627
; 
32'd22152: dataIn1 = 32'd641
; 
32'd22153: dataIn1 = 32'd675
; 
32'd22154: dataIn1 = 32'd676
; 
32'd22155: dataIn1 = 32'd690
; 
32'd22156: dataIn1 = 32'd700
; 
32'd22157: dataIn1 = 32'd702
; 
32'd22158: dataIn1 = 32'd704
; 
32'd22159: dataIn1 = 32'd708
; 
32'd22160: dataIn1 = 32'd713
; 
32'd22161: dataIn1 = 32'd724
; 
32'd22162: dataIn1 = 32'd728
; 
32'd22163: dataIn1 = 32'd730
; 
32'd22164: dataIn1 = 32'd734
; 
32'd22165: dataIn1 = 32'd751
; 
32'd22166: dataIn1 = 32'd781
; 
32'd22167: dataIn1 = 32'd795
; 
32'd22168: dataIn1 = 32'd397
; 
32'd22169: dataIn1 = 32'd404
; 
32'd22170: dataIn1 = 32'd415
; 
32'd22171: dataIn1 = 32'd423
; 
32'd22172: dataIn1 = 32'd433
; 
32'd22173: dataIn1 = 32'd457
; 
32'd22174: dataIn1 = 32'd506
; 
32'd22175: dataIn1 = 32'd543
; 
32'd22176: dataIn1 = 32'd546
; 
32'd22177: dataIn1 = 32'd569
; 
32'd22178: dataIn1 = 32'd578
; 
32'd22179: dataIn1 = 32'd584
; 
32'd22180: dataIn1 = 32'd618
; 
32'd22181: dataIn1 = 32'd637
; 
32'd22182: dataIn1 = 32'd639
; 
32'd22183: dataIn1 = 32'd646
; 
32'd22184: dataIn1 = 32'd660
; 
32'd22185: dataIn1 = 32'd686
; 
32'd22186: dataIn1 = 32'd689
; 
32'd22187: dataIn1 = 32'd701
; 
32'd22188: dataIn1 = 32'd706
; 
32'd22189: dataIn1 = 32'd711
; 
32'd22190: dataIn1 = 32'd744
; 
32'd22191: dataIn1 = 32'd748
; 
32'd22192: dataIn1 = 32'd424
; 
32'd22193: dataIn1 = 32'd432
; 
32'd22194: dataIn1 = 32'd458
; 
32'd22195: dataIn1 = 32'd480
; 
32'd22196: dataIn1 = 32'd497
; 
32'd22197: dataIn1 = 32'd501
; 
32'd22198: dataIn1 = 32'd519
; 
32'd22199: dataIn1 = 32'd521
; 
32'd22200: dataIn1 = 32'd523
; 
32'd22201: dataIn1 = 32'd532
; 
32'd22202: dataIn1 = 32'd541
; 
32'd22203: dataIn1 = 32'd544
; 
32'd22204: dataIn1 = 32'd550
; 
32'd22205: dataIn1 = 32'd556
; 
32'd22206: dataIn1 = 32'd629
; 
32'd22207: dataIn1 = 32'd631
; 
32'd22208: dataIn1 = 32'd647
; 
32'd22209: dataIn1 = 32'd670
; 
32'd22210: dataIn1 = 32'd671
; 
32'd22211: dataIn1 = 32'd689
; 
32'd22212: dataIn1 = 32'd713
; 
32'd22213: dataIn1 = 32'd716
; 
32'd22214: dataIn1 = 32'd721
; 
32'd22215: dataIn1 = 32'd781
; 
32'd22216: dataIn1 = 32'd795
; 
32'd22217: dataIn1 = 32'd394
; 
32'd22218: dataIn1 = 32'd396
; 
32'd22219: dataIn1 = 32'd398
; 
32'd22220: dataIn1 = 32'd422
; 
32'd22221: dataIn1 = 32'd423
; 
32'd22222: dataIn1 = 32'd424
; 
32'd22223: dataIn1 = 32'd429
; 
32'd22224: dataIn1 = 32'd436
; 
32'd22225: dataIn1 = 32'd437
; 
32'd22226: dataIn1 = 32'd455
; 
32'd22227: dataIn1 = 32'd465
; 
32'd22228: dataIn1 = 32'd485
; 
32'd22229: dataIn1 = 32'd496
; 
32'd22230: dataIn1 = 32'd509
; 
32'd22231: dataIn1 = 32'd529
; 
32'd22232: dataIn1 = 32'd552
; 
32'd22233: dataIn1 = 32'd577
; 
32'd22234: dataIn1 = 32'd588
; 
32'd22235: dataIn1 = 32'd612
; 
32'd22236: dataIn1 = 32'd621
; 
32'd22237: dataIn1 = 32'd623
; 
32'd22238: dataIn1 = 32'd626
; 
32'd22239: dataIn1 = 32'd636
; 
32'd22240: dataIn1 = 32'd638
; 
32'd22241: dataIn1 = 32'd663
; 
32'd22242: dataIn1 = 32'd710
; 
32'd22243: dataIn1 = 32'd733
; 
32'd22244: dataIn1 = 32'd743
; 
32'd22245: dataIn1 = 32'd762
; 
32'd22246: dataIn1 = 32'd764
; 
32'd22247: dataIn1 = 32'd775
; 
32'd22248: dataIn1 = 32'd776
; 
32'd22249: dataIn1 = 32'd795
; 
32'd22250: dataIn1 = 32'd797
; 
32'd22251: dataIn1 = 32'd799
; 
32'd22252: dataIn1 = 32'd394
; 
32'd22253: dataIn1 = 32'd395
; 
32'd22254: dataIn1 = 32'd398
; 
32'd22255: dataIn1 = 32'd407
; 
32'd22256: dataIn1 = 32'd413
; 
32'd22257: dataIn1 = 32'd420
; 
32'd22258: dataIn1 = 32'd431
; 
32'd22259: dataIn1 = 32'd435
; 
32'd22260: dataIn1 = 32'd468
; 
32'd22261: dataIn1 = 32'd477
; 
32'd22262: dataIn1 = 32'd478
; 
32'd22263: dataIn1 = 32'd486
; 
32'd22264: dataIn1 = 32'd488
; 
32'd22265: dataIn1 = 32'd489
; 
32'd22266: dataIn1 = 32'd511
; 
32'd22267: dataIn1 = 32'd534
; 
32'd22268: dataIn1 = 32'd539
; 
32'd22269: dataIn1 = 32'd608
; 
32'd22270: dataIn1 = 32'd610
; 
32'd22271: dataIn1 = 32'd646
; 
32'd22272: dataIn1 = 32'd666
; 
32'd22273: dataIn1 = 32'd710
; 
32'd22274: dataIn1 = 32'd736
; 
32'd22275: dataIn1 = 32'd742
; 
32'd22276: dataIn1 = 32'd411
; 
32'd22277: dataIn1 = 32'd435
; 
32'd22278: dataIn1 = 32'd438
; 
32'd22279: dataIn1 = 32'd442
; 
32'd22280: dataIn1 = 32'd459
; 
32'd22281: dataIn1 = 32'd470
; 
32'd22282: dataIn1 = 32'd480
; 
32'd22283: dataIn1 = 32'd494
; 
32'd22284: dataIn1 = 32'd517
; 
32'd22285: dataIn1 = 32'd523
; 
32'd22286: dataIn1 = 32'd541
; 
32'd22287: dataIn1 = 32'd554
; 
32'd22288: dataIn1 = 32'd561
; 
32'd22289: dataIn1 = 32'd574
; 
32'd22290: dataIn1 = 32'd587
; 
32'd22291: dataIn1 = 32'd601
; 
32'd22292: dataIn1 = 32'd606
; 
32'd22293: dataIn1 = 32'd625
; 
32'd22294: dataIn1 = 32'd647
; 
32'd22295: dataIn1 = 32'd687
; 
32'd22296: dataIn1 = 32'd692
; 
32'd22297: dataIn1 = 32'd742
; 
32'd22298: dataIn1 = 32'd765
; 
32'd22299: dataIn1 = 32'd767
; 
32'd22300: dataIn1 = 32'd408
; 
32'd22301: dataIn1 = 32'd419
; 
32'd22302: dataIn1 = 32'd421
; 
32'd22303: dataIn1 = 32'd425
; 
32'd22304: dataIn1 = 32'd436
; 
32'd22305: dataIn1 = 32'd437
; 
32'd22306: dataIn1 = 32'd442
; 
32'd22307: dataIn1 = 32'd462
; 
32'd22308: dataIn1 = 32'd468
; 
32'd22309: dataIn1 = 32'd480
; 
32'd22310: dataIn1 = 32'd518
; 
32'd22311: dataIn1 = 32'd543
; 
32'd22312: dataIn1 = 32'd564
; 
32'd22313: dataIn1 = 32'd573
; 
32'd22314: dataIn1 = 32'd580
; 
32'd22315: dataIn1 = 32'd615
; 
32'd22316: dataIn1 = 32'd619
; 
32'd22317: dataIn1 = 32'd625
; 
32'd22318: dataIn1 = 32'd652
; 
32'd22319: dataIn1 = 32'd654
; 
32'd22320: dataIn1 = 32'd698
; 
32'd22321: dataIn1 = 32'd778
; 
32'd22322: dataIn1 = 32'd400
; 
32'd22323: dataIn1 = 32'd405
; 
32'd22324: dataIn1 = 32'd413
; 
32'd22325: dataIn1 = 32'd450
; 
32'd22326: dataIn1 = 32'd453
; 
32'd22327: dataIn1 = 32'd490
; 
32'd22328: dataIn1 = 32'd512
; 
32'd22329: dataIn1 = 32'd552
; 
32'd22330: dataIn1 = 32'd602
; 
32'd22331: dataIn1 = 32'd603
; 
32'd22332: dataIn1 = 32'd604
; 
32'd22333: dataIn1 = 32'd614
; 
32'd22334: dataIn1 = 32'd621
; 
32'd22335: dataIn1 = 32'd634
; 
32'd22336: dataIn1 = 32'd640
; 
32'd22337: dataIn1 = 32'd656
; 
32'd22338: dataIn1 = 32'd658
; 
32'd22339: dataIn1 = 32'd660
; 
32'd22340: dataIn1 = 32'd677
; 
32'd22341: dataIn1 = 32'd697
; 
32'd22342: dataIn1 = 32'd701
; 
32'd22343: dataIn1 = 32'd709
; 
32'd22344: dataIn1 = 32'd718
; 
32'd22345: dataIn1 = 32'd719
; 
32'd22346: dataIn1 = 32'd727
; 
32'd22347: dataIn1 = 32'd740
; 
32'd22348: dataIn1 = 32'd763
; 
32'd22349: dataIn1 = 32'd767
; 
32'd22350: dataIn1 = 32'd770
; 
32'd22351: dataIn1 = 32'd774
; 
32'd22352: dataIn1 = 32'd405
; 
32'd22353: dataIn1 = 32'd409
; 
32'd22354: dataIn1 = 32'd412
; 
32'd22355: dataIn1 = 32'd432
; 
32'd22356: dataIn1 = 32'd435
; 
32'd22357: dataIn1 = 32'd449
; 
32'd22358: dataIn1 = 32'd491
; 
32'd22359: dataIn1 = 32'd500
; 
32'd22360: dataIn1 = 32'd545
; 
32'd22361: dataIn1 = 32'd598
; 
32'd22362: dataIn1 = 32'd611
; 
32'd22363: dataIn1 = 32'd630
; 
32'd22364: dataIn1 = 32'd631
; 
32'd22365: dataIn1 = 32'd632
; 
32'd22366: dataIn1 = 32'd660
; 
32'd22367: dataIn1 = 32'd680
; 
32'd22368: dataIn1 = 32'd707
; 
32'd22369: dataIn1 = 32'd720
; 
32'd22370: dataIn1 = 32'd723
; 
32'd22371: dataIn1 = 32'd725
; 
32'd22372: dataIn1 = 32'd728
; 
32'd22373: dataIn1 = 32'd775
; 
32'd22374: dataIn1 = 32'd789
; 
32'd22375: dataIn1 = 32'd796
; 
32'd22376: dataIn1 = 32'd423
; 
32'd22377: dataIn1 = 32'd436
; 
32'd22378: dataIn1 = 32'd480
; 
32'd22379: dataIn1 = 32'd508
; 
32'd22380: dataIn1 = 32'd519
; 
32'd22381: dataIn1 = 32'd562
; 
32'd22382: dataIn1 = 32'd566
; 
32'd22383: dataIn1 = 32'd605
; 
32'd22384: dataIn1 = 32'd613
; 
32'd22385: dataIn1 = 32'd673
; 
32'd22386: dataIn1 = 32'd686
; 
32'd22387: dataIn1 = 32'd759
; 
32'd22388: dataIn1 = 32'd771
; 
32'd22389: dataIn1 = 32'd787
; 
32'd22390: dataIn1 = 32'd434
; 
32'd22391: dataIn1 = 32'd454
; 
32'd22392: dataIn1 = 32'd524
; 
32'd22393: dataIn1 = 32'd544
; 
32'd22394: dataIn1 = 32'd555
; 
32'd22395: dataIn1 = 32'd578
; 
32'd22396: dataIn1 = 32'd581
; 
32'd22397: dataIn1 = 32'd585
; 
32'd22398: dataIn1 = 32'd602
; 
32'd22399: dataIn1 = 32'd605
; 
32'd22400: dataIn1 = 32'd612
; 
32'd22401: dataIn1 = 32'd623
; 
32'd22402: dataIn1 = 32'd629
; 
32'd22403: dataIn1 = 32'd646
; 
32'd22404: dataIn1 = 32'd688
; 
32'd22405: dataIn1 = 32'd699
; 
32'd22406: dataIn1 = 32'd728
; 
32'd22407: dataIn1 = 32'd740
; 
32'd22408: dataIn1 = 32'd755
; 
32'd22409: dataIn1 = 32'd788
; 
32'd22410: dataIn1 = 32'd463
; 
32'd22411: dataIn1 = 32'd482
; 
32'd22412: dataIn1 = 32'd487
; 
32'd22413: dataIn1 = 32'd506
; 
32'd22414: dataIn1 = 32'd509
; 
32'd22415: dataIn1 = 32'd533
; 
32'd22416: dataIn1 = 32'd564
; 
32'd22417: dataIn1 = 32'd585
; 
32'd22418: dataIn1 = 32'd588
; 
32'd22419: dataIn1 = 32'd590
; 
32'd22420: dataIn1 = 32'd601
; 
32'd22421: dataIn1 = 32'd603
; 
32'd22422: dataIn1 = 32'd613
; 
32'd22423: dataIn1 = 32'd620
; 
32'd22424: dataIn1 = 32'd647
; 
32'd22425: dataIn1 = 32'd716
; 
32'd22426: dataIn1 = 32'd724
; 
32'd22427: dataIn1 = 32'd749
; 
32'd22428: dataIn1 = 32'd762
; 
32'd22429: dataIn1 = 32'd763
; 
32'd22430: dataIn1 = 32'd778
; 
32'd22431: dataIn1 = 32'd783
; 
32'd22432: dataIn1 = 32'd402
; 
32'd22433: dataIn1 = 32'd424
; 
32'd22434: dataIn1 = 32'd431
; 
32'd22435: dataIn1 = 32'd452
; 
32'd22436: dataIn1 = 32'd454
; 
32'd22437: dataIn1 = 32'd485
; 
32'd22438: dataIn1 = 32'd488
; 
32'd22439: dataIn1 = 32'd492
; 
32'd22440: dataIn1 = 32'd509
; 
32'd22441: dataIn1 = 32'd512
; 
32'd22442: dataIn1 = 32'd515
; 
32'd22443: dataIn1 = 32'd517
; 
32'd22444: dataIn1 = 32'd527
; 
32'd22445: dataIn1 = 32'd537
; 
32'd22446: dataIn1 = 32'd542
; 
32'd22447: dataIn1 = 32'd569
; 
32'd22448: dataIn1 = 32'd574
; 
32'd22449: dataIn1 = 32'd576
; 
32'd22450: dataIn1 = 32'd604
; 
32'd22451: dataIn1 = 32'd636
; 
32'd22452: dataIn1 = 32'd642
; 
32'd22453: dataIn1 = 32'd651
; 
32'd22454: dataIn1 = 32'd652
; 
32'd22455: dataIn1 = 32'd653
; 
32'd22456: dataIn1 = 32'd657
; 
32'd22457: dataIn1 = 32'd665
; 
32'd22458: dataIn1 = 32'd676
; 
32'd22459: dataIn1 = 32'd703
; 
32'd22460: dataIn1 = 32'd732
; 
32'd22461: dataIn1 = 32'd744
; 
32'd22462: dataIn1 = 32'd746
; 
32'd22463: dataIn1 = 32'd761
; 
32'd22464: dataIn1 = 32'd771
; 
32'd22465: dataIn1 = 32'd784
; 
32'd22466: dataIn1 = 32'd405
; 
32'd22467: dataIn1 = 32'd409
; 
32'd22468: dataIn1 = 32'd410
; 
32'd22469: dataIn1 = 32'd414
; 
32'd22470: dataIn1 = 32'd422
; 
32'd22471: dataIn1 = 32'd443
; 
32'd22472: dataIn1 = 32'd448
; 
32'd22473: dataIn1 = 32'd456
; 
32'd22474: dataIn1 = 32'd463
; 
32'd22475: dataIn1 = 32'd480
; 
32'd22476: dataIn1 = 32'd501
; 
32'd22477: dataIn1 = 32'd553
; 
32'd22478: dataIn1 = 32'd566
; 
32'd22479: dataIn1 = 32'd585
; 
32'd22480: dataIn1 = 32'd625
; 
32'd22481: dataIn1 = 32'd657
; 
32'd22482: dataIn1 = 32'd658
; 
32'd22483: dataIn1 = 32'd668
; 
32'd22484: dataIn1 = 32'd672
; 
32'd22485: dataIn1 = 32'd683
; 
32'd22486: dataIn1 = 32'd684
; 
32'd22487: dataIn1 = 32'd685
; 
32'd22488: dataIn1 = 32'd690
; 
32'd22489: dataIn1 = 32'd715
; 
32'd22490: dataIn1 = 32'd746
; 
32'd22491: dataIn1 = 32'd750
; 
32'd22492: dataIn1 = 32'd761
; 
32'd22493: dataIn1 = 32'd772
; 
32'd22494: dataIn1 = 32'd773
; 
32'd22495: dataIn1 = 32'd796
; 
32'd22496: dataIn1 = 32'd421
; 
32'd22497: dataIn1 = 32'd428
; 
32'd22498: dataIn1 = 32'd444
; 
32'd22499: dataIn1 = 32'd489
; 
32'd22500: dataIn1 = 32'd520
; 
32'd22501: dataIn1 = 32'd521
; 
32'd22502: dataIn1 = 32'd543
; 
32'd22503: dataIn1 = 32'd545
; 
32'd22504: dataIn1 = 32'd565
; 
32'd22505: dataIn1 = 32'd605
; 
32'd22506: dataIn1 = 32'd614
; 
32'd22507: dataIn1 = 32'd619
; 
32'd22508: dataIn1 = 32'd626
; 
32'd22509: dataIn1 = 32'd639
; 
32'd22510: dataIn1 = 32'd645
; 
32'd22511: dataIn1 = 32'd652
; 
32'd22512: dataIn1 = 32'd660
; 
32'd22513: dataIn1 = 32'd668
; 
32'd22514: dataIn1 = 32'd677
; 
32'd22515: dataIn1 = 32'd680
; 
32'd22516: dataIn1 = 32'd691
; 
32'd22517: dataIn1 = 32'd729
; 
32'd22518: dataIn1 = 32'd730
; 
32'd22519: dataIn1 = 32'd749
; 
32'd22520: dataIn1 = 32'd761
; 
32'd22521: dataIn1 = 32'd767
; 
32'd22522: dataIn1 = 32'd776
; 
32'd22523: dataIn1 = 32'd796
; 
32'd22524: dataIn1 = 32'd432
; 
32'd22525: dataIn1 = 32'd434
; 
32'd22526: dataIn1 = 32'd445
; 
32'd22527: dataIn1 = 32'd448
; 
32'd22528: dataIn1 = 32'd458
; 
32'd22529: dataIn1 = 32'd478
; 
32'd22530: dataIn1 = 32'd535
; 
32'd22531: dataIn1 = 32'd538
; 
32'd22532: dataIn1 = 32'd581
; 
32'd22533: dataIn1 = 32'd620
; 
32'd22534: dataIn1 = 32'd628
; 
32'd22535: dataIn1 = 32'd630
; 
32'd22536: dataIn1 = 32'd636
; 
32'd22537: dataIn1 = 32'd680
; 
32'd22538: dataIn1 = 32'd704
; 
32'd22539: dataIn1 = 32'd441
; 
32'd22540: dataIn1 = 32'd460
; 
32'd22541: dataIn1 = 32'd463
; 
32'd22542: dataIn1 = 32'd483
; 
32'd22543: dataIn1 = 32'd518
; 
32'd22544: dataIn1 = 32'd541
; 
32'd22545: dataIn1 = 32'd551
; 
32'd22546: dataIn1 = 32'd580
; 
32'd22547: dataIn1 = 32'd589
; 
32'd22548: dataIn1 = 32'd606
; 
32'd22549: dataIn1 = 32'd635
; 
32'd22550: dataIn1 = 32'd636
; 
32'd22551: dataIn1 = 32'd651
; 
32'd22552: dataIn1 = 32'd663
; 
32'd22553: dataIn1 = 32'd685
; 
32'd22554: dataIn1 = 32'd708
; 
32'd22555: dataIn1 = 32'd753
; 
32'd22556: dataIn1 = 32'd757
; 
32'd22557: dataIn1 = 32'd758
; 
32'd22558: dataIn1 = 32'd762
; 
32'd22559: dataIn1 = 32'd775
; 
32'd22560: dataIn1 = 32'd434
; 
32'd22561: dataIn1 = 32'd451
; 
32'd22562: dataIn1 = 32'd466
; 
32'd22563: dataIn1 = 32'd467
; 
32'd22564: dataIn1 = 32'd480
; 
32'd22565: dataIn1 = 32'd482
; 
32'd22566: dataIn1 = 32'd484
; 
32'd22567: dataIn1 = 32'd490
; 
32'd22568: dataIn1 = 32'd511
; 
32'd22569: dataIn1 = 32'd555
; 
32'd22570: dataIn1 = 32'd573
; 
32'd22571: dataIn1 = 32'd576
; 
32'd22572: dataIn1 = 32'd584
; 
32'd22573: dataIn1 = 32'd616
; 
32'd22574: dataIn1 = 32'd678
; 
32'd22575: dataIn1 = 32'd679
; 
32'd22576: dataIn1 = 32'd703
; 
32'd22577: dataIn1 = 32'd721
; 
32'd22578: dataIn1 = 32'd731
; 
32'd22579: dataIn1 = 32'd753
; 
32'd22580: dataIn1 = 32'd761
; 
32'd22581: dataIn1 = 32'd785
; 
32'd22582: dataIn1 = 32'd795
; 
32'd22583: dataIn1 = 32'd411
; 
32'd22584: dataIn1 = 32'd422
; 
32'd22585: dataIn1 = 32'd425
; 
32'd22586: dataIn1 = 32'd476
; 
32'd22587: dataIn1 = 32'd495
; 
32'd22588: dataIn1 = 32'd512
; 
32'd22589: dataIn1 = 32'd532
; 
32'd22590: dataIn1 = 32'd536
; 
32'd22591: dataIn1 = 32'd543
; 
32'd22592: dataIn1 = 32'd547
; 
32'd22593: dataIn1 = 32'd552
; 
32'd22594: dataIn1 = 32'd555
; 
32'd22595: dataIn1 = 32'd588
; 
32'd22596: dataIn1 = 32'd593
; 
32'd22597: dataIn1 = 32'd596
; 
32'd22598: dataIn1 = 32'd601
; 
32'd22599: dataIn1 = 32'd617
; 
32'd22600: dataIn1 = 32'd618
; 
32'd22601: dataIn1 = 32'd630
; 
32'd22602: dataIn1 = 32'd634
; 
32'd22603: dataIn1 = 32'd670
; 
32'd22604: dataIn1 = 32'd691
; 
32'd22605: dataIn1 = 32'd697
; 
32'd22606: dataIn1 = 32'd705
; 
32'd22607: dataIn1 = 32'd727
; 
32'd22608: dataIn1 = 32'd746
; 
32'd22609: dataIn1 = 32'd761
; 
32'd22610: dataIn1 = 32'd774
; 
32'd22611: dataIn1 = 32'd423
; 
32'd22612: dataIn1 = 32'd504
; 
32'd22613: dataIn1 = 32'd532
; 
32'd22614: dataIn1 = 32'd547
; 
32'd22615: dataIn1 = 32'd551
; 
32'd22616: dataIn1 = 32'd552
; 
32'd22617: dataIn1 = 32'd553
; 
32'd22618: dataIn1 = 32'd571
; 
32'd22619: dataIn1 = 32'd577
; 
32'd22620: dataIn1 = 32'd603
; 
32'd22621: dataIn1 = 32'd633
; 
32'd22622: dataIn1 = 32'd644
; 
32'd22623: dataIn1 = 32'd656
; 
32'd22624: dataIn1 = 32'd672
; 
32'd22625: dataIn1 = 32'd703
; 
32'd22626: dataIn1 = 32'd719
; 
32'd22627: dataIn1 = 32'd731
; 
32'd22628: dataIn1 = 32'd749
; 
32'd22629: dataIn1 = 32'd754
; 
32'd22630: dataIn1 = 32'd755
; 
32'd22631: dataIn1 = 32'd764
; 
32'd22632: dataIn1 = 32'd769
; 
32'd22633: dataIn1 = 32'd782
; 
32'd22634: dataIn1 = 32'd412
; 
32'd22635: dataIn1 = 32'd433
; 
32'd22636: dataIn1 = 32'd444
; 
32'd22637: dataIn1 = 32'd450
; 
32'd22638: dataIn1 = 32'd455
; 
32'd22639: dataIn1 = 32'd457
; 
32'd22640: dataIn1 = 32'd465
; 
32'd22641: dataIn1 = 32'd518
; 
32'd22642: dataIn1 = 32'd524
; 
32'd22643: dataIn1 = 32'd530
; 
32'd22644: dataIn1 = 32'd531
; 
32'd22645: dataIn1 = 32'd537
; 
32'd22646: dataIn1 = 32'd541
; 
32'd22647: dataIn1 = 32'd568
; 
32'd22648: dataIn1 = 32'd575
; 
32'd22649: dataIn1 = 32'd616
; 
32'd22650: dataIn1 = 32'd638
; 
32'd22651: dataIn1 = 32'd651
; 
32'd22652: dataIn1 = 32'd660
; 
32'd22653: dataIn1 = 32'd661
; 
32'd22654: dataIn1 = 32'd690
; 
32'd22655: dataIn1 = 32'd695
; 
32'd22656: dataIn1 = 32'd758
; 
32'd22657: dataIn1 = 32'd782
; 
32'd22658: dataIn1 = 32'd798
; 
32'd22659: dataIn1 = 32'd799
; 
32'd22660: dataIn1 = 32'd426
; 
32'd22661: dataIn1 = 32'd435
; 
32'd22662: dataIn1 = 32'd456
; 
32'd22663: dataIn1 = 32'd460
; 
32'd22664: dataIn1 = 32'd489
; 
32'd22665: dataIn1 = 32'd491
; 
32'd22666: dataIn1 = 32'd492
; 
32'd22667: dataIn1 = 32'd500
; 
32'd22668: dataIn1 = 32'd543
; 
32'd22669: dataIn1 = 32'd568
; 
32'd22670: dataIn1 = 32'd574
; 
32'd22671: dataIn1 = 32'd577
; 
32'd22672: dataIn1 = 32'd638
; 
32'd22673: dataIn1 = 32'd677
; 
32'd22674: dataIn1 = 32'd678
; 
32'd22675: dataIn1 = 32'd681
; 
32'd22676: dataIn1 = 32'd688
; 
32'd22677: dataIn1 = 32'd697
; 
32'd22678: dataIn1 = 32'd705
; 
32'd22679: dataIn1 = 32'd726
; 
32'd22680: dataIn1 = 32'd756
; 
32'd22681: dataIn1 = 32'd770
; 
32'd22682: dataIn1 = 32'd792
; 
32'd22683: dataIn1 = 32'd799
; 
32'd22684: dataIn1 = 32'd412
; 
32'd22685: dataIn1 = 32'd455
; 
32'd22686: dataIn1 = 32'd475
; 
32'd22687: dataIn1 = 32'd476
; 
32'd22688: dataIn1 = 32'd479
; 
32'd22689: dataIn1 = 32'd482
; 
32'd22690: dataIn1 = 32'd528
; 
32'd22691: dataIn1 = 32'd554
; 
32'd22692: dataIn1 = 32'd571
; 
32'd22693: dataIn1 = 32'd591
; 
32'd22694: dataIn1 = 32'd606
; 
32'd22695: dataIn1 = 32'd620
; 
32'd22696: dataIn1 = 32'd654
; 
32'd22697: dataIn1 = 32'd670
; 
32'd22698: dataIn1 = 32'd672
; 
32'd22699: dataIn1 = 32'd720
; 
32'd22700: dataIn1 = 32'd753
; 
32'd22701: dataIn1 = 32'd777
; 
32'd22702: dataIn1 = 32'd785
; 
32'd22703: dataIn1 = 32'd789
; 
32'd22704: dataIn1 = 32'd795
; 
32'd22705: dataIn1 = 32'd798
; 
32'd22706: dataIn1 = 32'd443
; 
32'd22707: dataIn1 = 32'd444
; 
32'd22708: dataIn1 = 32'd448
; 
32'd22709: dataIn1 = 32'd459
; 
32'd22710: dataIn1 = 32'd482
; 
32'd22711: dataIn1 = 32'd499
; 
32'd22712: dataIn1 = 32'd501
; 
32'd22713: dataIn1 = 32'd506
; 
32'd22714: dataIn1 = 32'd516
; 
32'd22715: dataIn1 = 32'd522
; 
32'd22716: dataIn1 = 32'd532
; 
32'd22717: dataIn1 = 32'd533
; 
32'd22718: dataIn1 = 32'd545
; 
32'd22719: dataIn1 = 32'd548
; 
32'd22720: dataIn1 = 32'd586
; 
32'd22721: dataIn1 = 32'd610
; 
32'd22722: dataIn1 = 32'd632
; 
32'd22723: dataIn1 = 32'd638
; 
32'd22724: dataIn1 = 32'd642
; 
32'd22725: dataIn1 = 32'd663
; 
32'd22726: dataIn1 = 32'd689
; 
32'd22727: dataIn1 = 32'd706
; 
32'd22728: dataIn1 = 32'd726
; 
32'd22729: dataIn1 = 32'd755
; 
32'd22730: dataIn1 = 32'd772
; 
32'd22731: dataIn1 = 32'd773
; 
32'd22732: dataIn1 = 32'd455
; 
32'd22733: dataIn1 = 32'd464
; 
32'd22734: dataIn1 = 32'd467
; 
32'd22735: dataIn1 = 32'd490
; 
32'd22736: dataIn1 = 32'd503
; 
32'd22737: dataIn1 = 32'd519
; 
32'd22738: dataIn1 = 32'd522
; 
32'd22739: dataIn1 = 32'd530
; 
32'd22740: dataIn1 = 32'd533
; 
32'd22741: dataIn1 = 32'd535
; 
32'd22742: dataIn1 = 32'd558
; 
32'd22743: dataIn1 = 32'd607
; 
32'd22744: dataIn1 = 32'd616
; 
32'd22745: dataIn1 = 32'd643
; 
32'd22746: dataIn1 = 32'd665
; 
32'd22747: dataIn1 = 32'd667
; 
32'd22748: dataIn1 = 32'd673
; 
32'd22749: dataIn1 = 32'd717
; 
32'd22750: dataIn1 = 32'd726
; 
32'd22751: dataIn1 = 32'd784
; 
32'd22752: dataIn1 = 32'd799
; 
32'd22753: dataIn1 = 32'd800
; 
32'd22754: dataIn1 = 32'd416
; 
32'd22755: dataIn1 = 32'd456
; 
32'd22756: dataIn1 = 32'd477
; 
32'd22757: dataIn1 = 32'd503
; 
32'd22758: dataIn1 = 32'd511
; 
32'd22759: dataIn1 = 32'd519
; 
32'd22760: dataIn1 = 32'd529
; 
32'd22761: dataIn1 = 32'd677
; 
32'd22762: dataIn1 = 32'd687
; 
32'd22763: dataIn1 = 32'd715
; 
32'd22764: dataIn1 = 32'd722
; 
32'd22765: dataIn1 = 32'd723
; 
32'd22766: dataIn1 = 32'd748
; 
32'd22767: dataIn1 = 32'd750
; 
32'd22768: dataIn1 = 32'd751
; 
32'd22769: dataIn1 = 32'd768
; 
32'd22770: dataIn1 = 32'd416
; 
32'd22771: dataIn1 = 32'd421
; 
32'd22772: dataIn1 = 32'd425
; 
32'd22773: dataIn1 = 32'd453
; 
32'd22774: dataIn1 = 32'd501
; 
32'd22775: dataIn1 = 32'd523
; 
32'd22776: dataIn1 = 32'd532
; 
32'd22777: dataIn1 = 32'd534
; 
32'd22778: dataIn1 = 32'd552
; 
32'd22779: dataIn1 = 32'd561
; 
32'd22780: dataIn1 = 32'd579
; 
32'd22781: dataIn1 = 32'd629
; 
32'd22782: dataIn1 = 32'd648
; 
32'd22783: dataIn1 = 32'd668
; 
32'd22784: dataIn1 = 32'd673
; 
32'd22785: dataIn1 = 32'd680
; 
32'd22786: dataIn1 = 32'd682
; 
32'd22787: dataIn1 = 32'd686
; 
32'd22788: dataIn1 = 32'd690
; 
32'd22789: dataIn1 = 32'd709
; 
32'd22790: dataIn1 = 32'd715
; 
32'd22791: dataIn1 = 32'd733
; 
32'd22792: dataIn1 = 32'd741
; 
32'd22793: dataIn1 = 32'd750
; 
32'd22794: dataIn1 = 32'd757
; 
32'd22795: dataIn1 = 32'd769
; 
32'd22796: dataIn1 = 32'd777
; 
32'd22797: dataIn1 = 32'd793
; 
32'd22798: dataIn1 = 32'd800
; 
32'd22799: dataIn1 = 32'd419
; 
32'd22800: dataIn1 = 32'd421
; 
32'd22801: dataIn1 = 32'd459
; 
32'd22802: dataIn1 = 32'd486
; 
32'd22803: dataIn1 = 32'd487
; 
32'd22804: dataIn1 = 32'd507
; 
32'd22805: dataIn1 = 32'd514
; 
32'd22806: dataIn1 = 32'd538
; 
32'd22807: dataIn1 = 32'd539
; 
32'd22808: dataIn1 = 32'd558
; 
32'd22809: dataIn1 = 32'd564
; 
32'd22810: dataIn1 = 32'd576
; 
32'd22811: dataIn1 = 32'd610
; 
32'd22812: dataIn1 = 32'd612
; 
32'd22813: dataIn1 = 32'd662
; 
32'd22814: dataIn1 = 32'd687
; 
32'd22815: dataIn1 = 32'd419
; 
32'd22816: dataIn1 = 32'd431
; 
32'd22817: dataIn1 = 32'd435
; 
32'd22818: dataIn1 = 32'd446
; 
32'd22819: dataIn1 = 32'd453
; 
32'd22820: dataIn1 = 32'd458
; 
32'd22821: dataIn1 = 32'd463
; 
32'd22822: dataIn1 = 32'd469
; 
32'd22823: dataIn1 = 32'd485
; 
32'd22824: dataIn1 = 32'd500
; 
32'd22825: dataIn1 = 32'd504
; 
32'd22826: dataIn1 = 32'd512
; 
32'd22827: dataIn1 = 32'd538
; 
32'd22828: dataIn1 = 32'd541
; 
32'd22829: dataIn1 = 32'd561
; 
32'd22830: dataIn1 = 32'd568
; 
32'd22831: dataIn1 = 32'd574
; 
32'd22832: dataIn1 = 32'd612
; 
32'd22833: dataIn1 = 32'd613
; 
32'd22834: dataIn1 = 32'd636
; 
32'd22835: dataIn1 = 32'd658
; 
32'd22836: dataIn1 = 32'd703
; 
32'd22837: dataIn1 = 32'd707
; 
32'd22838: dataIn1 = 32'd746
; 
32'd22839: dataIn1 = 32'd758
; 
32'd22840: dataIn1 = 32'd768
; 
32'd22841: dataIn1 = 32'd777
; 
32'd22842: dataIn1 = 32'd791
; 
32'd22843: dataIn1 = 32'd420
; 
32'd22844: dataIn1 = 32'd421
; 
32'd22845: dataIn1 = 32'd430
; 
32'd22846: dataIn1 = 32'd432
; 
32'd22847: dataIn1 = 32'd449
; 
32'd22848: dataIn1 = 32'd459
; 
32'd22849: dataIn1 = 32'd468
; 
32'd22850: dataIn1 = 32'd483
; 
32'd22851: dataIn1 = 32'd501
; 
32'd22852: dataIn1 = 32'd519
; 
32'd22853: dataIn1 = 32'd542
; 
32'd22854: dataIn1 = 32'd555
; 
32'd22855: dataIn1 = 32'd556
; 
32'd22856: dataIn1 = 32'd558
; 
32'd22857: dataIn1 = 32'd571
; 
32'd22858: dataIn1 = 32'd604
; 
32'd22859: dataIn1 = 32'd606
; 
32'd22860: dataIn1 = 32'd613
; 
32'd22861: dataIn1 = 32'd627
; 
32'd22862: dataIn1 = 32'd650
; 
32'd22863: dataIn1 = 32'd652
; 
32'd22864: dataIn1 = 32'd655
; 
32'd22865: dataIn1 = 32'd659
; 
32'd22866: dataIn1 = 32'd660
; 
32'd22867: dataIn1 = 32'd689
; 
32'd22868: dataIn1 = 32'd698
; 
32'd22869: dataIn1 = 32'd703
; 
32'd22870: dataIn1 = 32'd709
; 
32'd22871: dataIn1 = 32'd734
; 
32'd22872: dataIn1 = 32'd747
; 
32'd22873: dataIn1 = 32'd752
; 
32'd22874: dataIn1 = 32'd760
; 
32'd22875: dataIn1 = 32'd764
; 
32'd22876: dataIn1 = 32'd789
; 
32'd22877: dataIn1 = 32'd799
; 
32'd22878: dataIn1 = 32'd800
; 
32'd22879: dataIn1 = 32'd424
; 
32'd22880: dataIn1 = 32'd445
; 
32'd22881: dataIn1 = 32'd456
; 
32'd22882: dataIn1 = 32'd471
; 
32'd22883: dataIn1 = 32'd508
; 
32'd22884: dataIn1 = 32'd560
; 
32'd22885: dataIn1 = 32'd568
; 
32'd22886: dataIn1 = 32'd595
; 
32'd22887: dataIn1 = 32'd644
; 
32'd22888: dataIn1 = 32'd670
; 
32'd22889: dataIn1 = 32'd672
; 
32'd22890: dataIn1 = 32'd700
; 
32'd22891: dataIn1 = 32'd716
; 
32'd22892: dataIn1 = 32'd723
; 
32'd22893: dataIn1 = 32'd759
; 
32'd22894: dataIn1 = 32'd770
; 
32'd22895: dataIn1 = 32'd440
; 
32'd22896: dataIn1 = 32'd478
; 
32'd22897: dataIn1 = 32'd484
; 
32'd22898: dataIn1 = 32'd487
; 
32'd22899: dataIn1 = 32'd506
; 
32'd22900: dataIn1 = 32'd513
; 
32'd22901: dataIn1 = 32'd544
; 
32'd22902: dataIn1 = 32'd546
; 
32'd22903: dataIn1 = 32'd579
; 
32'd22904: dataIn1 = 32'd607
; 
32'd22905: dataIn1 = 32'd609
; 
32'd22906: dataIn1 = 32'd627
; 
32'd22907: dataIn1 = 32'd662
; 
32'd22908: dataIn1 = 32'd663
; 
32'd22909: dataIn1 = 32'd664
; 
32'd22910: dataIn1 = 32'd730
; 
32'd22911: dataIn1 = 32'd732
; 
32'd22912: dataIn1 = 32'd751
; 
32'd22913: dataIn1 = 32'd433
; 
32'd22914: dataIn1 = 32'd442
; 
32'd22915: dataIn1 = 32'd445
; 
32'd22916: dataIn1 = 32'd454
; 
32'd22917: dataIn1 = 32'd459
; 
32'd22918: dataIn1 = 32'd464
; 
32'd22919: dataIn1 = 32'd468
; 
32'd22920: dataIn1 = 32'd481
; 
32'd22921: dataIn1 = 32'd499
; 
32'd22922: dataIn1 = 32'd506
; 
32'd22923: dataIn1 = 32'd517
; 
32'd22924: dataIn1 = 32'd519
; 
32'd22925: dataIn1 = 32'd541
; 
32'd22926: dataIn1 = 32'd543
; 
32'd22927: dataIn1 = 32'd546
; 
32'd22928: dataIn1 = 32'd549
; 
32'd22929: dataIn1 = 32'd560
; 
32'd22930: dataIn1 = 32'd588
; 
32'd22931: dataIn1 = 32'd608
; 
32'd22932: dataIn1 = 32'd620
; 
32'd22933: dataIn1 = 32'd624
; 
32'd22934: dataIn1 = 32'd636
; 
32'd22935: dataIn1 = 32'd674
; 
32'd22936: dataIn1 = 32'd685
; 
32'd22937: dataIn1 = 32'd686
; 
32'd22938: dataIn1 = 32'd687
; 
32'd22939: dataIn1 = 32'd688
; 
32'd22940: dataIn1 = 32'd727
; 
32'd22941: dataIn1 = 32'd737
; 
32'd22942: dataIn1 = 32'd744
; 
32'd22943: dataIn1 = 32'd747
; 
32'd22944: dataIn1 = 32'd755
; 
32'd22945: dataIn1 = 32'd778
; 
32'd22946: dataIn1 = 32'd466
; 
32'd22947: dataIn1 = 32'd492
; 
32'd22948: dataIn1 = 32'd541
; 
32'd22949: dataIn1 = 32'd590
; 
32'd22950: dataIn1 = 32'd597
; 
32'd22951: dataIn1 = 32'd613
; 
32'd22952: dataIn1 = 32'd614
; 
32'd22953: dataIn1 = 32'd629
; 
32'd22954: dataIn1 = 32'd640
; 
32'd22955: dataIn1 = 32'd644
; 
32'd22956: dataIn1 = 32'd701
; 
32'd22957: dataIn1 = 32'd702
; 
32'd22958: dataIn1 = 32'd738
; 
32'd22959: dataIn1 = 32'd742
; 
32'd22960: dataIn1 = 32'd765
; 
32'd22961: dataIn1 = 32'd770
; 
32'd22962: dataIn1 = 32'd772
; 
32'd22963: dataIn1 = 32'd794
; 
32'd22964: dataIn1 = 32'd431
; 
32'd22965: dataIn1 = 32'd499
; 
32'd22966: dataIn1 = 32'd515
; 
32'd22967: dataIn1 = 32'd522
; 
32'd22968: dataIn1 = 32'd537
; 
32'd22969: dataIn1 = 32'd539
; 
32'd22970: dataIn1 = 32'd561
; 
32'd22971: dataIn1 = 32'd567
; 
32'd22972: dataIn1 = 32'd577
; 
32'd22973: dataIn1 = 32'd599
; 
32'd22974: dataIn1 = 32'd647
; 
32'd22975: dataIn1 = 32'd657
; 
32'd22976: dataIn1 = 32'd672
; 
32'd22977: dataIn1 = 32'd679
; 
32'd22978: dataIn1 = 32'd695
; 
32'd22979: dataIn1 = 32'd754
; 
32'd22980: dataIn1 = 32'd775
; 
32'd22981: dataIn1 = 32'd776
; 
32'd22982: dataIn1 = 32'd777
; 
32'd22983: dataIn1 = 32'd799
; 
32'd22984: dataIn1 = 32'd434
; 
32'd22985: dataIn1 = 32'd454
; 
32'd22986: dataIn1 = 32'd456
; 
32'd22987: dataIn1 = 32'd464
; 
32'd22988: dataIn1 = 32'd470
; 
32'd22989: dataIn1 = 32'd472
; 
32'd22990: dataIn1 = 32'd490
; 
32'd22991: dataIn1 = 32'd509
; 
32'd22992: dataIn1 = 32'd528
; 
32'd22993: dataIn1 = 32'd556
; 
32'd22994: dataIn1 = 32'd558
; 
32'd22995: dataIn1 = 32'd609
; 
32'd22996: dataIn1 = 32'd620
; 
32'd22997: dataIn1 = 32'd624
; 
32'd22998: dataIn1 = 32'd711
; 
32'd22999: dataIn1 = 32'd720
; 
32'd23000: dataIn1 = 32'd733
; 
32'd23001: dataIn1 = 32'd768
; 
32'd23002: dataIn1 = 32'd789
; 
32'd23003: dataIn1 = 32'd475
; 
32'd23004: dataIn1 = 32'd509
; 
32'd23005: dataIn1 = 32'd517
; 
32'd23006: dataIn1 = 32'd527
; 
32'd23007: dataIn1 = 32'd530
; 
32'd23008: dataIn1 = 32'd571
; 
32'd23009: dataIn1 = 32'd573
; 
32'd23010: dataIn1 = 32'd575
; 
32'd23011: dataIn1 = 32'd577
; 
32'd23012: dataIn1 = 32'd585
; 
32'd23013: dataIn1 = 32'd642
; 
32'd23014: dataIn1 = 32'd690
; 
32'd23015: dataIn1 = 32'd701
; 
32'd23016: dataIn1 = 32'd706
; 
32'd23017: dataIn1 = 32'd754
; 
32'd23018: dataIn1 = 32'd757
; 
32'd23019: dataIn1 = 32'd773
; 
32'd23020: dataIn1 = 32'd774
; 
32'd23021: dataIn1 = 32'd778
; 
32'd23022: dataIn1 = 32'd783
; 
32'd23023: dataIn1 = 32'd795
; 
32'd23024: dataIn1 = 32'd800
; 
32'd23025: dataIn1 = 32'd434
; 
32'd23026: dataIn1 = 32'd448
; 
32'd23027: dataIn1 = 32'd454
; 
32'd23028: dataIn1 = 32'd455
; 
32'd23029: dataIn1 = 32'd461
; 
32'd23030: dataIn1 = 32'd464
; 
32'd23031: dataIn1 = 32'd477
; 
32'd23032: dataIn1 = 32'd480
; 
32'd23033: dataIn1 = 32'd481
; 
32'd23034: dataIn1 = 32'd515
; 
32'd23035: dataIn1 = 32'd524
; 
32'd23036: dataIn1 = 32'd566
; 
32'd23037: dataIn1 = 32'd614
; 
32'd23038: dataIn1 = 32'd666
; 
32'd23039: dataIn1 = 32'd675
; 
32'd23040: dataIn1 = 32'd681
; 
32'd23041: dataIn1 = 32'd697
; 
32'd23042: dataIn1 = 32'd718
; 
32'd23043: dataIn1 = 32'd746
; 
32'd23044: dataIn1 = 32'd758
; 
32'd23045: dataIn1 = 32'd766
; 
32'd23046: dataIn1 = 32'd770
; 
32'd23047: dataIn1 = 32'd772
; 
32'd23048: dataIn1 = 32'd775
; 
32'd23049: dataIn1 = 32'd778
; 
32'd23050: dataIn1 = 32'd448
; 
32'd23051: dataIn1 = 32'd472
; 
32'd23052: dataIn1 = 32'd496
; 
32'd23053: dataIn1 = 32'd501
; 
32'd23054: dataIn1 = 32'd526
; 
32'd23055: dataIn1 = 32'd541
; 
32'd23056: dataIn1 = 32'd566
; 
32'd23057: dataIn1 = 32'd573
; 
32'd23058: dataIn1 = 32'd590
; 
32'd23059: dataIn1 = 32'd591
; 
32'd23060: dataIn1 = 32'd610
; 
32'd23061: dataIn1 = 32'd618
; 
32'd23062: dataIn1 = 32'd621
; 
32'd23063: dataIn1 = 32'd627
; 
32'd23064: dataIn1 = 32'd640
; 
32'd23065: dataIn1 = 32'd668
; 
32'd23066: dataIn1 = 32'd674
; 
32'd23067: dataIn1 = 32'd675
; 
32'd23068: dataIn1 = 32'd683
; 
32'd23069: dataIn1 = 32'd694
; 
32'd23070: dataIn1 = 32'd701
; 
32'd23071: dataIn1 = 32'd703
; 
32'd23072: dataIn1 = 32'd732
; 
32'd23073: dataIn1 = 32'd763
; 
32'd23074: dataIn1 = 32'd773
; 
32'd23075: dataIn1 = 32'd796
; 
32'd23076: dataIn1 = 32'd437
; 
32'd23077: dataIn1 = 32'd454
; 
32'd23078: dataIn1 = 32'd467
; 
32'd23079: dataIn1 = 32'd479
; 
32'd23080: dataIn1 = 32'd500
; 
32'd23081: dataIn1 = 32'd519
; 
32'd23082: dataIn1 = 32'd526
; 
32'd23083: dataIn1 = 32'd550
; 
32'd23084: dataIn1 = 32'd576
; 
32'd23085: dataIn1 = 32'd595
; 
32'd23086: dataIn1 = 32'd611
; 
32'd23087: dataIn1 = 32'd632
; 
32'd23088: dataIn1 = 32'd645
; 
32'd23089: dataIn1 = 32'd649
; 
32'd23090: dataIn1 = 32'd656
; 
32'd23091: dataIn1 = 32'd719
; 
32'd23092: dataIn1 = 32'd723
; 
32'd23093: dataIn1 = 32'd736
; 
32'd23094: dataIn1 = 32'd751
; 
32'd23095: dataIn1 = 32'd761
; 
32'd23096: dataIn1 = 32'd770
; 
32'd23097: dataIn1 = 32'd786
; 
32'd23098: dataIn1 = 32'd791
; 
32'd23099: dataIn1 = 32'd449
; 
32'd23100: dataIn1 = 32'd456
; 
32'd23101: dataIn1 = 32'd467
; 
32'd23102: dataIn1 = 32'd475
; 
32'd23103: dataIn1 = 32'd494
; 
32'd23104: dataIn1 = 32'd508
; 
32'd23105: dataIn1 = 32'd512
; 
32'd23106: dataIn1 = 32'd581
; 
32'd23107: dataIn1 = 32'd606
; 
32'd23108: dataIn1 = 32'd623
; 
32'd23109: dataIn1 = 32'd638
; 
32'd23110: dataIn1 = 32'd660
; 
32'd23111: dataIn1 = 32'd662
; 
32'd23112: dataIn1 = 32'd678
; 
32'd23113: dataIn1 = 32'd679
; 
32'd23114: dataIn1 = 32'd721
; 
32'd23115: dataIn1 = 32'd723
; 
32'd23116: dataIn1 = 32'd762
; 
32'd23117: dataIn1 = 32'd782
; 
32'd23118: dataIn1 = 32'd786
; 
32'd23119: dataIn1 = 32'd462
; 
32'd23120: dataIn1 = 32'd477
; 
32'd23121: dataIn1 = 32'd480
; 
32'd23122: dataIn1 = 32'd483
; 
32'd23123: dataIn1 = 32'd526
; 
32'd23124: dataIn1 = 32'd529
; 
32'd23125: dataIn1 = 32'd536
; 
32'd23126: dataIn1 = 32'd568
; 
32'd23127: dataIn1 = 32'd574
; 
32'd23128: dataIn1 = 32'd611
; 
32'd23129: dataIn1 = 32'd645
; 
32'd23130: dataIn1 = 32'd661
; 
32'd23131: dataIn1 = 32'd691
; 
32'd23132: dataIn1 = 32'd700
; 
32'd23133: dataIn1 = 32'd723
; 
32'd23134: dataIn1 = 32'd757
; 
32'd23135: dataIn1 = 32'd780
; 
32'd23136: dataIn1 = 32'd437
; 
32'd23137: dataIn1 = 32'd443
; 
32'd23138: dataIn1 = 32'd447
; 
32'd23139: dataIn1 = 32'd449
; 
32'd23140: dataIn1 = 32'd458
; 
32'd23141: dataIn1 = 32'd466
; 
32'd23142: dataIn1 = 32'd478
; 
32'd23143: dataIn1 = 32'd523
; 
32'd23144: dataIn1 = 32'd537
; 
32'd23145: dataIn1 = 32'd539
; 
32'd23146: dataIn1 = 32'd586
; 
32'd23147: dataIn1 = 32'd588
; 
32'd23148: dataIn1 = 32'd630
; 
32'd23149: dataIn1 = 32'd631
; 
32'd23150: dataIn1 = 32'd684
; 
32'd23151: dataIn1 = 32'd693
; 
32'd23152: dataIn1 = 32'd713
; 
32'd23153: dataIn1 = 32'd728
; 
32'd23154: dataIn1 = 32'd740
; 
32'd23155: dataIn1 = 32'd759
; 
32'd23156: dataIn1 = 32'd784
; 
32'd23157: dataIn1 = 32'd788
; 
32'd23158: dataIn1 = 32'd799
; 
32'd23159: dataIn1 = 32'd433
; 
32'd23160: dataIn1 = 32'd436
; 
32'd23161: dataIn1 = 32'd463
; 
32'd23162: dataIn1 = 32'd504
; 
32'd23163: dataIn1 = 32'd522
; 
32'd23164: dataIn1 = 32'd575
; 
32'd23165: dataIn1 = 32'd581
; 
32'd23166: dataIn1 = 32'd601
; 
32'd23167: dataIn1 = 32'd610
; 
32'd23168: dataIn1 = 32'd657
; 
32'd23169: dataIn1 = 32'd666
; 
32'd23170: dataIn1 = 32'd677
; 
32'd23171: dataIn1 = 32'd680
; 
32'd23172: dataIn1 = 32'd699
; 
32'd23173: dataIn1 = 32'd701
; 
32'd23174: dataIn1 = 32'd704
; 
32'd23175: dataIn1 = 32'd727
; 
32'd23176: dataIn1 = 32'd748
; 
32'd23177: dataIn1 = 32'd764
; 
32'd23178: dataIn1 = 32'd434
; 
32'd23179: dataIn1 = 32'd448
; 
32'd23180: dataIn1 = 32'd532
; 
32'd23181: dataIn1 = 32'd535
; 
32'd23182: dataIn1 = 32'd559
; 
32'd23183: dataIn1 = 32'd570
; 
32'd23184: dataIn1 = 32'd579
; 
32'd23185: dataIn1 = 32'd608
; 
32'd23186: dataIn1 = 32'd627
; 
32'd23187: dataIn1 = 32'd651
; 
32'd23188: dataIn1 = 32'd664
; 
32'd23189: dataIn1 = 32'd727
; 
32'd23190: dataIn1 = 32'd740
; 
32'd23191: dataIn1 = 32'd745
; 
32'd23192: dataIn1 = 32'd747
; 
32'd23193: dataIn1 = 32'd753
; 
32'd23194: dataIn1 = 32'd459
; 
32'd23195: dataIn1 = 32'd462
; 
32'd23196: dataIn1 = 32'd495
; 
32'd23197: dataIn1 = 32'd523
; 
32'd23198: dataIn1 = 32'd531
; 
32'd23199: dataIn1 = 32'd547
; 
32'd23200: dataIn1 = 32'd551
; 
32'd23201: dataIn1 = 32'd590
; 
32'd23202: dataIn1 = 32'd607
; 
32'd23203: dataIn1 = 32'd621
; 
32'd23204: dataIn1 = 32'd643
; 
32'd23205: dataIn1 = 32'd655
; 
32'd23206: dataIn1 = 32'd656
; 
32'd23207: dataIn1 = 32'd661
; 
32'd23208: dataIn1 = 32'd670
; 
32'd23209: dataIn1 = 32'd676
; 
32'd23210: dataIn1 = 32'd691
; 
32'd23211: dataIn1 = 32'd710
; 
32'd23212: dataIn1 = 32'd716
; 
32'd23213: dataIn1 = 32'd727
; 
32'd23214: dataIn1 = 32'd734
; 
32'd23215: dataIn1 = 32'd739
; 
32'd23216: dataIn1 = 32'd770
; 
32'd23217: dataIn1 = 32'd793
; 
32'd23218: dataIn1 = 32'd443
; 
32'd23219: dataIn1 = 32'd477
; 
32'd23220: dataIn1 = 32'd533
; 
32'd23221: dataIn1 = 32'd542
; 
32'd23222: dataIn1 = 32'd555
; 
32'd23223: dataIn1 = 32'd557
; 
32'd23224: dataIn1 = 32'd561
; 
32'd23225: dataIn1 = 32'd587
; 
32'd23226: dataIn1 = 32'd610
; 
32'd23227: dataIn1 = 32'd611
; 
32'd23228: dataIn1 = 32'd621
; 
32'd23229: dataIn1 = 32'd622
; 
32'd23230: dataIn1 = 32'd650
; 
32'd23231: dataIn1 = 32'd653
; 
32'd23232: dataIn1 = 32'd654
; 
32'd23233: dataIn1 = 32'd673
; 
32'd23234: dataIn1 = 32'd698
; 
32'd23235: dataIn1 = 32'd759
; 
32'd23236: dataIn1 = 32'd766
; 
32'd23237: dataIn1 = 32'd794
; 
32'd23238: dataIn1 = 32'd799
; 
32'd23239: dataIn1 = 32'd443
; 
32'd23240: dataIn1 = 32'd455
; 
32'd23241: dataIn1 = 32'd463
; 
32'd23242: dataIn1 = 32'd465
; 
32'd23243: dataIn1 = 32'd478
; 
32'd23244: dataIn1 = 32'd479
; 
32'd23245: dataIn1 = 32'd495
; 
32'd23246: dataIn1 = 32'd523
; 
32'd23247: dataIn1 = 32'd534
; 
32'd23248: dataIn1 = 32'd545
; 
32'd23249: dataIn1 = 32'd563
; 
32'd23250: dataIn1 = 32'd574
; 
32'd23251: dataIn1 = 32'd576
; 
32'd23252: dataIn1 = 32'd610
; 
32'd23253: dataIn1 = 32'd615
; 
32'd23254: dataIn1 = 32'd616
; 
32'd23255: dataIn1 = 32'd649
; 
32'd23256: dataIn1 = 32'd650
; 
32'd23257: dataIn1 = 32'd656
; 
32'd23258: dataIn1 = 32'd668
; 
32'd23259: dataIn1 = 32'd681
; 
32'd23260: dataIn1 = 32'd691
; 
32'd23261: dataIn1 = 32'd709
; 
32'd23262: dataIn1 = 32'd768
; 
32'd23263: dataIn1 = 32'd772
; 
32'd23264: dataIn1 = 32'd773
; 
32'd23265: dataIn1 = 32'd777
; 
32'd23266: dataIn1 = 32'd441
; 
32'd23267: dataIn1 = 32'd446
; 
32'd23268: dataIn1 = 32'd470
; 
32'd23269: dataIn1 = 32'd496
; 
32'd23270: dataIn1 = 32'd513
; 
32'd23271: dataIn1 = 32'd517
; 
32'd23272: dataIn1 = 32'd524
; 
32'd23273: dataIn1 = 32'd538
; 
32'd23274: dataIn1 = 32'd552
; 
32'd23275: dataIn1 = 32'd556
; 
32'd23276: dataIn1 = 32'd580
; 
32'd23277: dataIn1 = 32'd581
; 
32'd23278: dataIn1 = 32'd587
; 
32'd23279: dataIn1 = 32'd590
; 
32'd23280: dataIn1 = 32'd596
; 
32'd23281: dataIn1 = 32'd598
; 
32'd23282: dataIn1 = 32'd619
; 
32'd23283: dataIn1 = 32'd621
; 
32'd23284: dataIn1 = 32'd670
; 
32'd23285: dataIn1 = 32'd690
; 
32'd23286: dataIn1 = 32'd734
; 
32'd23287: dataIn1 = 32'd738
; 
32'd23288: dataIn1 = 32'd747
; 
32'd23289: dataIn1 = 32'd759
; 
32'd23290: dataIn1 = 32'd764
; 
32'd23291: dataIn1 = 32'd786
; 
32'd23292: dataIn1 = 32'd561
; 
32'd23293: dataIn1 = 32'd591
; 
32'd23294: dataIn1 = 32'd625
; 
32'd23295: dataIn1 = 32'd627
; 
32'd23296: dataIn1 = 32'd628
; 
32'd23297: dataIn1 = 32'd634
; 
32'd23298: dataIn1 = 32'd679
; 
32'd23299: dataIn1 = 32'd681
; 
32'd23300: dataIn1 = 32'd689
; 
32'd23301: dataIn1 = 32'd703
; 
32'd23302: dataIn1 = 32'd771
; 
32'd23303: dataIn1 = 32'd778
; 
32'd23304: dataIn1 = 32'd443
; 
32'd23305: dataIn1 = 32'd448
; 
32'd23306: dataIn1 = 32'd455
; 
32'd23307: dataIn1 = 32'd456
; 
32'd23308: dataIn1 = 32'd464
; 
32'd23309: dataIn1 = 32'd565
; 
32'd23310: dataIn1 = 32'd573
; 
32'd23311: dataIn1 = 32'd580
; 
32'd23312: dataIn1 = 32'd617
; 
32'd23313: dataIn1 = 32'd618
; 
32'd23314: dataIn1 = 32'd638
; 
32'd23315: dataIn1 = 32'd640
; 
32'd23316: dataIn1 = 32'd676
; 
32'd23317: dataIn1 = 32'd692
; 
32'd23318: dataIn1 = 32'd693
; 
32'd23319: dataIn1 = 32'd769
; 
32'd23320: dataIn1 = 32'd452
; 
32'd23321: dataIn1 = 32'd467
; 
32'd23322: dataIn1 = 32'd491
; 
32'd23323: dataIn1 = 32'd496
; 
32'd23324: dataIn1 = 32'd505
; 
32'd23325: dataIn1 = 32'd534
; 
32'd23326: dataIn1 = 32'd544
; 
32'd23327: dataIn1 = 32'd545
; 
32'd23328: dataIn1 = 32'd563
; 
32'd23329: dataIn1 = 32'd565
; 
32'd23330: dataIn1 = 32'd606
; 
32'd23331: dataIn1 = 32'd616
; 
32'd23332: dataIn1 = 32'd642
; 
32'd23333: dataIn1 = 32'd650
; 
32'd23334: dataIn1 = 32'd657
; 
32'd23335: dataIn1 = 32'd659
; 
32'd23336: dataIn1 = 32'd671
; 
32'd23337: dataIn1 = 32'd675
; 
32'd23338: dataIn1 = 32'd682
; 
32'd23339: dataIn1 = 32'd689
; 
32'd23340: dataIn1 = 32'd700
; 
32'd23341: dataIn1 = 32'd732
; 
32'd23342: dataIn1 = 32'd746
; 
32'd23343: dataIn1 = 32'd748
; 
32'd23344: dataIn1 = 32'd770
; 
32'd23345: dataIn1 = 32'd787
; 
32'd23346: dataIn1 = 32'd799
; 
32'd23347: dataIn1 = 32'd443
; 
32'd23348: dataIn1 = 32'd449
; 
32'd23349: dataIn1 = 32'd459
; 
32'd23350: dataIn1 = 32'd473
; 
32'd23351: dataIn1 = 32'd496
; 
32'd23352: dataIn1 = 32'd511
; 
32'd23353: dataIn1 = 32'd525
; 
32'd23354: dataIn1 = 32'd598
; 
32'd23355: dataIn1 = 32'd647
; 
32'd23356: dataIn1 = 32'd660
; 
32'd23357: dataIn1 = 32'd690
; 
32'd23358: dataIn1 = 32'd696
; 
32'd23359: dataIn1 = 32'd705
; 
32'd23360: dataIn1 = 32'd706
; 
32'd23361: dataIn1 = 32'd750
; 
32'd23362: dataIn1 = 32'd781
; 
32'd23363: dataIn1 = 32'd785
; 
32'd23364: dataIn1 = 32'd445
; 
32'd23365: dataIn1 = 32'd460
; 
32'd23366: dataIn1 = 32'd495
; 
32'd23367: dataIn1 = 32'd499
; 
32'd23368: dataIn1 = 32'd519
; 
32'd23369: dataIn1 = 32'd528
; 
32'd23370: dataIn1 = 32'd539
; 
32'd23371: dataIn1 = 32'd547
; 
32'd23372: dataIn1 = 32'd562
; 
32'd23373: dataIn1 = 32'd576
; 
32'd23374: dataIn1 = 32'd586
; 
32'd23375: dataIn1 = 32'd590
; 
32'd23376: dataIn1 = 32'd601
; 
32'd23377: dataIn1 = 32'd658
; 
32'd23378: dataIn1 = 32'd660
; 
32'd23379: dataIn1 = 32'd661
; 
32'd23380: dataIn1 = 32'd692
; 
32'd23381: dataIn1 = 32'd697
; 
32'd23382: dataIn1 = 32'd713
; 
32'd23383: dataIn1 = 32'd718
; 
32'd23384: dataIn1 = 32'd724
; 
32'd23385: dataIn1 = 32'd741
; 
32'd23386: dataIn1 = 32'd744
; 
32'd23387: dataIn1 = 32'd746
; 
32'd23388: dataIn1 = 32'd756
; 
32'd23389: dataIn1 = 32'd772
; 
32'd23390: dataIn1 = 32'd778
; 
32'd23391: dataIn1 = 32'd783
; 
32'd23392: dataIn1 = 32'd446
; 
32'd23393: dataIn1 = 32'd472
; 
32'd23394: dataIn1 = 32'd484
; 
32'd23395: dataIn1 = 32'd512
; 
32'd23396: dataIn1 = 32'd520
; 
32'd23397: dataIn1 = 32'd540
; 
32'd23398: dataIn1 = 32'd578
; 
32'd23399: dataIn1 = 32'd641
; 
32'd23400: dataIn1 = 32'd644
; 
32'd23401: dataIn1 = 32'd685
; 
32'd23402: dataIn1 = 32'd718
; 
32'd23403: dataIn1 = 32'd720
; 
32'd23404: dataIn1 = 32'd738
; 
32'd23405: dataIn1 = 32'd740
; 
32'd23406: dataIn1 = 32'd458
; 
32'd23407: dataIn1 = 32'd490
; 
32'd23408: dataIn1 = 32'd493
; 
32'd23409: dataIn1 = 32'd504
; 
32'd23410: dataIn1 = 32'd521
; 
32'd23411: dataIn1 = 32'd527
; 
32'd23412: dataIn1 = 32'd552
; 
32'd23413: dataIn1 = 32'd577
; 
32'd23414: dataIn1 = 32'd583
; 
32'd23415: dataIn1 = 32'd605
; 
32'd23416: dataIn1 = 32'd607
; 
32'd23417: dataIn1 = 32'd618
; 
32'd23418: dataIn1 = 32'd624
; 
32'd23419: dataIn1 = 32'd630
; 
32'd23420: dataIn1 = 32'd647
; 
32'd23421: dataIn1 = 32'd650
; 
32'd23422: dataIn1 = 32'd683
; 
32'd23423: dataIn1 = 32'd694
; 
32'd23424: dataIn1 = 32'd716
; 
32'd23425: dataIn1 = 32'd718
; 
32'd23426: dataIn1 = 32'd727
; 
32'd23427: dataIn1 = 32'd734
; 
32'd23428: dataIn1 = 32'd743
; 
32'd23429: dataIn1 = 32'd746
; 
32'd23430: dataIn1 = 32'd751
; 
32'd23431: dataIn1 = 32'd769
; 
32'd23432: dataIn1 = 32'd772
; 
32'd23433: dataIn1 = 32'd788
; 
32'd23434: dataIn1 = 32'd448
; 
32'd23435: dataIn1 = 32'd454
; 
32'd23436: dataIn1 = 32'd458
; 
32'd23437: dataIn1 = 32'd483
; 
32'd23438: dataIn1 = 32'd487
; 
32'd23439: dataIn1 = 32'd521
; 
32'd23440: dataIn1 = 32'd526
; 
32'd23441: dataIn1 = 32'd531
; 
32'd23442: dataIn1 = 32'd540
; 
32'd23443: dataIn1 = 32'd561
; 
32'd23444: dataIn1 = 32'd562
; 
32'd23445: dataIn1 = 32'd581
; 
32'd23446: dataIn1 = 32'd588
; 
32'd23447: dataIn1 = 32'd592
; 
32'd23448: dataIn1 = 32'd599
; 
32'd23449: dataIn1 = 32'd609
; 
32'd23450: dataIn1 = 32'd612
; 
32'd23451: dataIn1 = 32'd613
; 
32'd23452: dataIn1 = 32'd620
; 
32'd23453: dataIn1 = 32'd623
; 
32'd23454: dataIn1 = 32'd641
; 
32'd23455: dataIn1 = 32'd675
; 
32'd23456: dataIn1 = 32'd676
; 
32'd23457: dataIn1 = 32'd694
; 
32'd23458: dataIn1 = 32'd707
; 
32'd23459: dataIn1 = 32'd710
; 
32'd23460: dataIn1 = 32'd717
; 
32'd23461: dataIn1 = 32'd719
; 
32'd23462: dataIn1 = 32'd737
; 
32'd23463: dataIn1 = 32'd739
; 
32'd23464: dataIn1 = 32'd757
; 
32'd23465: dataIn1 = 32'd775
; 
32'd23466: dataIn1 = 32'd777
; 
32'd23467: dataIn1 = 32'd785
; 
32'd23468: dataIn1 = 32'd799
; 
32'd23469: dataIn1 = 32'd487
; 
32'd23470: dataIn1 = 32'd536
; 
32'd23471: dataIn1 = 32'd549
; 
32'd23472: dataIn1 = 32'd623
; 
32'd23473: dataIn1 = 32'd630
; 
32'd23474: dataIn1 = 32'd650
; 
32'd23475: dataIn1 = 32'd664
; 
32'd23476: dataIn1 = 32'd668
; 
32'd23477: dataIn1 = 32'd700
; 
32'd23478: dataIn1 = 32'd723
; 
32'd23479: dataIn1 = 32'd737
; 
32'd23480: dataIn1 = 32'd747
; 
32'd23481: dataIn1 = 32'd748
; 
32'd23482: dataIn1 = 32'd752
; 
32'd23483: dataIn1 = 32'd759
; 
32'd23484: dataIn1 = 32'd781
; 
32'd23485: dataIn1 = 32'd789
; 
32'd23486: dataIn1 = 32'd474
; 
32'd23487: dataIn1 = 32'd475
; 
32'd23488: dataIn1 = 32'd504
; 
32'd23489: dataIn1 = 32'd506
; 
32'd23490: dataIn1 = 32'd514
; 
32'd23491: dataIn1 = 32'd517
; 
32'd23492: dataIn1 = 32'd518
; 
32'd23493: dataIn1 = 32'd520
; 
32'd23494: dataIn1 = 32'd540
; 
32'd23495: dataIn1 = 32'd552
; 
32'd23496: dataIn1 = 32'd561
; 
32'd23497: dataIn1 = 32'd563
; 
32'd23498: dataIn1 = 32'd577
; 
32'd23499: dataIn1 = 32'd613
; 
32'd23500: dataIn1 = 32'd614
; 
32'd23501: dataIn1 = 32'd621
; 
32'd23502: dataIn1 = 32'd623
; 
32'd23503: dataIn1 = 32'd639
; 
32'd23504: dataIn1 = 32'd667
; 
32'd23505: dataIn1 = 32'd689
; 
32'd23506: dataIn1 = 32'd702
; 
32'd23507: dataIn1 = 32'd708
; 
32'd23508: dataIn1 = 32'd770
; 
32'd23509: dataIn1 = 32'd776
; 
32'd23510: dataIn1 = 32'd783
; 
32'd23511: dataIn1 = 32'd792
; 
32'd23512: dataIn1 = 32'd797
; 
32'd23513: dataIn1 = 32'd469
; 
32'd23514: dataIn1 = 32'd476
; 
32'd23515: dataIn1 = 32'd486
; 
32'd23516: dataIn1 = 32'd492
; 
32'd23517: dataIn1 = 32'd509
; 
32'd23518: dataIn1 = 32'd510
; 
32'd23519: dataIn1 = 32'd521
; 
32'd23520: dataIn1 = 32'd545
; 
32'd23521: dataIn1 = 32'd560
; 
32'd23522: dataIn1 = 32'd584
; 
32'd23523: dataIn1 = 32'd595
; 
32'd23524: dataIn1 = 32'd603
; 
32'd23525: dataIn1 = 32'd618
; 
32'd23526: dataIn1 = 32'd629
; 
32'd23527: dataIn1 = 32'd651
; 
32'd23528: dataIn1 = 32'd652
; 
32'd23529: dataIn1 = 32'd656
; 
32'd23530: dataIn1 = 32'd657
; 
32'd23531: dataIn1 = 32'd662
; 
32'd23532: dataIn1 = 32'd664
; 
32'd23533: dataIn1 = 32'd767
; 
32'd23534: dataIn1 = 32'd786
; 
32'd23535: dataIn1 = 32'd469
; 
32'd23536: dataIn1 = 32'd494
; 
32'd23537: dataIn1 = 32'd543
; 
32'd23538: dataIn1 = 32'd561
; 
32'd23539: dataIn1 = 32'd575
; 
32'd23540: dataIn1 = 32'd595
; 
32'd23541: dataIn1 = 32'd605
; 
32'd23542: dataIn1 = 32'd612
; 
32'd23543: dataIn1 = 32'd618
; 
32'd23544: dataIn1 = 32'd619
; 
32'd23545: dataIn1 = 32'd627
; 
32'd23546: dataIn1 = 32'd657
; 
32'd23547: dataIn1 = 32'd662
; 
32'd23548: dataIn1 = 32'd664
; 
32'd23549: dataIn1 = 32'd679
; 
32'd23550: dataIn1 = 32'd682
; 
32'd23551: dataIn1 = 32'd709
; 
32'd23552: dataIn1 = 32'd715
; 
32'd23553: dataIn1 = 32'd719
; 
32'd23554: dataIn1 = 32'd721
; 
32'd23555: dataIn1 = 32'd736
; 
32'd23556: dataIn1 = 32'd740
; 
32'd23557: dataIn1 = 32'd748
; 
32'd23558: dataIn1 = 32'd784
; 
32'd23559: dataIn1 = 32'd798
; 
32'd23560: dataIn1 = 32'd479
; 
32'd23561: dataIn1 = 32'd508
; 
32'd23562: dataIn1 = 32'd520
; 
32'd23563: dataIn1 = 32'd524
; 
32'd23564: dataIn1 = 32'd525
; 
32'd23565: dataIn1 = 32'd529
; 
32'd23566: dataIn1 = 32'd532
; 
32'd23567: dataIn1 = 32'd549
; 
32'd23568: dataIn1 = 32'd572
; 
32'd23569: dataIn1 = 32'd573
; 
32'd23570: dataIn1 = 32'd595
; 
32'd23571: dataIn1 = 32'd596
; 
32'd23572: dataIn1 = 32'd597
; 
32'd23573: dataIn1 = 32'd646
; 
32'd23574: dataIn1 = 32'd668
; 
32'd23575: dataIn1 = 32'd676
; 
32'd23576: dataIn1 = 32'd678
; 
32'd23577: dataIn1 = 32'd681
; 
32'd23578: dataIn1 = 32'd709
; 
32'd23579: dataIn1 = 32'd757
; 
32'd23580: dataIn1 = 32'd776
; 
32'd23581: dataIn1 = 32'd793
; 
32'd23582: dataIn1 = 32'd465
; 
32'd23583: dataIn1 = 32'd481
; 
32'd23584: dataIn1 = 32'd491
; 
32'd23585: dataIn1 = 32'd499
; 
32'd23586: dataIn1 = 32'd512
; 
32'd23587: dataIn1 = 32'd515
; 
32'd23588: dataIn1 = 32'd544
; 
32'd23589: dataIn1 = 32'd594
; 
32'd23590: dataIn1 = 32'd596
; 
32'd23591: dataIn1 = 32'd610
; 
32'd23592: dataIn1 = 32'd636
; 
32'd23593: dataIn1 = 32'd648
; 
32'd23594: dataIn1 = 32'd650
; 
32'd23595: dataIn1 = 32'd651
; 
32'd23596: dataIn1 = 32'd678
; 
32'd23597: dataIn1 = 32'd681
; 
32'd23598: dataIn1 = 32'd690
; 
32'd23599: dataIn1 = 32'd694
; 
32'd23600: dataIn1 = 32'd752
; 
32'd23601: dataIn1 = 32'd796
; 
32'd23602: dataIn1 = 32'd453
; 
32'd23603: dataIn1 = 32'd463
; 
32'd23604: dataIn1 = 32'd507
; 
32'd23605: dataIn1 = 32'd519
; 
32'd23606: dataIn1 = 32'd559
; 
32'd23607: dataIn1 = 32'd562
; 
32'd23608: dataIn1 = 32'd584
; 
32'd23609: dataIn1 = 32'd591
; 
32'd23610: dataIn1 = 32'd624
; 
32'd23611: dataIn1 = 32'd637
; 
32'd23612: dataIn1 = 32'd651
; 
32'd23613: dataIn1 = 32'd652
; 
32'd23614: dataIn1 = 32'd671
; 
32'd23615: dataIn1 = 32'd724
; 
32'd23616: dataIn1 = 32'd744
; 
32'd23617: dataIn1 = 32'd770
; 
32'd23618: dataIn1 = 32'd798
; 
32'd23619: dataIn1 = 32'd800
; 
32'd23620: dataIn1 = 32'd494
; 
32'd23621: dataIn1 = 32'd498
; 
32'd23622: dataIn1 = 32'd508
; 
32'd23623: dataIn1 = 32'd509
; 
32'd23624: dataIn1 = 32'd512
; 
32'd23625: dataIn1 = 32'd554
; 
32'd23626: dataIn1 = 32'd557
; 
32'd23627: dataIn1 = 32'd578
; 
32'd23628: dataIn1 = 32'd623
; 
32'd23629: dataIn1 = 32'd624
; 
32'd23630: dataIn1 = 32'd629
; 
32'd23631: dataIn1 = 32'd633
; 
32'd23632: dataIn1 = 32'd637
; 
32'd23633: dataIn1 = 32'd650
; 
32'd23634: dataIn1 = 32'd664
; 
32'd23635: dataIn1 = 32'd693
; 
32'd23636: dataIn1 = 32'd694
; 
32'd23637: dataIn1 = 32'd697
; 
32'd23638: dataIn1 = 32'd701
; 
32'd23639: dataIn1 = 32'd709
; 
32'd23640: dataIn1 = 32'd727
; 
32'd23641: dataIn1 = 32'd728
; 
32'd23642: dataIn1 = 32'd741
; 
32'd23643: dataIn1 = 32'd758
; 
32'd23644: dataIn1 = 32'd760
; 
32'd23645: dataIn1 = 32'd779
; 
32'd23646: dataIn1 = 32'd784
; 
32'd23647: dataIn1 = 32'd789
; 
32'd23648: dataIn1 = 32'd473
; 
32'd23649: dataIn1 = 32'd479
; 
32'd23650: dataIn1 = 32'd491
; 
32'd23651: dataIn1 = 32'd567
; 
32'd23652: dataIn1 = 32'd573
; 
32'd23653: dataIn1 = 32'd600
; 
32'd23654: dataIn1 = 32'd629
; 
32'd23655: dataIn1 = 32'd645
; 
32'd23656: dataIn1 = 32'd684
; 
32'd23657: dataIn1 = 32'd712
; 
32'd23658: dataIn1 = 32'd752
; 
32'd23659: dataIn1 = 32'd772
; 
32'd23660: dataIn1 = 32'd793
; 
32'd23661: dataIn1 = 32'd459
; 
32'd23662: dataIn1 = 32'd500
; 
32'd23663: dataIn1 = 32'd520
; 
32'd23664: dataIn1 = 32'd540
; 
32'd23665: dataIn1 = 32'd550
; 
32'd23666: dataIn1 = 32'd587
; 
32'd23667: dataIn1 = 32'd613
; 
32'd23668: dataIn1 = 32'd621
; 
32'd23669: dataIn1 = 32'd643
; 
32'd23670: dataIn1 = 32'd658
; 
32'd23671: dataIn1 = 32'd669
; 
32'd23672: dataIn1 = 32'd673
; 
32'd23673: dataIn1 = 32'd686
; 
32'd23674: dataIn1 = 32'd694
; 
32'd23675: dataIn1 = 32'd725
; 
32'd23676: dataIn1 = 32'd774
; 
32'd23677: dataIn1 = 32'd781
; 
32'd23678: dataIn1 = 32'd787
; 
32'd23679: dataIn1 = 32'd797
; 
32'd23680: dataIn1 = 32'd495
; 
32'd23681: dataIn1 = 32'd502
; 
32'd23682: dataIn1 = 32'd523
; 
32'd23683: dataIn1 = 32'd547
; 
32'd23684: dataIn1 = 32'd553
; 
32'd23685: dataIn1 = 32'd571
; 
32'd23686: dataIn1 = 32'd575
; 
32'd23687: dataIn1 = 32'd597
; 
32'd23688: dataIn1 = 32'd598
; 
32'd23689: dataIn1 = 32'd600
; 
32'd23690: dataIn1 = 32'd607
; 
32'd23691: dataIn1 = 32'd614
; 
32'd23692: dataIn1 = 32'd653
; 
32'd23693: dataIn1 = 32'd669
; 
32'd23694: dataIn1 = 32'd682
; 
32'd23695: dataIn1 = 32'd688
; 
32'd23696: dataIn1 = 32'd689
; 
32'd23697: dataIn1 = 32'd692
; 
32'd23698: dataIn1 = 32'd723
; 
32'd23699: dataIn1 = 32'd754
; 
32'd23700: dataIn1 = 32'd761
; 
32'd23701: dataIn1 = 32'd768
; 
32'd23702: dataIn1 = 32'd772
; 
32'd23703: dataIn1 = 32'd799
; 
32'd23704: dataIn1 = 32'd460
; 
32'd23705: dataIn1 = 32'd464
; 
32'd23706: dataIn1 = 32'd469
; 
32'd23707: dataIn1 = 32'd496
; 
32'd23708: dataIn1 = 32'd504
; 
32'd23709: dataIn1 = 32'd509
; 
32'd23710: dataIn1 = 32'd548
; 
32'd23711: dataIn1 = 32'd568
; 
32'd23712: dataIn1 = 32'd587
; 
32'd23713: dataIn1 = 32'd591
; 
32'd23714: dataIn1 = 32'd594
; 
32'd23715: dataIn1 = 32'd611
; 
32'd23716: dataIn1 = 32'd621
; 
32'd23717: dataIn1 = 32'd656
; 
32'd23718: dataIn1 = 32'd664
; 
32'd23719: dataIn1 = 32'd719
; 
32'd23720: dataIn1 = 32'd765
; 
32'd23721: dataIn1 = 32'd770
; 
32'd23722: dataIn1 = 32'd460
; 
32'd23723: dataIn1 = 32'd506
; 
32'd23724: dataIn1 = 32'd529
; 
32'd23725: dataIn1 = 32'd533
; 
32'd23726: dataIn1 = 32'd548
; 
32'd23727: dataIn1 = 32'd553
; 
32'd23728: dataIn1 = 32'd629
; 
32'd23729: dataIn1 = 32'd662
; 
32'd23730: dataIn1 = 32'd674
; 
32'd23731: dataIn1 = 32'd675
; 
32'd23732: dataIn1 = 32'd689
; 
32'd23733: dataIn1 = 32'd713
; 
32'd23734: dataIn1 = 32'd461
; 
32'd23735: dataIn1 = 32'd482
; 
32'd23736: dataIn1 = 32'd512
; 
32'd23737: dataIn1 = 32'd519
; 
32'd23738: dataIn1 = 32'd554
; 
32'd23739: dataIn1 = 32'd569
; 
32'd23740: dataIn1 = 32'd589
; 
32'd23741: dataIn1 = 32'd600
; 
32'd23742: dataIn1 = 32'd717
; 
32'd23743: dataIn1 = 32'd732
; 
32'd23744: dataIn1 = 32'd782
; 
32'd23745: dataIn1 = 32'd462
; 
32'd23746: dataIn1 = 32'd467
; 
32'd23747: dataIn1 = 32'd483
; 
32'd23748: dataIn1 = 32'd490
; 
32'd23749: dataIn1 = 32'd491
; 
32'd23750: dataIn1 = 32'd544
; 
32'd23751: dataIn1 = 32'd551
; 
32'd23752: dataIn1 = 32'd553
; 
32'd23753: dataIn1 = 32'd611
; 
32'd23754: dataIn1 = 32'd639
; 
32'd23755: dataIn1 = 32'd647
; 
32'd23756: dataIn1 = 32'd671
; 
32'd23757: dataIn1 = 32'd681
; 
32'd23758: dataIn1 = 32'd691
; 
32'd23759: dataIn1 = 32'd755
; 
32'd23760: dataIn1 = 32'd758
; 
32'd23761: dataIn1 = 32'd768
; 
32'd23762: dataIn1 = 32'd773
; 
32'd23763: dataIn1 = 32'd784
; 
32'd23764: dataIn1 = 32'd790
; 
32'd23765: dataIn1 = 32'd482
; 
32'd23766: dataIn1 = 32'd483
; 
32'd23767: dataIn1 = 32'd500
; 
32'd23768: dataIn1 = 32'd502
; 
32'd23769: dataIn1 = 32'd507
; 
32'd23770: dataIn1 = 32'd534
; 
32'd23771: dataIn1 = 32'd553
; 
32'd23772: dataIn1 = 32'd589
; 
32'd23773: dataIn1 = 32'd598
; 
32'd23774: dataIn1 = 32'd628
; 
32'd23775: dataIn1 = 32'd632
; 
32'd23776: dataIn1 = 32'd656
; 
32'd23777: dataIn1 = 32'd720
; 
32'd23778: dataIn1 = 32'd741
; 
32'd23779: dataIn1 = 32'd746
; 
32'd23780: dataIn1 = 32'd750
; 
32'd23781: dataIn1 = 32'd770
; 
32'd23782: dataIn1 = 32'd486
; 
32'd23783: dataIn1 = 32'd489
; 
32'd23784: dataIn1 = 32'd513
; 
32'd23785: dataIn1 = 32'd531
; 
32'd23786: dataIn1 = 32'd537
; 
32'd23787: dataIn1 = 32'd545
; 
32'd23788: dataIn1 = 32'd548
; 
32'd23789: dataIn1 = 32'd557
; 
32'd23790: dataIn1 = 32'd569
; 
32'd23791: dataIn1 = 32'd586
; 
32'd23792: dataIn1 = 32'd588
; 
32'd23793: dataIn1 = 32'd596
; 
32'd23794: dataIn1 = 32'd604
; 
32'd23795: dataIn1 = 32'd613
; 
32'd23796: dataIn1 = 32'd655
; 
32'd23797: dataIn1 = 32'd668
; 
32'd23798: dataIn1 = 32'd669
; 
32'd23799: dataIn1 = 32'd687
; 
32'd23800: dataIn1 = 32'd689
; 
32'd23801: dataIn1 = 32'd696
; 
32'd23802: dataIn1 = 32'd705
; 
32'd23803: dataIn1 = 32'd709
; 
32'd23804: dataIn1 = 32'd762
; 
32'd23805: dataIn1 = 32'd764
; 
32'd23806: dataIn1 = 32'd469
; 
32'd23807: dataIn1 = 32'd588
; 
32'd23808: dataIn1 = 32'd686
; 
32'd23809: dataIn1 = 32'd691
; 
32'd23810: dataIn1 = 32'd746
; 
32'd23811: dataIn1 = 32'd772
; 
32'd23812: dataIn1 = 32'd778
; 
32'd23813: dataIn1 = 32'd795
; 
32'd23814: dataIn1 = 32'd475
; 
32'd23815: dataIn1 = 32'd484
; 
32'd23816: dataIn1 = 32'd486
; 
32'd23817: dataIn1 = 32'd505
; 
32'd23818: dataIn1 = 32'd506
; 
32'd23819: dataIn1 = 32'd517
; 
32'd23820: dataIn1 = 32'd540
; 
32'd23821: dataIn1 = 32'd560
; 
32'd23822: dataIn1 = 32'd571
; 
32'd23823: dataIn1 = 32'd585
; 
32'd23824: dataIn1 = 32'd595
; 
32'd23825: dataIn1 = 32'd719
; 
32'd23826: dataIn1 = 32'd727
; 
32'd23827: dataIn1 = 32'd735
; 
32'd23828: dataIn1 = 32'd743
; 
32'd23829: dataIn1 = 32'd783
; 
32'd23830: dataIn1 = 32'd787
; 
32'd23831: dataIn1 = 32'd796
; 
32'd23832: dataIn1 = 32'd469
; 
32'd23833: dataIn1 = 32'd485
; 
32'd23834: dataIn1 = 32'd487
; 
32'd23835: dataIn1 = 32'd490
; 
32'd23836: dataIn1 = 32'd494
; 
32'd23837: dataIn1 = 32'd503
; 
32'd23838: dataIn1 = 32'd506
; 
32'd23839: dataIn1 = 32'd551
; 
32'd23840: dataIn1 = 32'd556
; 
32'd23841: dataIn1 = 32'd560
; 
32'd23842: dataIn1 = 32'd565
; 
32'd23843: dataIn1 = 32'd569
; 
32'd23844: dataIn1 = 32'd573
; 
32'd23845: dataIn1 = 32'd577
; 
32'd23846: dataIn1 = 32'd601
; 
32'd23847: dataIn1 = 32'd610
; 
32'd23848: dataIn1 = 32'd626
; 
32'd23849: dataIn1 = 32'd636
; 
32'd23850: dataIn1 = 32'd662
; 
32'd23851: dataIn1 = 32'd679
; 
32'd23852: dataIn1 = 32'd690
; 
32'd23853: dataIn1 = 32'd697
; 
32'd23854: dataIn1 = 32'd725
; 
32'd23855: dataIn1 = 32'd783
; 
32'd23856: dataIn1 = 32'd788
; 
32'd23857: dataIn1 = 32'd507
; 
32'd23858: dataIn1 = 32'd515
; 
32'd23859: dataIn1 = 32'd539
; 
32'd23860: dataIn1 = 32'd552
; 
32'd23861: dataIn1 = 32'd561
; 
32'd23862: dataIn1 = 32'd573
; 
32'd23863: dataIn1 = 32'd589
; 
32'd23864: dataIn1 = 32'd596
; 
32'd23865: dataIn1 = 32'd601
; 
32'd23866: dataIn1 = 32'd646
; 
32'd23867: dataIn1 = 32'd650
; 
32'd23868: dataIn1 = 32'd652
; 
32'd23869: dataIn1 = 32'd678
; 
32'd23870: dataIn1 = 32'd680
; 
32'd23871: dataIn1 = 32'd715
; 
32'd23872: dataIn1 = 32'd718
; 
32'd23873: dataIn1 = 32'd740
; 
32'd23874: dataIn1 = 32'd742
; 
32'd23875: dataIn1 = 32'd756
; 
32'd23876: dataIn1 = 32'd780
; 
32'd23877: dataIn1 = 32'd786
; 
32'd23878: dataIn1 = 32'd487
; 
32'd23879: dataIn1 = 32'd516
; 
32'd23880: dataIn1 = 32'd528
; 
32'd23881: dataIn1 = 32'd542
; 
32'd23882: dataIn1 = 32'd543
; 
32'd23883: dataIn1 = 32'd605
; 
32'd23884: dataIn1 = 32'd611
; 
32'd23885: dataIn1 = 32'd630
; 
32'd23886: dataIn1 = 32'd632
; 
32'd23887: dataIn1 = 32'd707
; 
32'd23888: dataIn1 = 32'd730
; 
32'd23889: dataIn1 = 32'd739
; 
32'd23890: dataIn1 = 32'd746
; 
32'd23891: dataIn1 = 32'd764
; 
32'd23892: dataIn1 = 32'd771
; 
32'd23893: dataIn1 = 32'd772
; 
32'd23894: dataIn1 = 32'd780
; 
32'd23895: dataIn1 = 32'd787
; 
32'd23896: dataIn1 = 32'd789
; 
32'd23897: dataIn1 = 32'd790
; 
32'd23898: dataIn1 = 32'd794
; 
32'd23899: dataIn1 = 32'd492
; 
32'd23900: dataIn1 = 32'd500
; 
32'd23901: dataIn1 = 32'd534
; 
32'd23902: dataIn1 = 32'd565
; 
32'd23903: dataIn1 = 32'd568
; 
32'd23904: dataIn1 = 32'd617
; 
32'd23905: dataIn1 = 32'd618
; 
32'd23906: dataIn1 = 32'd621
; 
32'd23907: dataIn1 = 32'd643
; 
32'd23908: dataIn1 = 32'd670
; 
32'd23909: dataIn1 = 32'd682
; 
32'd23910: dataIn1 = 32'd695
; 
32'd23911: dataIn1 = 32'd724
; 
32'd23912: dataIn1 = 32'd799
; 
32'd23913: dataIn1 = 32'd487
; 
32'd23914: dataIn1 = 32'd491
; 
32'd23915: dataIn1 = 32'd533
; 
32'd23916: dataIn1 = 32'd545
; 
32'd23917: dataIn1 = 32'd563
; 
32'd23918: dataIn1 = 32'd574
; 
32'd23919: dataIn1 = 32'd579
; 
32'd23920: dataIn1 = 32'd600
; 
32'd23921: dataIn1 = 32'd613
; 
32'd23922: dataIn1 = 32'd623
; 
32'd23923: dataIn1 = 32'd624
; 
32'd23924: dataIn1 = 32'd626
; 
32'd23925: dataIn1 = 32'd629
; 
32'd23926: dataIn1 = 32'd631
; 
32'd23927: dataIn1 = 32'd636
; 
32'd23928: dataIn1 = 32'd640
; 
32'd23929: dataIn1 = 32'd644
; 
32'd23930: dataIn1 = 32'd671
; 
32'd23931: dataIn1 = 32'd673
; 
32'd23932: dataIn1 = 32'd678
; 
32'd23933: dataIn1 = 32'd688
; 
32'd23934: dataIn1 = 32'd707
; 
32'd23935: dataIn1 = 32'd749
; 
32'd23936: dataIn1 = 32'd751
; 
32'd23937: dataIn1 = 32'd760
; 
32'd23938: dataIn1 = 32'd763
; 
32'd23939: dataIn1 = 32'd768
; 
32'd23940: dataIn1 = 32'd771
; 
32'd23941: dataIn1 = 32'd796
; 
32'd23942: dataIn1 = 32'd482
; 
32'd23943: dataIn1 = 32'd491
; 
32'd23944: dataIn1 = 32'd493
; 
32'd23945: dataIn1 = 32'd498
; 
32'd23946: dataIn1 = 32'd512
; 
32'd23947: dataIn1 = 32'd520
; 
32'd23948: dataIn1 = 32'd535
; 
32'd23949: dataIn1 = 32'd541
; 
32'd23950: dataIn1 = 32'd543
; 
32'd23951: dataIn1 = 32'd565
; 
32'd23952: dataIn1 = 32'd589
; 
32'd23953: dataIn1 = 32'd599
; 
32'd23954: dataIn1 = 32'd659
; 
32'd23955: dataIn1 = 32'd680
; 
32'd23956: dataIn1 = 32'd688
; 
32'd23957: dataIn1 = 32'd693
; 
32'd23958: dataIn1 = 32'd698
; 
32'd23959: dataIn1 = 32'd731
; 
32'd23960: dataIn1 = 32'd739
; 
32'd23961: dataIn1 = 32'd763
; 
32'd23962: dataIn1 = 32'd788
; 
32'd23963: dataIn1 = 32'd507
; 
32'd23964: dataIn1 = 32'd519
; 
32'd23965: dataIn1 = 32'd526
; 
32'd23966: dataIn1 = 32'd532
; 
32'd23967: dataIn1 = 32'd565
; 
32'd23968: dataIn1 = 32'd650
; 
32'd23969: dataIn1 = 32'd658
; 
32'd23970: dataIn1 = 32'd662
; 
32'd23971: dataIn1 = 32'd671
; 
32'd23972: dataIn1 = 32'd679
; 
32'd23973: dataIn1 = 32'd681
; 
32'd23974: dataIn1 = 32'd721
; 
32'd23975: dataIn1 = 32'd736
; 
32'd23976: dataIn1 = 32'd753
; 
32'd23977: dataIn1 = 32'd756
; 
32'd23978: dataIn1 = 32'd758
; 
32'd23979: dataIn1 = 32'd790
; 
32'd23980: dataIn1 = 32'd791
; 
32'd23981: dataIn1 = 32'd477
; 
32'd23982: dataIn1 = 32'd498
; 
32'd23983: dataIn1 = 32'd504
; 
32'd23984: dataIn1 = 32'd537
; 
32'd23985: dataIn1 = 32'd576
; 
32'd23986: dataIn1 = 32'd580
; 
32'd23987: dataIn1 = 32'd581
; 
32'd23988: dataIn1 = 32'd594
; 
32'd23989: dataIn1 = 32'd602
; 
32'd23990: dataIn1 = 32'd630
; 
32'd23991: dataIn1 = 32'd657
; 
32'd23992: dataIn1 = 32'd674
; 
32'd23993: dataIn1 = 32'd676
; 
32'd23994: dataIn1 = 32'd681
; 
32'd23995: dataIn1 = 32'd695
; 
32'd23996: dataIn1 = 32'd702
; 
32'd23997: dataIn1 = 32'd716
; 
32'd23998: dataIn1 = 32'd720
; 
32'd23999: dataIn1 = 32'd751
; 
32'd24000: dataIn1 = 32'd799
; 
32'd24001: dataIn1 = 32'd479
; 
32'd24002: dataIn1 = 32'd497
; 
32'd24003: dataIn1 = 32'd514
; 
32'd24004: dataIn1 = 32'd536
; 
32'd24005: dataIn1 = 32'd553
; 
32'd24006: dataIn1 = 32'd567
; 
32'd24007: dataIn1 = 32'd568
; 
32'd24008: dataIn1 = 32'd595
; 
32'd24009: dataIn1 = 32'd617
; 
32'd24010: dataIn1 = 32'd669
; 
32'd24011: dataIn1 = 32'd687
; 
32'd24012: dataIn1 = 32'd689
; 
32'd24013: dataIn1 = 32'd701
; 
32'd24014: dataIn1 = 32'd714
; 
32'd24015: dataIn1 = 32'd489
; 
32'd24016: dataIn1 = 32'd499
; 
32'd24017: dataIn1 = 32'd502
; 
32'd24018: dataIn1 = 32'd504
; 
32'd24019: dataIn1 = 32'd528
; 
32'd24020: dataIn1 = 32'd552
; 
32'd24021: dataIn1 = 32'd557
; 
32'd24022: dataIn1 = 32'd578
; 
32'd24023: dataIn1 = 32'd583
; 
32'd24024: dataIn1 = 32'd585
; 
32'd24025: dataIn1 = 32'd624
; 
32'd24026: dataIn1 = 32'd646
; 
32'd24027: dataIn1 = 32'd670
; 
32'd24028: dataIn1 = 32'd701
; 
32'd24029: dataIn1 = 32'd707
; 
32'd24030: dataIn1 = 32'd751
; 
32'd24031: dataIn1 = 32'd755
; 
32'd24032: dataIn1 = 32'd764
; 
32'd24033: dataIn1 = 32'd771
; 
32'd24034: dataIn1 = 32'd793
; 
32'd24035: dataIn1 = 32'd496
; 
32'd24036: dataIn1 = 32'd521
; 
32'd24037: dataIn1 = 32'd527
; 
32'd24038: dataIn1 = 32'd540
; 
32'd24039: dataIn1 = 32'd544
; 
32'd24040: dataIn1 = 32'd602
; 
32'd24041: dataIn1 = 32'd609
; 
32'd24042: dataIn1 = 32'd611
; 
32'd24043: dataIn1 = 32'd621
; 
32'd24044: dataIn1 = 32'd634
; 
32'd24045: dataIn1 = 32'd641
; 
32'd24046: dataIn1 = 32'd654
; 
32'd24047: dataIn1 = 32'd674
; 
32'd24048: dataIn1 = 32'd675
; 
32'd24049: dataIn1 = 32'd699
; 
32'd24050: dataIn1 = 32'd704
; 
32'd24051: dataIn1 = 32'd720
; 
32'd24052: dataIn1 = 32'd732
; 
32'd24053: dataIn1 = 32'd759
; 
32'd24054: dataIn1 = 32'd761
; 
32'd24055: dataIn1 = 32'd765
; 
32'd24056: dataIn1 = 32'd768
; 
32'd24057: dataIn1 = 32'd770
; 
32'd24058: dataIn1 = 32'd522
; 
32'd24059: dataIn1 = 32'd533
; 
32'd24060: dataIn1 = 32'd538
; 
32'd24061: dataIn1 = 32'd569
; 
32'd24062: dataIn1 = 32'd585
; 
32'd24063: dataIn1 = 32'd647
; 
32'd24064: dataIn1 = 32'd685
; 
32'd24065: dataIn1 = 32'd690
; 
32'd24066: dataIn1 = 32'd693
; 
32'd24067: dataIn1 = 32'd694
; 
32'd24068: dataIn1 = 32'd695
; 
32'd24069: dataIn1 = 32'd707
; 
32'd24070: dataIn1 = 32'd731
; 
32'd24071: dataIn1 = 32'd738
; 
32'd24072: dataIn1 = 32'd763
; 
32'd24073: dataIn1 = 32'd784
; 
32'd24074: dataIn1 = 32'd480
; 
32'd24075: dataIn1 = 32'd498
; 
32'd24076: dataIn1 = 32'd512
; 
32'd24077: dataIn1 = 32'd519
; 
32'd24078: dataIn1 = 32'd573
; 
32'd24079: dataIn1 = 32'd574
; 
32'd24080: dataIn1 = 32'd576
; 
32'd24081: dataIn1 = 32'd592
; 
32'd24082: dataIn1 = 32'd612
; 
32'd24083: dataIn1 = 32'd627
; 
32'd24084: dataIn1 = 32'd631
; 
32'd24085: dataIn1 = 32'd635
; 
32'd24086: dataIn1 = 32'd658
; 
32'd24087: dataIn1 = 32'd673
; 
32'd24088: dataIn1 = 32'd687
; 
32'd24089: dataIn1 = 32'd688
; 
32'd24090: dataIn1 = 32'd723
; 
32'd24091: dataIn1 = 32'd724
; 
32'd24092: dataIn1 = 32'd726
; 
32'd24093: dataIn1 = 32'd728
; 
32'd24094: dataIn1 = 32'd736
; 
32'd24095: dataIn1 = 32'd789
; 
32'd24096: dataIn1 = 32'd790
; 
32'd24097: dataIn1 = 32'd794
; 
32'd24098: dataIn1 = 32'd502
; 
32'd24099: dataIn1 = 32'd509
; 
32'd24100: dataIn1 = 32'd513
; 
32'd24101: dataIn1 = 32'd518
; 
32'd24102: dataIn1 = 32'd529
; 
32'd24103: dataIn1 = 32'd547
; 
32'd24104: dataIn1 = 32'd584
; 
32'd24105: dataIn1 = 32'd585
; 
32'd24106: dataIn1 = 32'd592
; 
32'd24107: dataIn1 = 32'd605
; 
32'd24108: dataIn1 = 32'd607
; 
32'd24109: dataIn1 = 32'd608
; 
32'd24110: dataIn1 = 32'd629
; 
32'd24111: dataIn1 = 32'd693
; 
32'd24112: dataIn1 = 32'd754
; 
32'd24113: dataIn1 = 32'd777
; 
32'd24114: dataIn1 = 32'd484
; 
32'd24115: dataIn1 = 32'd486
; 
32'd24116: dataIn1 = 32'd492
; 
32'd24117: dataIn1 = 32'd512
; 
32'd24118: dataIn1 = 32'd568
; 
32'd24119: dataIn1 = 32'd570
; 
32'd24120: dataIn1 = 32'd580
; 
32'd24121: dataIn1 = 32'd584
; 
32'd24122: dataIn1 = 32'd591
; 
32'd24123: dataIn1 = 32'd663
; 
32'd24124: dataIn1 = 32'd675
; 
32'd24125: dataIn1 = 32'd688
; 
32'd24126: dataIn1 = 32'd712
; 
32'd24127: dataIn1 = 32'd739
; 
32'd24128: dataIn1 = 32'd757
; 
32'd24129: dataIn1 = 32'd780
; 
32'd24130: dataIn1 = 32'd785
; 
32'd24131: dataIn1 = 32'd484
; 
32'd24132: dataIn1 = 32'd502
; 
32'd24133: dataIn1 = 32'd519
; 
32'd24134: dataIn1 = 32'd546
; 
32'd24135: dataIn1 = 32'd555
; 
32'd24136: dataIn1 = 32'd559
; 
32'd24137: dataIn1 = 32'd566
; 
32'd24138: dataIn1 = 32'd569
; 
32'd24139: dataIn1 = 32'd574
; 
32'd24140: dataIn1 = 32'd575
; 
32'd24141: dataIn1 = 32'd587
; 
32'd24142: dataIn1 = 32'd606
; 
32'd24143: dataIn1 = 32'd662
; 
32'd24144: dataIn1 = 32'd677
; 
32'd24145: dataIn1 = 32'd688
; 
32'd24146: dataIn1 = 32'd708
; 
32'd24147: dataIn1 = 32'd721
; 
32'd24148: dataIn1 = 32'd726
; 
32'd24149: dataIn1 = 32'd736
; 
32'd24150: dataIn1 = 32'd744
; 
32'd24151: dataIn1 = 32'd749
; 
32'd24152: dataIn1 = 32'd750
; 
32'd24153: dataIn1 = 32'd766
; 
32'd24154: dataIn1 = 32'd767
; 
32'd24155: dataIn1 = 32'd789
; 
32'd24156: dataIn1 = 32'd791
; 
32'd24157: dataIn1 = 32'd794
; 
32'd24158: dataIn1 = 32'd492
; 
32'd24159: dataIn1 = 32'd556
; 
32'd24160: dataIn1 = 32'd577
; 
32'd24161: dataIn1 = 32'd584
; 
32'd24162: dataIn1 = 32'd596
; 
32'd24163: dataIn1 = 32'd597
; 
32'd24164: dataIn1 = 32'd615
; 
32'd24165: dataIn1 = 32'd630
; 
32'd24166: dataIn1 = 32'd680
; 
32'd24167: dataIn1 = 32'd687
; 
32'd24168: dataIn1 = 32'd693
; 
32'd24169: dataIn1 = 32'd717
; 
32'd24170: dataIn1 = 32'd746
; 
32'd24171: dataIn1 = 32'd759
; 
32'd24172: dataIn1 = 32'd768
; 
32'd24173: dataIn1 = 32'd783
; 
32'd24174: dataIn1 = 32'd795
; 
32'd24175: dataIn1 = 32'd488
; 
32'd24176: dataIn1 = 32'd492
; 
32'd24177: dataIn1 = 32'd503
; 
32'd24178: dataIn1 = 32'd519
; 
32'd24179: dataIn1 = 32'd541
; 
32'd24180: dataIn1 = 32'd563
; 
32'd24181: dataIn1 = 32'd566
; 
32'd24182: dataIn1 = 32'd613
; 
32'd24183: dataIn1 = 32'd627
; 
32'd24184: dataIn1 = 32'd652
; 
32'd24185: dataIn1 = 32'd664
; 
32'd24186: dataIn1 = 32'd684
; 
32'd24187: dataIn1 = 32'd719
; 
32'd24188: dataIn1 = 32'd741
; 
32'd24189: dataIn1 = 32'd754
; 
32'd24190: dataIn1 = 32'd774
; 
32'd24191: dataIn1 = 32'd781
; 
32'd24192: dataIn1 = 32'd505
; 
32'd24193: dataIn1 = 32'd517
; 
32'd24194: dataIn1 = 32'd518
; 
32'd24195: dataIn1 = 32'd531
; 
32'd24196: dataIn1 = 32'd552
; 
32'd24197: dataIn1 = 32'd571
; 
32'd24198: dataIn1 = 32'd572
; 
32'd24199: dataIn1 = 32'd592
; 
32'd24200: dataIn1 = 32'd605
; 
32'd24201: dataIn1 = 32'd642
; 
32'd24202: dataIn1 = 32'd647
; 
32'd24203: dataIn1 = 32'd654
; 
32'd24204: dataIn1 = 32'd656
; 
32'd24205: dataIn1 = 32'd701
; 
32'd24206: dataIn1 = 32'd704
; 
32'd24207: dataIn1 = 32'd711
; 
32'd24208: dataIn1 = 32'd735
; 
32'd24209: dataIn1 = 32'd742
; 
32'd24210: dataIn1 = 32'd795
; 
32'd24211: dataIn1 = 32'd515
; 
32'd24212: dataIn1 = 32'd537
; 
32'd24213: dataIn1 = 32'd571
; 
32'd24214: dataIn1 = 32'd575
; 
32'd24215: dataIn1 = 32'd584
; 
32'd24216: dataIn1 = 32'd595
; 
32'd24217: dataIn1 = 32'd603
; 
32'd24218: dataIn1 = 32'd608
; 
32'd24219: dataIn1 = 32'd614
; 
32'd24220: dataIn1 = 32'd620
; 
32'd24221: dataIn1 = 32'd631
; 
32'd24222: dataIn1 = 32'd632
; 
32'd24223: dataIn1 = 32'd634
; 
32'd24224: dataIn1 = 32'd644
; 
32'd24225: dataIn1 = 32'd660
; 
32'd24226: dataIn1 = 32'd688
; 
32'd24227: dataIn1 = 32'd713
; 
32'd24228: dataIn1 = 32'd723
; 
32'd24229: dataIn1 = 32'd758
; 
32'd24230: dataIn1 = 32'd765
; 
32'd24231: dataIn1 = 32'd767
; 
32'd24232: dataIn1 = 32'd503
; 
32'd24233: dataIn1 = 32'd525
; 
32'd24234: dataIn1 = 32'd537
; 
32'd24235: dataIn1 = 32'd553
; 
32'd24236: dataIn1 = 32'd555
; 
32'd24237: dataIn1 = 32'd586
; 
32'd24238: dataIn1 = 32'd600
; 
32'd24239: dataIn1 = 32'd628
; 
32'd24240: dataIn1 = 32'd637
; 
32'd24241: dataIn1 = 32'd648
; 
32'd24242: dataIn1 = 32'd662
; 
32'd24243: dataIn1 = 32'd665
; 
32'd24244: dataIn1 = 32'd678
; 
32'd24245: dataIn1 = 32'd686
; 
32'd24246: dataIn1 = 32'd692
; 
32'd24247: dataIn1 = 32'd730
; 
32'd24248: dataIn1 = 32'd762
; 
32'd24249: dataIn1 = 32'd768
; 
32'd24250: dataIn1 = 32'd775
; 
32'd24251: dataIn1 = 32'd777
; 
32'd24252: dataIn1 = 32'd787
; 
32'd24253: dataIn1 = 32'd789
; 
32'd24254: dataIn1 = 32'd507
; 
32'd24255: dataIn1 = 32'd527
; 
32'd24256: dataIn1 = 32'd529
; 
32'd24257: dataIn1 = 32'd533
; 
32'd24258: dataIn1 = 32'd536
; 
32'd24259: dataIn1 = 32'd538
; 
32'd24260: dataIn1 = 32'd547
; 
32'd24261: dataIn1 = 32'd548
; 
32'd24262: dataIn1 = 32'd558
; 
32'd24263: dataIn1 = 32'd562
; 
32'd24264: dataIn1 = 32'd597
; 
32'd24265: dataIn1 = 32'd601
; 
32'd24266: dataIn1 = 32'd614
; 
32'd24267: dataIn1 = 32'd623
; 
32'd24268: dataIn1 = 32'd649
; 
32'd24269: dataIn1 = 32'd656
; 
32'd24270: dataIn1 = 32'd699
; 
32'd24271: dataIn1 = 32'd705
; 
32'd24272: dataIn1 = 32'd718
; 
32'd24273: dataIn1 = 32'd727
; 
32'd24274: dataIn1 = 32'd732
; 
32'd24275: dataIn1 = 32'd733
; 
32'd24276: dataIn1 = 32'd782
; 
32'd24277: dataIn1 = 32'd524
; 
32'd24278: dataIn1 = 32'd527
; 
32'd24279: dataIn1 = 32'd539
; 
32'd24280: dataIn1 = 32'd553
; 
32'd24281: dataIn1 = 32'd555
; 
32'd24282: dataIn1 = 32'd579
; 
32'd24283: dataIn1 = 32'd580
; 
32'd24284: dataIn1 = 32'd599
; 
32'd24285: dataIn1 = 32'd615
; 
32'd24286: dataIn1 = 32'd620
; 
32'd24287: dataIn1 = 32'd631
; 
32'd24288: dataIn1 = 32'd637
; 
32'd24289: dataIn1 = 32'd659
; 
32'd24290: dataIn1 = 32'd663
; 
32'd24291: dataIn1 = 32'd666
; 
32'd24292: dataIn1 = 32'd680
; 
32'd24293: dataIn1 = 32'd705
; 
32'd24294: dataIn1 = 32'd711
; 
32'd24295: dataIn1 = 32'd725
; 
32'd24296: dataIn1 = 32'd737
; 
32'd24297: dataIn1 = 32'd761
; 
32'd24298: dataIn1 = 32'd771
; 
32'd24299: dataIn1 = 32'd790
; 
32'd24300: dataIn1 = 32'd494
; 
32'd24301: dataIn1 = 32'd502
; 
32'd24302: dataIn1 = 32'd505
; 
32'd24303: dataIn1 = 32'd510
; 
32'd24304: dataIn1 = 32'd521
; 
32'd24305: dataIn1 = 32'd538
; 
32'd24306: dataIn1 = 32'd556
; 
32'd24307: dataIn1 = 32'd570
; 
32'd24308: dataIn1 = 32'd592
; 
32'd24309: dataIn1 = 32'd614
; 
32'd24310: dataIn1 = 32'd640
; 
32'd24311: dataIn1 = 32'd651
; 
32'd24312: dataIn1 = 32'd655
; 
32'd24313: dataIn1 = 32'd677
; 
32'd24314: dataIn1 = 32'd680
; 
32'd24315: dataIn1 = 32'd683
; 
32'd24316: dataIn1 = 32'd698
; 
32'd24317: dataIn1 = 32'd703
; 
32'd24318: dataIn1 = 32'd724
; 
32'd24319: dataIn1 = 32'd728
; 
32'd24320: dataIn1 = 32'd742
; 
32'd24321: dataIn1 = 32'd753
; 
32'd24322: dataIn1 = 32'd786
; 
32'd24323: dataIn1 = 32'd535
; 
32'd24324: dataIn1 = 32'd551
; 
32'd24325: dataIn1 = 32'd576
; 
32'd24326: dataIn1 = 32'd616
; 
32'd24327: dataIn1 = 32'd623
; 
32'd24328: dataIn1 = 32'd640
; 
32'd24329: dataIn1 = 32'd653
; 
32'd24330: dataIn1 = 32'd683
; 
32'd24331: dataIn1 = 32'd690
; 
32'd24332: dataIn1 = 32'd698
; 
32'd24333: dataIn1 = 32'd721
; 
32'd24334: dataIn1 = 32'd750
; 
32'd24335: dataIn1 = 32'd763
; 
32'd24336: dataIn1 = 32'd500
; 
32'd24337: dataIn1 = 32'd507
; 
32'd24338: dataIn1 = 32'd510
; 
32'd24339: dataIn1 = 32'd553
; 
32'd24340: dataIn1 = 32'd562
; 
32'd24341: dataIn1 = 32'd579
; 
32'd24342: dataIn1 = 32'd588
; 
32'd24343: dataIn1 = 32'd591
; 
32'd24344: dataIn1 = 32'd598
; 
32'd24345: dataIn1 = 32'd629
; 
32'd24346: dataIn1 = 32'd646
; 
32'd24347: dataIn1 = 32'd660
; 
32'd24348: dataIn1 = 32'd661
; 
32'd24349: dataIn1 = 32'd681
; 
32'd24350: dataIn1 = 32'd687
; 
32'd24351: dataIn1 = 32'd702
; 
32'd24352: dataIn1 = 32'd724
; 
32'd24353: dataIn1 = 32'd738
; 
32'd24354: dataIn1 = 32'd753
; 
32'd24355: dataIn1 = 32'd788
; 
32'd24356: dataIn1 = 32'd799
; 
32'd24357: dataIn1 = 32'd500
; 
32'd24358: dataIn1 = 32'd515
; 
32'd24359: dataIn1 = 32'd525
; 
32'd24360: dataIn1 = 32'd531
; 
32'd24361: dataIn1 = 32'd545
; 
32'd24362: dataIn1 = 32'd553
; 
32'd24363: dataIn1 = 32'd558
; 
32'd24364: dataIn1 = 32'd572
; 
32'd24365: dataIn1 = 32'd577
; 
32'd24366: dataIn1 = 32'd585
; 
32'd24367: dataIn1 = 32'd636
; 
32'd24368: dataIn1 = 32'd641
; 
32'd24369: dataIn1 = 32'd647
; 
32'd24370: dataIn1 = 32'd648
; 
32'd24371: dataIn1 = 32'd656
; 
32'd24372: dataIn1 = 32'd659
; 
32'd24373: dataIn1 = 32'd678
; 
32'd24374: dataIn1 = 32'd742
; 
32'd24375: dataIn1 = 32'd779
; 
32'd24376: dataIn1 = 32'd791
; 
32'd24377: dataIn1 = 32'd794
; 
32'd24378: dataIn1 = 32'd796
; 
32'd24379: dataIn1 = 32'd499
; 
32'd24380: dataIn1 = 32'd506
; 
32'd24381: dataIn1 = 32'd521
; 
32'd24382: dataIn1 = 32'd522
; 
32'd24383: dataIn1 = 32'd533
; 
32'd24384: dataIn1 = 32'd544
; 
32'd24385: dataIn1 = 32'd567
; 
32'd24386: dataIn1 = 32'd581
; 
32'd24387: dataIn1 = 32'd582
; 
32'd24388: dataIn1 = 32'd607
; 
32'd24389: dataIn1 = 32'd610
; 
32'd24390: dataIn1 = 32'd637
; 
32'd24391: dataIn1 = 32'd673
; 
32'd24392: dataIn1 = 32'd685
; 
32'd24393: dataIn1 = 32'd696
; 
32'd24394: dataIn1 = 32'd704
; 
32'd24395: dataIn1 = 32'd710
; 
32'd24396: dataIn1 = 32'd726
; 
32'd24397: dataIn1 = 32'd730
; 
32'd24398: dataIn1 = 32'd741
; 
32'd24399: dataIn1 = 32'd764
; 
32'd24400: dataIn1 = 32'd765
; 
32'd24401: dataIn1 = 32'd771
; 
32'd24402: dataIn1 = 32'd786
; 
32'd24403: dataIn1 = 32'd794
; 
32'd24404: dataIn1 = 32'd526
; 
32'd24405: dataIn1 = 32'd541
; 
32'd24406: dataIn1 = 32'd552
; 
32'd24407: dataIn1 = 32'd564
; 
32'd24408: dataIn1 = 32'd567
; 
32'd24409: dataIn1 = 32'd596
; 
32'd24410: dataIn1 = 32'd608
; 
32'd24411: dataIn1 = 32'd625
; 
32'd24412: dataIn1 = 32'd646
; 
32'd24413: dataIn1 = 32'd655
; 
32'd24414: dataIn1 = 32'd668
; 
32'd24415: dataIn1 = 32'd685
; 
32'd24416: dataIn1 = 32'd705
; 
32'd24417: dataIn1 = 32'd708
; 
32'd24418: dataIn1 = 32'd712
; 
32'd24419: dataIn1 = 32'd713
; 
32'd24420: dataIn1 = 32'd720
; 
32'd24421: dataIn1 = 32'd730
; 
32'd24422: dataIn1 = 32'd734
; 
32'd24423: dataIn1 = 32'd736
; 
32'd24424: dataIn1 = 32'd739
; 
32'd24425: dataIn1 = 32'd749
; 
32'd24426: dataIn1 = 32'd758
; 
32'd24427: dataIn1 = 32'd779
; 
32'd24428: dataIn1 = 32'd785
; 
32'd24429: dataIn1 = 32'd510
; 
32'd24430: dataIn1 = 32'd530
; 
32'd24431: dataIn1 = 32'd537
; 
32'd24432: dataIn1 = 32'd596
; 
32'd24433: dataIn1 = 32'd597
; 
32'd24434: dataIn1 = 32'd599
; 
32'd24435: dataIn1 = 32'd617
; 
32'd24436: dataIn1 = 32'd619
; 
32'd24437: dataIn1 = 32'd633
; 
32'd24438: dataIn1 = 32'd635
; 
32'd24439: dataIn1 = 32'd646
; 
32'd24440: dataIn1 = 32'd731
; 
32'd24441: dataIn1 = 32'd737
; 
32'd24442: dataIn1 = 32'd789
; 
32'd24443: dataIn1 = 32'd515
; 
32'd24444: dataIn1 = 32'd554
; 
32'd24445: dataIn1 = 32'd568
; 
32'd24446: dataIn1 = 32'd570
; 
32'd24447: dataIn1 = 32'd601
; 
32'd24448: dataIn1 = 32'd605
; 
32'd24449: dataIn1 = 32'd617
; 
32'd24450: dataIn1 = 32'd618
; 
32'd24451: dataIn1 = 32'd635
; 
32'd24452: dataIn1 = 32'd645
; 
32'd24453: dataIn1 = 32'd677
; 
32'd24454: dataIn1 = 32'd742
; 
32'd24455: dataIn1 = 32'd743
; 
32'd24456: dataIn1 = 32'd745
; 
32'd24457: dataIn1 = 32'd782
; 
32'd24458: dataIn1 = 32'd517
; 
32'd24459: dataIn1 = 32'd553
; 
32'd24460: dataIn1 = 32'd556
; 
32'd24461: dataIn1 = 32'd600
; 
32'd24462: dataIn1 = 32'd613
; 
32'd24463: dataIn1 = 32'd621
; 
32'd24464: dataIn1 = 32'd626
; 
32'd24465: dataIn1 = 32'd627
; 
32'd24466: dataIn1 = 32'd657
; 
32'd24467: dataIn1 = 32'd725
; 
32'd24468: dataIn1 = 32'd775
; 
32'd24469: dataIn1 = 32'd794
; 
32'd24470: dataIn1 = 32'd797
; 
32'd24471: dataIn1 = 32'd511
; 
32'd24472: dataIn1 = 32'd531
; 
32'd24473: dataIn1 = 32'd532
; 
32'd24474: dataIn1 = 32'd536
; 
32'd24475: dataIn1 = 32'd542
; 
32'd24476: dataIn1 = 32'd594
; 
32'd24477: dataIn1 = 32'd624
; 
32'd24478: dataIn1 = 32'd649
; 
32'd24479: dataIn1 = 32'd652
; 
32'd24480: dataIn1 = 32'd671
; 
32'd24481: dataIn1 = 32'd678
; 
32'd24482: dataIn1 = 32'd691
; 
32'd24483: dataIn1 = 32'd721
; 
32'd24484: dataIn1 = 32'd725
; 
32'd24485: dataIn1 = 32'd731
; 
32'd24486: dataIn1 = 32'd767
; 
32'd24487: dataIn1 = 32'd769
; 
32'd24488: dataIn1 = 32'd783
; 
32'd24489: dataIn1 = 32'd511
; 
32'd24490: dataIn1 = 32'd516
; 
32'd24491: dataIn1 = 32'd519
; 
32'd24492: dataIn1 = 32'd552
; 
32'd24493: dataIn1 = 32'd561
; 
32'd24494: dataIn1 = 32'd562
; 
32'd24495: dataIn1 = 32'd582
; 
32'd24496: dataIn1 = 32'd594
; 
32'd24497: dataIn1 = 32'd601
; 
32'd24498: dataIn1 = 32'd610
; 
32'd24499: dataIn1 = 32'd619
; 
32'd24500: dataIn1 = 32'd622
; 
32'd24501: dataIn1 = 32'd642
; 
32'd24502: dataIn1 = 32'd662
; 
32'd24503: dataIn1 = 32'd663
; 
32'd24504: dataIn1 = 32'd669
; 
32'd24505: dataIn1 = 32'd704
; 
32'd24506: dataIn1 = 32'd724
; 
32'd24507: dataIn1 = 32'd735
; 
32'd24508: dataIn1 = 32'd772
; 
32'd24509: dataIn1 = 32'd780
; 
32'd24510: dataIn1 = 32'd514
; 
32'd24511: dataIn1 = 32'd560
; 
32'd24512: dataIn1 = 32'd568
; 
32'd24513: dataIn1 = 32'd584
; 
32'd24514: dataIn1 = 32'd617
; 
32'd24515: dataIn1 = 32'd624
; 
32'd24516: dataIn1 = 32'd660
; 
32'd24517: dataIn1 = 32'd666
; 
32'd24518: dataIn1 = 32'd682
; 
32'd24519: dataIn1 = 32'd684
; 
32'd24520: dataIn1 = 32'd687
; 
32'd24521: dataIn1 = 32'd690
; 
32'd24522: dataIn1 = 32'd708
; 
32'd24523: dataIn1 = 32'd747
; 
32'd24524: dataIn1 = 32'd754
; 
32'd24525: dataIn1 = 32'd758
; 
32'd24526: dataIn1 = 32'd780
; 
32'd24527: dataIn1 = 32'd788
; 
32'd24528: dataIn1 = 32'd560
; 
32'd24529: dataIn1 = 32'd568
; 
32'd24530: dataIn1 = 32'd572
; 
32'd24531: dataIn1 = 32'd574
; 
32'd24532: dataIn1 = 32'd588
; 
32'd24533: dataIn1 = 32'd598
; 
32'd24534: dataIn1 = 32'd622
; 
32'd24535: dataIn1 = 32'd645
; 
32'd24536: dataIn1 = 32'd661
; 
32'd24537: dataIn1 = 32'd684
; 
32'd24538: dataIn1 = 32'd687
; 
32'd24539: dataIn1 = 32'd696
; 
32'd24540: dataIn1 = 32'd702
; 
32'd24541: dataIn1 = 32'd739
; 
32'd24542: dataIn1 = 32'd751
; 
32'd24543: dataIn1 = 32'd761
; 
32'd24544: dataIn1 = 32'd775
; 
32'd24545: dataIn1 = 32'd540
; 
32'd24546: dataIn1 = 32'd549
; 
32'd24547: dataIn1 = 32'd566
; 
32'd24548: dataIn1 = 32'd619
; 
32'd24549: dataIn1 = 32'd656
; 
32'd24550: dataIn1 = 32'd691
; 
32'd24551: dataIn1 = 32'd693
; 
32'd24552: dataIn1 = 32'd719
; 
32'd24553: dataIn1 = 32'd728
; 
32'd24554: dataIn1 = 32'd731
; 
32'd24555: dataIn1 = 32'd769
; 
32'd24556: dataIn1 = 32'd782
; 
32'd24557: dataIn1 = 32'd783
; 
32'd24558: dataIn1 = 32'd790
; 
32'd24559: dataIn1 = 32'd523
; 
32'd24560: dataIn1 = 32'd543
; 
32'd24561: dataIn1 = 32'd580
; 
32'd24562: dataIn1 = 32'd587
; 
32'd24563: dataIn1 = 32'd599
; 
32'd24564: dataIn1 = 32'd612
; 
32'd24565: dataIn1 = 32'd614
; 
32'd24566: dataIn1 = 32'd632
; 
32'd24567: dataIn1 = 32'd665
; 
32'd24568: dataIn1 = 32'd681
; 
32'd24569: dataIn1 = 32'd696
; 
32'd24570: dataIn1 = 32'd706
; 
32'd24571: dataIn1 = 32'd778
; 
32'd24572: dataIn1 = 32'd789
; 
32'd24573: dataIn1 = 32'd510
; 
32'd24574: dataIn1 = 32'd538
; 
32'd24575: dataIn1 = 32'd544
; 
32'd24576: dataIn1 = 32'd563
; 
32'd24577: dataIn1 = 32'd587
; 
32'd24578: dataIn1 = 32'd596
; 
32'd24579: dataIn1 = 32'd601
; 
32'd24580: dataIn1 = 32'd603
; 
32'd24581: dataIn1 = 32'd647
; 
32'd24582: dataIn1 = 32'd657
; 
32'd24583: dataIn1 = 32'd669
; 
32'd24584: dataIn1 = 32'd673
; 
32'd24585: dataIn1 = 32'd701
; 
32'd24586: dataIn1 = 32'd713
; 
32'd24587: dataIn1 = 32'd716
; 
32'd24588: dataIn1 = 32'd720
; 
32'd24589: dataIn1 = 32'd736
; 
32'd24590: dataIn1 = 32'd747
; 
32'd24591: dataIn1 = 32'd757
; 
32'd24592: dataIn1 = 32'd523
; 
32'd24593: dataIn1 = 32'd544
; 
32'd24594: dataIn1 = 32'd569
; 
32'd24595: dataIn1 = 32'd585
; 
32'd24596: dataIn1 = 32'd640
; 
32'd24597: dataIn1 = 32'd704
; 
32'd24598: dataIn1 = 32'd707
; 
32'd24599: dataIn1 = 32'd719
; 
32'd24600: dataIn1 = 32'd726
; 
32'd24601: dataIn1 = 32'd733
; 
32'd24602: dataIn1 = 32'd769
; 
32'd24603: dataIn1 = 32'd788
; 
32'd24604: dataIn1 = 32'd789
; 
32'd24605: dataIn1 = 32'd794
; 
32'd24606: dataIn1 = 32'd513
; 
32'd24607: dataIn1 = 32'd522
; 
32'd24608: dataIn1 = 32'd541
; 
32'd24609: dataIn1 = 32'd557
; 
32'd24610: dataIn1 = 32'd568
; 
32'd24611: dataIn1 = 32'd587
; 
32'd24612: dataIn1 = 32'd596
; 
32'd24613: dataIn1 = 32'd605
; 
32'd24614: dataIn1 = 32'd633
; 
32'd24615: dataIn1 = 32'd646
; 
32'd24616: dataIn1 = 32'd666
; 
32'd24617: dataIn1 = 32'd717
; 
32'd24618: dataIn1 = 32'd732
; 
32'd24619: dataIn1 = 32'd744
; 
32'd24620: dataIn1 = 32'd761
; 
32'd24621: dataIn1 = 32'd785
; 
32'd24622: dataIn1 = 32'd540
; 
32'd24623: dataIn1 = 32'd545
; 
32'd24624: dataIn1 = 32'd554
; 
32'd24625: dataIn1 = 32'd578
; 
32'd24626: dataIn1 = 32'd588
; 
32'd24627: dataIn1 = 32'd589
; 
32'd24628: dataIn1 = 32'd595
; 
32'd24629: dataIn1 = 32'd613
; 
32'd24630: dataIn1 = 32'd627
; 
32'd24631: dataIn1 = 32'd643
; 
32'd24632: dataIn1 = 32'd671
; 
32'd24633: dataIn1 = 32'd679
; 
32'd24634: dataIn1 = 32'd683
; 
32'd24635: dataIn1 = 32'd684
; 
32'd24636: dataIn1 = 32'd688
; 
32'd24637: dataIn1 = 32'd702
; 
32'd24638: dataIn1 = 32'd708
; 
32'd24639: dataIn1 = 32'd720
; 
32'd24640: dataIn1 = 32'd729
; 
32'd24641: dataIn1 = 32'd774
; 
32'd24642: dataIn1 = 32'd781
; 
32'd24643: dataIn1 = 32'd512
; 
32'd24644: dataIn1 = 32'd533
; 
32'd24645: dataIn1 = 32'd549
; 
32'd24646: dataIn1 = 32'd572
; 
32'd24647: dataIn1 = 32'd583
; 
32'd24648: dataIn1 = 32'd593
; 
32'd24649: dataIn1 = 32'd610
; 
32'd24650: dataIn1 = 32'd613
; 
32'd24651: dataIn1 = 32'd629
; 
32'd24652: dataIn1 = 32'd645
; 
32'd24653: dataIn1 = 32'd721
; 
32'd24654: dataIn1 = 32'd724
; 
32'd24655: dataIn1 = 32'd731
; 
32'd24656: dataIn1 = 32'd742
; 
32'd24657: dataIn1 = 32'd746
; 
32'd24658: dataIn1 = 32'd777
; 
32'd24659: dataIn1 = 32'd778
; 
32'd24660: dataIn1 = 32'd523
; 
32'd24661: dataIn1 = 32'd535
; 
32'd24662: dataIn1 = 32'd536
; 
32'd24663: dataIn1 = 32'd544
; 
32'd24664: dataIn1 = 32'd564
; 
32'd24665: dataIn1 = 32'd574
; 
32'd24666: dataIn1 = 32'd591
; 
32'd24667: dataIn1 = 32'd593
; 
32'd24668: dataIn1 = 32'd610
; 
32'd24669: dataIn1 = 32'd617
; 
32'd24670: dataIn1 = 32'd646
; 
32'd24671: dataIn1 = 32'd667
; 
32'd24672: dataIn1 = 32'd680
; 
32'd24673: dataIn1 = 32'd698
; 
32'd24674: dataIn1 = 32'd734
; 
32'd24675: dataIn1 = 32'd755
; 
32'd24676: dataIn1 = 32'd770
; 
32'd24677: dataIn1 = 32'd799
; 
32'd24678: dataIn1 = 32'd536
; 
32'd24679: dataIn1 = 32'd548
; 
32'd24680: dataIn1 = 32'd579
; 
32'd24681: dataIn1 = 32'd616
; 
32'd24682: dataIn1 = 32'd659
; 
32'd24683: dataIn1 = 32'd671
; 
32'd24684: dataIn1 = 32'd722
; 
32'd24685: dataIn1 = 32'd771
; 
32'd24686: dataIn1 = 32'd775
; 
32'd24687: dataIn1 = 32'd787
; 
32'd24688: dataIn1 = 32'd520
; 
32'd24689: dataIn1 = 32'd521
; 
32'd24690: dataIn1 = 32'd545
; 
32'd24691: dataIn1 = 32'd607
; 
32'd24692: dataIn1 = 32'd615
; 
32'd24693: dataIn1 = 32'd665
; 
32'd24694: dataIn1 = 32'd686
; 
32'd24695: dataIn1 = 32'd690
; 
32'd24696: dataIn1 = 32'd691
; 
32'd24697: dataIn1 = 32'd710
; 
32'd24698: dataIn1 = 32'd711
; 
32'd24699: dataIn1 = 32'd713
; 
32'd24700: dataIn1 = 32'd715
; 
32'd24701: dataIn1 = 32'd724
; 
32'd24702: dataIn1 = 32'd737
; 
32'd24703: dataIn1 = 32'd751
; 
32'd24704: dataIn1 = 32'd752
; 
32'd24705: dataIn1 = 32'd766
; 
32'd24706: dataIn1 = 32'd788
; 
32'd24707: dataIn1 = 32'd530
; 
32'd24708: dataIn1 = 32'd546
; 
32'd24709: dataIn1 = 32'd550
; 
32'd24710: dataIn1 = 32'd556
; 
32'd24711: dataIn1 = 32'd577
; 
32'd24712: dataIn1 = 32'd597
; 
32'd24713: dataIn1 = 32'd647
; 
32'd24714: dataIn1 = 32'd654
; 
32'd24715: dataIn1 = 32'd702
; 
32'd24716: dataIn1 = 32'd717
; 
32'd24717: dataIn1 = 32'd732
; 
32'd24718: dataIn1 = 32'd736
; 
32'd24719: dataIn1 = 32'd746
; 
32'd24720: dataIn1 = 32'd758
; 
32'd24721: dataIn1 = 32'd763
; 
32'd24722: dataIn1 = 32'd775
; 
32'd24723: dataIn1 = 32'd795
; 
32'd24724: dataIn1 = 32'd558
; 
32'd24725: dataIn1 = 32'd565
; 
32'd24726: dataIn1 = 32'd605
; 
32'd24727: dataIn1 = 32'd608
; 
32'd24728: dataIn1 = 32'd621
; 
32'd24729: dataIn1 = 32'd657
; 
32'd24730: dataIn1 = 32'd679
; 
32'd24731: dataIn1 = 32'd686
; 
32'd24732: dataIn1 = 32'd719
; 
32'd24733: dataIn1 = 32'd734
; 
32'd24734: dataIn1 = 32'd531
; 
32'd24735: dataIn1 = 32'd541
; 
32'd24736: dataIn1 = 32'd550
; 
32'd24737: dataIn1 = 32'd570
; 
32'd24738: dataIn1 = 32'd576
; 
32'd24739: dataIn1 = 32'd582
; 
32'd24740: dataIn1 = 32'd601
; 
32'd24741: dataIn1 = 32'd606
; 
32'd24742: dataIn1 = 32'd625
; 
32'd24743: dataIn1 = 32'd628
; 
32'd24744: dataIn1 = 32'd637
; 
32'd24745: dataIn1 = 32'd644
; 
32'd24746: dataIn1 = 32'd646
; 
32'd24747: dataIn1 = 32'd674
; 
32'd24748: dataIn1 = 32'd681
; 
32'd24749: dataIn1 = 32'd697
; 
32'd24750: dataIn1 = 32'd703
; 
32'd24751: dataIn1 = 32'd713
; 
32'd24752: dataIn1 = 32'd720
; 
32'd24753: dataIn1 = 32'd745
; 
32'd24754: dataIn1 = 32'd749
; 
32'd24755: dataIn1 = 32'd772
; 
32'd24756: dataIn1 = 32'd776
; 
32'd24757: dataIn1 = 32'd777
; 
32'd24758: dataIn1 = 32'd518
; 
32'd24759: dataIn1 = 32'd551
; 
32'd24760: dataIn1 = 32'd584
; 
32'd24761: dataIn1 = 32'd604
; 
32'd24762: dataIn1 = 32'd615
; 
32'd24763: dataIn1 = 32'd622
; 
32'd24764: dataIn1 = 32'd638
; 
32'd24765: dataIn1 = 32'd655
; 
32'd24766: dataIn1 = 32'd681
; 
32'd24767: dataIn1 = 32'd691
; 
32'd24768: dataIn1 = 32'd694
; 
32'd24769: dataIn1 = 32'd713
; 
32'd24770: dataIn1 = 32'd740
; 
32'd24771: dataIn1 = 32'd760
; 
32'd24772: dataIn1 = 32'd775
; 
32'd24773: dataIn1 = 32'd573
; 
32'd24774: dataIn1 = 32'd595
; 
32'd24775: dataIn1 = 32'd610
; 
32'd24776: dataIn1 = 32'd613
; 
32'd24777: dataIn1 = 32'd621
; 
32'd24778: dataIn1 = 32'd632
; 
32'd24779: dataIn1 = 32'd671
; 
32'd24780: dataIn1 = 32'd681
; 
32'd24781: dataIn1 = 32'd688
; 
32'd24782: dataIn1 = 32'd710
; 
32'd24783: dataIn1 = 32'd714
; 
32'd24784: dataIn1 = 32'd749
; 
32'd24785: dataIn1 = 32'd753
; 
32'd24786: dataIn1 = 32'd755
; 
32'd24787: dataIn1 = 32'd777
; 
32'd24788: dataIn1 = 32'd785
; 
32'd24789: dataIn1 = 32'd796
; 
32'd24790: dataIn1 = 32'd799
; 
32'd24791: dataIn1 = 32'd535
; 
32'd24792: dataIn1 = 32'd571
; 
32'd24793: dataIn1 = 32'd593
; 
32'd24794: dataIn1 = 32'd594
; 
32'd24795: dataIn1 = 32'd600
; 
32'd24796: dataIn1 = 32'd604
; 
32'd24797: dataIn1 = 32'd614
; 
32'd24798: dataIn1 = 32'd618
; 
32'd24799: dataIn1 = 32'd620
; 
32'd24800: dataIn1 = 32'd633
; 
32'd24801: dataIn1 = 32'd637
; 
32'd24802: dataIn1 = 32'd642
; 
32'd24803: dataIn1 = 32'd683
; 
32'd24804: dataIn1 = 32'd702
; 
32'd24805: dataIn1 = 32'd720
; 
32'd24806: dataIn1 = 32'd725
; 
32'd24807: dataIn1 = 32'd742
; 
32'd24808: dataIn1 = 32'd758
; 
32'd24809: dataIn1 = 32'd759
; 
32'd24810: dataIn1 = 32'd789
; 
32'd24811: dataIn1 = 32'd526
; 
32'd24812: dataIn1 = 32'd529
; 
32'd24813: dataIn1 = 32'd534
; 
32'd24814: dataIn1 = 32'd547
; 
32'd24815: dataIn1 = 32'd551
; 
32'd24816: dataIn1 = 32'd558
; 
32'd24817: dataIn1 = 32'd573
; 
32'd24818: dataIn1 = 32'd580
; 
32'd24819: dataIn1 = 32'd585
; 
32'd24820: dataIn1 = 32'd587
; 
32'd24821: dataIn1 = 32'd593
; 
32'd24822: dataIn1 = 32'd599
; 
32'd24823: dataIn1 = 32'd636
; 
32'd24824: dataIn1 = 32'd656
; 
32'd24825: dataIn1 = 32'd680
; 
32'd24826: dataIn1 = 32'd683
; 
32'd24827: dataIn1 = 32'd695
; 
32'd24828: dataIn1 = 32'd699
; 
32'd24829: dataIn1 = 32'd700
; 
32'd24830: dataIn1 = 32'd714
; 
32'd24831: dataIn1 = 32'd718
; 
32'd24832: dataIn1 = 32'd753
; 
32'd24833: dataIn1 = 32'd786
; 
32'd24834: dataIn1 = 32'd791
; 
32'd24835: dataIn1 = 32'd793
; 
32'd24836: dataIn1 = 32'd545
; 
32'd24837: dataIn1 = 32'd579
; 
32'd24838: dataIn1 = 32'd602
; 
32'd24839: dataIn1 = 32'd623
; 
32'd24840: dataIn1 = 32'd634
; 
32'd24841: dataIn1 = 32'd671
; 
32'd24842: dataIn1 = 32'd699
; 
32'd24843: dataIn1 = 32'd701
; 
32'd24844: dataIn1 = 32'd715
; 
32'd24845: dataIn1 = 32'd728
; 
32'd24846: dataIn1 = 32'd743
; 
32'd24847: dataIn1 = 32'd521
; 
32'd24848: dataIn1 = 32'd529
; 
32'd24849: dataIn1 = 32'd534
; 
32'd24850: dataIn1 = 32'd540
; 
32'd24851: dataIn1 = 32'd547
; 
32'd24852: dataIn1 = 32'd556
; 
32'd24853: dataIn1 = 32'd607
; 
32'd24854: dataIn1 = 32'd648
; 
32'd24855: dataIn1 = 32'd658
; 
32'd24856: dataIn1 = 32'd675
; 
32'd24857: dataIn1 = 32'd680
; 
32'd24858: dataIn1 = 32'd701
; 
32'd24859: dataIn1 = 32'd738
; 
32'd24860: dataIn1 = 32'd742
; 
32'd24861: dataIn1 = 32'd754
; 
32'd24862: dataIn1 = 32'd762
; 
32'd24863: dataIn1 = 32'd768
; 
32'd24864: dataIn1 = 32'd769
; 
32'd24865: dataIn1 = 32'd779
; 
32'd24866: dataIn1 = 32'd521
; 
32'd24867: dataIn1 = 32'd538
; 
32'd24868: dataIn1 = 32'd555
; 
32'd24869: dataIn1 = 32'd569
; 
32'd24870: dataIn1 = 32'd570
; 
32'd24871: dataIn1 = 32'd572
; 
32'd24872: dataIn1 = 32'd628
; 
32'd24873: dataIn1 = 32'd631
; 
32'd24874: dataIn1 = 32'd641
; 
32'd24875: dataIn1 = 32'd659
; 
32'd24876: dataIn1 = 32'd673
; 
32'd24877: dataIn1 = 32'd694
; 
32'd24878: dataIn1 = 32'd697
; 
32'd24879: dataIn1 = 32'd718
; 
32'd24880: dataIn1 = 32'd722
; 
32'd24881: dataIn1 = 32'd748
; 
32'd24882: dataIn1 = 32'd758
; 
32'd24883: dataIn1 = 32'd761
; 
32'd24884: dataIn1 = 32'd767
; 
32'd24885: dataIn1 = 32'd800
; 
32'd24886: dataIn1 = 32'd527
; 
32'd24887: dataIn1 = 32'd528
; 
32'd24888: dataIn1 = 32'd531
; 
32'd24889: dataIn1 = 32'd548
; 
32'd24890: dataIn1 = 32'd556
; 
32'd24891: dataIn1 = 32'd579
; 
32'd24892: dataIn1 = 32'd614
; 
32'd24893: dataIn1 = 32'd624
; 
32'd24894: dataIn1 = 32'd656
; 
32'd24895: dataIn1 = 32'd671
; 
32'd24896: dataIn1 = 32'd734
; 
32'd24897: dataIn1 = 32'd786
; 
32'd24898: dataIn1 = 32'd796
; 
32'd24899: dataIn1 = 32'd799
; 
32'd24900: dataIn1 = 32'd534
; 
32'd24901: dataIn1 = 32'd586
; 
32'd24902: dataIn1 = 32'd598
; 
32'd24903: dataIn1 = 32'd604
; 
32'd24904: dataIn1 = 32'd618
; 
32'd24905: dataIn1 = 32'd622
; 
32'd24906: dataIn1 = 32'd624
; 
32'd24907: dataIn1 = 32'd628
; 
32'd24908: dataIn1 = 32'd648
; 
32'd24909: dataIn1 = 32'd659
; 
32'd24910: dataIn1 = 32'd661
; 
32'd24911: dataIn1 = 32'd674
; 
32'd24912: dataIn1 = 32'd734
; 
32'd24913: dataIn1 = 32'd737
; 
32'd24914: dataIn1 = 32'd738
; 
32'd24915: dataIn1 = 32'd747
; 
32'd24916: dataIn1 = 32'd770
; 
32'd24917: dataIn1 = 32'd789
; 
32'd24918: dataIn1 = 32'd525
; 
32'd24919: dataIn1 = 32'd541
; 
32'd24920: dataIn1 = 32'd549
; 
32'd24921: dataIn1 = 32'd565
; 
32'd24922: dataIn1 = 32'd577
; 
32'd24923: dataIn1 = 32'd582
; 
32'd24924: dataIn1 = 32'd588
; 
32'd24925: dataIn1 = 32'd635
; 
32'd24926: dataIn1 = 32'd637
; 
32'd24927: dataIn1 = 32'd652
; 
32'd24928: dataIn1 = 32'd667
; 
32'd24929: dataIn1 = 32'd721
; 
32'd24930: dataIn1 = 32'd726
; 
32'd24931: dataIn1 = 32'd749
; 
32'd24932: dataIn1 = 32'd761
; 
32'd24933: dataIn1 = 32'd762
; 
32'd24934: dataIn1 = 32'd771
; 
32'd24935: dataIn1 = 32'd773
; 
32'd24936: dataIn1 = 32'd799
; 
32'd24937: dataIn1 = 32'd529
; 
32'd24938: dataIn1 = 32'd536
; 
32'd24939: dataIn1 = 32'd541
; 
32'd24940: dataIn1 = 32'd552
; 
32'd24941: dataIn1 = 32'd556
; 
32'd24942: dataIn1 = 32'd600
; 
32'd24943: dataIn1 = 32'd666
; 
32'd24944: dataIn1 = 32'd669
; 
32'd24945: dataIn1 = 32'd717
; 
32'd24946: dataIn1 = 32'd741
; 
32'd24947: dataIn1 = 32'd749
; 
32'd24948: dataIn1 = 32'd755
; 
32'd24949: dataIn1 = 32'd794
; 
32'd24950: dataIn1 = 32'd526
; 
32'd24951: dataIn1 = 32'd532
; 
32'd24952: dataIn1 = 32'd539
; 
32'd24953: dataIn1 = 32'd540
; 
32'd24954: dataIn1 = 32'd566
; 
32'd24955: dataIn1 = 32'd588
; 
32'd24956: dataIn1 = 32'd598
; 
32'd24957: dataIn1 = 32'd610
; 
32'd24958: dataIn1 = 32'd615
; 
32'd24959: dataIn1 = 32'd631
; 
32'd24960: dataIn1 = 32'd636
; 
32'd24961: dataIn1 = 32'd642
; 
32'd24962: dataIn1 = 32'd684
; 
32'd24963: dataIn1 = 32'd696
; 
32'd24964: dataIn1 = 32'd704
; 
32'd24965: dataIn1 = 32'd764
; 
32'd24966: dataIn1 = 32'd776
; 
32'd24967: dataIn1 = 32'd779
; 
32'd24968: dataIn1 = 32'd793
; 
32'd24969: dataIn1 = 32'd539
; 
32'd24970: dataIn1 = 32'd541
; 
32'd24971: dataIn1 = 32'd547
; 
32'd24972: dataIn1 = 32'd552
; 
32'd24973: dataIn1 = 32'd570
; 
32'd24974: dataIn1 = 32'd580
; 
32'd24975: dataIn1 = 32'd595
; 
32'd24976: dataIn1 = 32'd632
; 
32'd24977: dataIn1 = 32'd640
; 
32'd24978: dataIn1 = 32'd647
; 
32'd24979: dataIn1 = 32'd697
; 
32'd24980: dataIn1 = 32'd703
; 
32'd24981: dataIn1 = 32'd726
; 
32'd24982: dataIn1 = 32'd743
; 
32'd24983: dataIn1 = 32'd747
; 
32'd24984: dataIn1 = 32'd770
; 
32'd24985: dataIn1 = 32'd533
; 
32'd24986: dataIn1 = 32'd564
; 
32'd24987: dataIn1 = 32'd567
; 
32'd24988: dataIn1 = 32'd586
; 
32'd24989: dataIn1 = 32'd594
; 
32'd24990: dataIn1 = 32'd595
; 
32'd24991: dataIn1 = 32'd635
; 
32'd24992: dataIn1 = 32'd658
; 
32'd24993: dataIn1 = 32'd668
; 
32'd24994: dataIn1 = 32'd714
; 
32'd24995: dataIn1 = 32'd720
; 
32'd24996: dataIn1 = 32'd769
; 
32'd24997: dataIn1 = 32'd548
; 
32'd24998: dataIn1 = 32'd561
; 
32'd24999: dataIn1 = 32'd578
; 
32'd25000: dataIn1 = 32'd587
; 
32'd25001: dataIn1 = 32'd592
; 
32'd25002: dataIn1 = 32'd612
; 
32'd25003: dataIn1 = 32'd619
; 
32'd25004: dataIn1 = 32'd648
; 
32'd25005: dataIn1 = 32'd652
; 
32'd25006: dataIn1 = 32'd665
; 
32'd25007: dataIn1 = 32'd693
; 
32'd25008: dataIn1 = 32'd710
; 
32'd25009: dataIn1 = 32'd721
; 
32'd25010: dataIn1 = 32'd742
; 
32'd25011: dataIn1 = 32'd745
; 
32'd25012: dataIn1 = 32'd781
; 
32'd25013: dataIn1 = 32'd783
; 
32'd25014: dataIn1 = 32'd787
; 
32'd25015: dataIn1 = 32'd532
; 
32'd25016: dataIn1 = 32'd546
; 
32'd25017: dataIn1 = 32'd548
; 
32'd25018: dataIn1 = 32'd552
; 
32'd25019: dataIn1 = 32'd573
; 
32'd25020: dataIn1 = 32'd579
; 
32'd25021: dataIn1 = 32'd616
; 
32'd25022: dataIn1 = 32'd628
; 
32'd25023: dataIn1 = 32'd629
; 
32'd25024: dataIn1 = 32'd648
; 
32'd25025: dataIn1 = 32'd678
; 
32'd25026: dataIn1 = 32'd714
; 
32'd25027: dataIn1 = 32'd718
; 
32'd25028: dataIn1 = 32'd724
; 
32'd25029: dataIn1 = 32'd728
; 
32'd25030: dataIn1 = 32'd734
; 
32'd25031: dataIn1 = 32'd754
; 
32'd25032: dataIn1 = 32'd766
; 
32'd25033: dataIn1 = 32'd777
; 
32'd25034: dataIn1 = 32'd536
; 
32'd25035: dataIn1 = 32'd556
; 
32'd25036: dataIn1 = 32'd565
; 
32'd25037: dataIn1 = 32'd643
; 
32'd25038: dataIn1 = 32'd656
; 
32'd25039: dataIn1 = 32'd658
; 
32'd25040: dataIn1 = 32'd680
; 
32'd25041: dataIn1 = 32'd683
; 
32'd25042: dataIn1 = 32'd685
; 
32'd25043: dataIn1 = 32'd699
; 
32'd25044: dataIn1 = 32'd728
; 
32'd25045: dataIn1 = 32'd758
; 
32'd25046: dataIn1 = 32'd778
; 
32'd25047: dataIn1 = 32'd800
; 
32'd25048: dataIn1 = 32'd554
; 
32'd25049: dataIn1 = 32'd555
; 
32'd25050: dataIn1 = 32'd558
; 
32'd25051: dataIn1 = 32'd566
; 
32'd25052: dataIn1 = 32'd575
; 
32'd25053: dataIn1 = 32'd577
; 
32'd25054: dataIn1 = 32'd595
; 
32'd25055: dataIn1 = 32'd609
; 
32'd25056: dataIn1 = 32'd665
; 
32'd25057: dataIn1 = 32'd696
; 
32'd25058: dataIn1 = 32'd721
; 
32'd25059: dataIn1 = 32'd725
; 
32'd25060: dataIn1 = 32'd733
; 
32'd25061: dataIn1 = 32'd752
; 
32'd25062: dataIn1 = 32'd797
; 
32'd25063: dataIn1 = 32'd799
; 
32'd25064: dataIn1 = 32'd541
; 
32'd25065: dataIn1 = 32'd556
; 
32'd25066: dataIn1 = 32'd562
; 
32'd25067: dataIn1 = 32'd580
; 
32'd25068: dataIn1 = 32'd604
; 
32'd25069: dataIn1 = 32'd614
; 
32'd25070: dataIn1 = 32'd635
; 
32'd25071: dataIn1 = 32'd641
; 
32'd25072: dataIn1 = 32'd657
; 
32'd25073: dataIn1 = 32'd662
; 
32'd25074: dataIn1 = 32'd718
; 
32'd25075: dataIn1 = 32'd763
; 
32'd25076: dataIn1 = 32'd784
; 
32'd25077: dataIn1 = 32'd534
; 
32'd25078: dataIn1 = 32'd564
; 
32'd25079: dataIn1 = 32'd584
; 
32'd25080: dataIn1 = 32'd596
; 
32'd25081: dataIn1 = 32'd607
; 
32'd25082: dataIn1 = 32'd609
; 
32'd25083: dataIn1 = 32'd628
; 
32'd25084: dataIn1 = 32'd639
; 
32'd25085: dataIn1 = 32'd643
; 
32'd25086: dataIn1 = 32'd651
; 
32'd25087: dataIn1 = 32'd679
; 
32'd25088: dataIn1 = 32'd684
; 
32'd25089: dataIn1 = 32'd685
; 
32'd25090: dataIn1 = 32'd687
; 
32'd25091: dataIn1 = 32'd695
; 
32'd25092: dataIn1 = 32'd705
; 
32'd25093: dataIn1 = 32'd707
; 
32'd25094: dataIn1 = 32'd719
; 
32'd25095: dataIn1 = 32'd720
; 
32'd25096: dataIn1 = 32'd786
; 
32'd25097: dataIn1 = 32'd548
; 
32'd25098: dataIn1 = 32'd550
; 
32'd25099: dataIn1 = 32'd630
; 
32'd25100: dataIn1 = 32'd682
; 
32'd25101: dataIn1 = 32'd690
; 
32'd25102: dataIn1 = 32'd695
; 
32'd25103: dataIn1 = 32'd696
; 
32'd25104: dataIn1 = 32'd701
; 
32'd25105: dataIn1 = 32'd729
; 
32'd25106: dataIn1 = 32'd740
; 
32'd25107: dataIn1 = 32'd745
; 
32'd25108: dataIn1 = 32'd766
; 
32'd25109: dataIn1 = 32'd772
; 
32'd25110: dataIn1 = 32'd540
; 
32'd25111: dataIn1 = 32'd541
; 
32'd25112: dataIn1 = 32'd572
; 
32'd25113: dataIn1 = 32'd619
; 
32'd25114: dataIn1 = 32'd633
; 
32'd25115: dataIn1 = 32'd655
; 
32'd25116: dataIn1 = 32'd669
; 
32'd25117: dataIn1 = 32'd677
; 
32'd25118: dataIn1 = 32'd693
; 
32'd25119: dataIn1 = 32'd721
; 
32'd25120: dataIn1 = 32'd723
; 
32'd25121: dataIn1 = 32'd785
; 
32'd25122: dataIn1 = 32'd560
; 
32'd25123: dataIn1 = 32'd587
; 
32'd25124: dataIn1 = 32'd600
; 
32'd25125: dataIn1 = 32'd603
; 
32'd25126: dataIn1 = 32'd604
; 
32'd25127: dataIn1 = 32'd610
; 
32'd25128: dataIn1 = 32'd619
; 
32'd25129: dataIn1 = 32'd624
; 
32'd25130: dataIn1 = 32'd636
; 
32'd25131: dataIn1 = 32'd640
; 
32'd25132: dataIn1 = 32'd651
; 
32'd25133: dataIn1 = 32'd669
; 
32'd25134: dataIn1 = 32'd714
; 
32'd25135: dataIn1 = 32'd740
; 
32'd25136: dataIn1 = 32'd744
; 
32'd25137: dataIn1 = 32'd747
; 
32'd25138: dataIn1 = 32'd751
; 
32'd25139: dataIn1 = 32'd771
; 
32'd25140: dataIn1 = 32'd772
; 
32'd25141: dataIn1 = 32'd787
; 
32'd25142: dataIn1 = 32'd542
; 
32'd25143: dataIn1 = 32'd545
; 
32'd25144: dataIn1 = 32'd581
; 
32'd25145: dataIn1 = 32'd600
; 
32'd25146: dataIn1 = 32'd619
; 
32'd25147: dataIn1 = 32'd643
; 
32'd25148: dataIn1 = 32'd659
; 
32'd25149: dataIn1 = 32'd664
; 
32'd25150: dataIn1 = 32'd693
; 
32'd25151: dataIn1 = 32'd740
; 
32'd25152: dataIn1 = 32'd762
; 
32'd25153: dataIn1 = 32'd796
; 
32'd25154: dataIn1 = 32'd555
; 
32'd25155: dataIn1 = 32'd560
; 
32'd25156: dataIn1 = 32'd563
; 
32'd25157: dataIn1 = 32'd573
; 
32'd25158: dataIn1 = 32'd583
; 
32'd25159: dataIn1 = 32'd597
; 
32'd25160: dataIn1 = 32'd599
; 
32'd25161: dataIn1 = 32'd626
; 
32'd25162: dataIn1 = 32'd683
; 
32'd25163: dataIn1 = 32'd700
; 
32'd25164: dataIn1 = 32'd712
; 
32'd25165: dataIn1 = 32'd741
; 
32'd25166: dataIn1 = 32'd742
; 
32'd25167: dataIn1 = 32'd776
; 
32'd25168: dataIn1 = 32'd790
; 
32'd25169: dataIn1 = 32'd792
; 
32'd25170: dataIn1 = 32'd557
; 
32'd25171: dataIn1 = 32'd581
; 
32'd25172: dataIn1 = 32'd586
; 
32'd25173: dataIn1 = 32'd601
; 
32'd25174: dataIn1 = 32'd606
; 
32'd25175: dataIn1 = 32'd630
; 
32'd25176: dataIn1 = 32'd638
; 
32'd25177: dataIn1 = 32'd646
; 
32'd25178: dataIn1 = 32'd653
; 
32'd25179: dataIn1 = 32'd663
; 
32'd25180: dataIn1 = 32'd675
; 
32'd25181: dataIn1 = 32'd714
; 
32'd25182: dataIn1 = 32'd751
; 
32'd25183: dataIn1 = 32'd756
; 
32'd25184: dataIn1 = 32'd776
; 
32'd25185: dataIn1 = 32'd778
; 
32'd25186: dataIn1 = 32'd789
; 
32'd25187: dataIn1 = 32'd790
; 
32'd25188: dataIn1 = 32'd793
; 
32'd25189: dataIn1 = 32'd549
; 
32'd25190: dataIn1 = 32'd583
; 
32'd25191: dataIn1 = 32'd596
; 
32'd25192: dataIn1 = 32'd606
; 
32'd25193: dataIn1 = 32'd614
; 
32'd25194: dataIn1 = 32'd617
; 
32'd25195: dataIn1 = 32'd644
; 
32'd25196: dataIn1 = 32'd649
; 
32'd25197: dataIn1 = 32'd652
; 
32'd25198: dataIn1 = 32'd661
; 
32'd25199: dataIn1 = 32'd723
; 
32'd25200: dataIn1 = 32'd746
; 
32'd25201: dataIn1 = 32'd550
; 
32'd25202: dataIn1 = 32'd560
; 
32'd25203: dataIn1 = 32'd573
; 
32'd25204: dataIn1 = 32'd653
; 
32'd25205: dataIn1 = 32'd655
; 
32'd25206: dataIn1 = 32'd783
; 
32'd25207: dataIn1 = 32'd793
; 
32'd25208: dataIn1 = 32'd544
; 
32'd25209: dataIn1 = 32'd546
; 
32'd25210: dataIn1 = 32'd549
; 
32'd25211: dataIn1 = 32'd570
; 
32'd25212: dataIn1 = 32'd586
; 
32'd25213: dataIn1 = 32'd616
; 
32'd25214: dataIn1 = 32'd625
; 
32'd25215: dataIn1 = 32'd633
; 
32'd25216: dataIn1 = 32'd648
; 
32'd25217: dataIn1 = 32'd654
; 
32'd25218: dataIn1 = 32'd677
; 
32'd25219: dataIn1 = 32'd706
; 
32'd25220: dataIn1 = 32'd739
; 
32'd25221: dataIn1 = 32'd751
; 
32'd25222: dataIn1 = 32'd762
; 
32'd25223: dataIn1 = 32'd778
; 
32'd25224: dataIn1 = 32'd551
; 
32'd25225: dataIn1 = 32'd564
; 
32'd25226: dataIn1 = 32'd574
; 
32'd25227: dataIn1 = 32'd575
; 
32'd25228: dataIn1 = 32'd603
; 
32'd25229: dataIn1 = 32'd604
; 
32'd25230: dataIn1 = 32'd626
; 
32'd25231: dataIn1 = 32'd631
; 
32'd25232: dataIn1 = 32'd636
; 
32'd25233: dataIn1 = 32'd649
; 
32'd25234: dataIn1 = 32'd651
; 
32'd25235: dataIn1 = 32'd661
; 
32'd25236: dataIn1 = 32'd689
; 
32'd25237: dataIn1 = 32'd705
; 
32'd25238: dataIn1 = 32'd729
; 
32'd25239: dataIn1 = 32'd768
; 
32'd25240: dataIn1 = 32'd788
; 
32'd25241: dataIn1 = 32'd565
; 
32'd25242: dataIn1 = 32'd583
; 
32'd25243: dataIn1 = 32'd592
; 
32'd25244: dataIn1 = 32'd607
; 
32'd25245: dataIn1 = 32'd632
; 
32'd25246: dataIn1 = 32'd658
; 
32'd25247: dataIn1 = 32'd674
; 
32'd25248: dataIn1 = 32'd728
; 
32'd25249: dataIn1 = 32'd729
; 
32'd25250: dataIn1 = 32'd732
; 
32'd25251: dataIn1 = 32'd749
; 
32'd25252: dataIn1 = 32'd765
; 
32'd25253: dataIn1 = 32'd785
; 
32'd25254: dataIn1 = 32'd576
; 
32'd25255: dataIn1 = 32'd600
; 
32'd25256: dataIn1 = 32'd616
; 
32'd25257: dataIn1 = 32'd638
; 
32'd25258: dataIn1 = 32'd664
; 
32'd25259: dataIn1 = 32'd702
; 
32'd25260: dataIn1 = 32'd706
; 
32'd25261: dataIn1 = 32'd719
; 
32'd25262: dataIn1 = 32'd730
; 
32'd25263: dataIn1 = 32'd749
; 
32'd25264: dataIn1 = 32'd781
; 
32'd25265: dataIn1 = 32'd793
; 
32'd25266: dataIn1 = 32'd565
; 
32'd25267: dataIn1 = 32'd575
; 
32'd25268: dataIn1 = 32'd579
; 
32'd25269: dataIn1 = 32'd600
; 
32'd25270: dataIn1 = 32'd614
; 
32'd25271: dataIn1 = 32'd619
; 
32'd25272: dataIn1 = 32'd631
; 
32'd25273: dataIn1 = 32'd660
; 
32'd25274: dataIn1 = 32'd661
; 
32'd25275: dataIn1 = 32'd672
; 
32'd25276: dataIn1 = 32'd674
; 
32'd25277: dataIn1 = 32'd678
; 
32'd25278: dataIn1 = 32'd690
; 
32'd25279: dataIn1 = 32'd695
; 
32'd25280: dataIn1 = 32'd700
; 
32'd25281: dataIn1 = 32'd704
; 
32'd25282: dataIn1 = 32'd737
; 
32'd25283: dataIn1 = 32'd757
; 
32'd25284: dataIn1 = 32'd787
; 
32'd25285: dataIn1 = 32'd788
; 
32'd25286: dataIn1 = 32'd555
; 
32'd25287: dataIn1 = 32'd556
; 
32'd25288: dataIn1 = 32'd561
; 
32'd25289: dataIn1 = 32'd566
; 
32'd25290: dataIn1 = 32'd581
; 
32'd25291: dataIn1 = 32'd646
; 
32'd25292: dataIn1 = 32'd648
; 
32'd25293: dataIn1 = 32'd655
; 
32'd25294: dataIn1 = 32'd772
; 
32'd25295: dataIn1 = 32'd774
; 
32'd25296: dataIn1 = 32'd777
; 
32'd25297: dataIn1 = 32'd786
; 
32'd25298: dataIn1 = 32'd789
; 
32'd25299: dataIn1 = 32'd791
; 
32'd25300: dataIn1 = 32'd792
; 
32'd25301: dataIn1 = 32'd568
; 
32'd25302: dataIn1 = 32'd571
; 
32'd25303: dataIn1 = 32'd578
; 
32'd25304: dataIn1 = 32'd584
; 
32'd25305: dataIn1 = 32'd598
; 
32'd25306: dataIn1 = 32'd600
; 
32'd25307: dataIn1 = 32'd608
; 
32'd25308: dataIn1 = 32'd615
; 
32'd25309: dataIn1 = 32'd618
; 
32'd25310: dataIn1 = 32'd682
; 
32'd25311: dataIn1 = 32'd691
; 
32'd25312: dataIn1 = 32'd703
; 
32'd25313: dataIn1 = 32'd735
; 
32'd25314: dataIn1 = 32'd758
; 
32'd25315: dataIn1 = 32'd798
; 
32'd25316: dataIn1 = 32'd558
; 
32'd25317: dataIn1 = 32'd563
; 
32'd25318: dataIn1 = 32'd581
; 
32'd25319: dataIn1 = 32'd605
; 
32'd25320: dataIn1 = 32'd617
; 
32'd25321: dataIn1 = 32'd622
; 
32'd25322: dataIn1 = 32'd634
; 
32'd25323: dataIn1 = 32'd657
; 
32'd25324: dataIn1 = 32'd682
; 
32'd25325: dataIn1 = 32'd683
; 
32'd25326: dataIn1 = 32'd693
; 
32'd25327: dataIn1 = 32'd698
; 
32'd25328: dataIn1 = 32'd713
; 
32'd25329: dataIn1 = 32'd714
; 
32'd25330: dataIn1 = 32'd722
; 
32'd25331: dataIn1 = 32'd729
; 
32'd25332: dataIn1 = 32'd732
; 
32'd25333: dataIn1 = 32'd762
; 
32'd25334: dataIn1 = 32'd765
; 
32'd25335: dataIn1 = 32'd564
; 
32'd25336: dataIn1 = 32'd572
; 
32'd25337: dataIn1 = 32'd574
; 
32'd25338: dataIn1 = 32'd579
; 
32'd25339: dataIn1 = 32'd610
; 
32'd25340: dataIn1 = 32'd702
; 
32'd25341: dataIn1 = 32'd712
; 
32'd25342: dataIn1 = 32'd724
; 
32'd25343: dataIn1 = 32'd729
; 
32'd25344: dataIn1 = 32'd738
; 
32'd25345: dataIn1 = 32'd743
; 
32'd25346: dataIn1 = 32'd760
; 
32'd25347: dataIn1 = 32'd773
; 
32'd25348: dataIn1 = 32'd774
; 
32'd25349: dataIn1 = 32'd565
; 
32'd25350: dataIn1 = 32'd571
; 
32'd25351: dataIn1 = 32'd581
; 
32'd25352: dataIn1 = 32'd591
; 
32'd25353: dataIn1 = 32'd609
; 
32'd25354: dataIn1 = 32'd612
; 
32'd25355: dataIn1 = 32'd626
; 
32'd25356: dataIn1 = 32'd647
; 
32'd25357: dataIn1 = 32'd648
; 
32'd25358: dataIn1 = 32'd672
; 
32'd25359: dataIn1 = 32'd691
; 
32'd25360: dataIn1 = 32'd742
; 
32'd25361: dataIn1 = 32'd763
; 
32'd25362: dataIn1 = 32'd791
; 
32'd25363: dataIn1 = 32'd562
; 
32'd25364: dataIn1 = 32'd568
; 
32'd25365: dataIn1 = 32'd572
; 
32'd25366: dataIn1 = 32'd581
; 
32'd25367: dataIn1 = 32'd582
; 
32'd25368: dataIn1 = 32'd633
; 
32'd25369: dataIn1 = 32'd641
; 
32'd25370: dataIn1 = 32'd643
; 
32'd25371: dataIn1 = 32'd671
; 
32'd25372: dataIn1 = 32'd695
; 
32'd25373: dataIn1 = 32'd706
; 
32'd25374: dataIn1 = 32'd720
; 
32'd25375: dataIn1 = 32'd728
; 
32'd25376: dataIn1 = 32'd759
; 
32'd25377: dataIn1 = 32'd782
; 
32'd25378: dataIn1 = 32'd788
; 
32'd25379: dataIn1 = 32'd584
; 
32'd25380: dataIn1 = 32'd598
; 
32'd25381: dataIn1 = 32'd607
; 
32'd25382: dataIn1 = 32'd654
; 
32'd25383: dataIn1 = 32'd677
; 
32'd25384: dataIn1 = 32'd686
; 
32'd25385: dataIn1 = 32'd722
; 
32'd25386: dataIn1 = 32'd737
; 
32'd25387: dataIn1 = 32'd740
; 
32'd25388: dataIn1 = 32'd742
; 
32'd25389: dataIn1 = 32'd756
; 
32'd25390: dataIn1 = 32'd762
; 
32'd25391: dataIn1 = 32'd793
; 
32'd25392: dataIn1 = 32'd796
; 
32'd25393: dataIn1 = 32'd590
; 
32'd25394: dataIn1 = 32'd601
; 
32'd25395: dataIn1 = 32'd656
; 
32'd25396: dataIn1 = 32'd669
; 
32'd25397: dataIn1 = 32'd687
; 
32'd25398: dataIn1 = 32'd700
; 
32'd25399: dataIn1 = 32'd719
; 
32'd25400: dataIn1 = 32'd728
; 
32'd25401: dataIn1 = 32'd753
; 
32'd25402: dataIn1 = 32'd776
; 
32'd25403: dataIn1 = 32'd799
; 
32'd25404: dataIn1 = 32'd628
; 
32'd25405: dataIn1 = 32'd642
; 
32'd25406: dataIn1 = 32'd653
; 
32'd25407: dataIn1 = 32'd684
; 
32'd25408: dataIn1 = 32'd704
; 
32'd25409: dataIn1 = 32'd742
; 
32'd25410: dataIn1 = 32'd752
; 
32'd25411: dataIn1 = 32'd766
; 
32'd25412: dataIn1 = 32'd772
; 
32'd25413: dataIn1 = 32'd557
; 
32'd25414: dataIn1 = 32'd558
; 
32'd25415: dataIn1 = 32'd576
; 
32'd25416: dataIn1 = 32'd579
; 
32'd25417: dataIn1 = 32'd616
; 
32'd25418: dataIn1 = 32'd655
; 
32'd25419: dataIn1 = 32'd659
; 
32'd25420: dataIn1 = 32'd663
; 
32'd25421: dataIn1 = 32'd674
; 
32'd25422: dataIn1 = 32'd677
; 
32'd25423: dataIn1 = 32'd686
; 
32'd25424: dataIn1 = 32'd688
; 
32'd25425: dataIn1 = 32'd705
; 
32'd25426: dataIn1 = 32'd721
; 
32'd25427: dataIn1 = 32'd734
; 
32'd25428: dataIn1 = 32'd760
; 
32'd25429: dataIn1 = 32'd794
; 
32'd25430: dataIn1 = 32'd800
; 
32'd25431: dataIn1 = 32'd567
; 
32'd25432: dataIn1 = 32'd582
; 
32'd25433: dataIn1 = 32'd590
; 
32'd25434: dataIn1 = 32'd591
; 
32'd25435: dataIn1 = 32'd608
; 
32'd25436: dataIn1 = 32'd629
; 
32'd25437: dataIn1 = 32'd644
; 
32'd25438: dataIn1 = 32'd688
; 
32'd25439: dataIn1 = 32'd694
; 
32'd25440: dataIn1 = 32'd701
; 
32'd25441: dataIn1 = 32'd712
; 
32'd25442: dataIn1 = 32'd713
; 
32'd25443: dataIn1 = 32'd714
; 
32'd25444: dataIn1 = 32'd719
; 
32'd25445: dataIn1 = 32'd784
; 
32'd25446: dataIn1 = 32'd793
; 
32'd25447: dataIn1 = 32'd798
; 
32'd25448: dataIn1 = 32'd585
; 
32'd25449: dataIn1 = 32'd586
; 
32'd25450: dataIn1 = 32'd597
; 
32'd25451: dataIn1 = 32'd616
; 
32'd25452: dataIn1 = 32'd620
; 
32'd25453: dataIn1 = 32'd635
; 
32'd25454: dataIn1 = 32'd652
; 
32'd25455: dataIn1 = 32'd660
; 
32'd25456: dataIn1 = 32'd735
; 
32'd25457: dataIn1 = 32'd741
; 
32'd25458: dataIn1 = 32'd773
; 
32'd25459: dataIn1 = 32'd785
; 
32'd25460: dataIn1 = 32'd799
; 
32'd25461: dataIn1 = 32'd565
; 
32'd25462: dataIn1 = 32'd600
; 
32'd25463: dataIn1 = 32'd605
; 
32'd25464: dataIn1 = 32'd609
; 
32'd25465: dataIn1 = 32'd622
; 
32'd25466: dataIn1 = 32'd650
; 
32'd25467: dataIn1 = 32'd683
; 
32'd25468: dataIn1 = 32'd719
; 
32'd25469: dataIn1 = 32'd736
; 
32'd25470: dataIn1 = 32'd739
; 
32'd25471: dataIn1 = 32'd753
; 
32'd25472: dataIn1 = 32'd769
; 
32'd25473: dataIn1 = 32'd773
; 
32'd25474: dataIn1 = 32'd775
; 
32'd25475: dataIn1 = 32'd563
; 
32'd25476: dataIn1 = 32'd586
; 
32'd25477: dataIn1 = 32'd596
; 
32'd25478: dataIn1 = 32'd636
; 
32'd25479: dataIn1 = 32'd639
; 
32'd25480: dataIn1 = 32'd702
; 
32'd25481: dataIn1 = 32'd734
; 
32'd25482: dataIn1 = 32'd749
; 
32'd25483: dataIn1 = 32'd759
; 
32'd25484: dataIn1 = 32'd772
; 
32'd25485: dataIn1 = 32'd785
; 
32'd25486: dataIn1 = 32'd793
; 
32'd25487: dataIn1 = 32'd796
; 
32'd25488: dataIn1 = 32'd569
; 
32'd25489: dataIn1 = 32'd572
; 
32'd25490: dataIn1 = 32'd578
; 
32'd25491: dataIn1 = 32'd583
; 
32'd25492: dataIn1 = 32'd586
; 
32'd25493: dataIn1 = 32'd601
; 
32'd25494: dataIn1 = 32'd632
; 
32'd25495: dataIn1 = 32'd681
; 
32'd25496: dataIn1 = 32'd682
; 
32'd25497: dataIn1 = 32'd687
; 
32'd25498: dataIn1 = 32'd699
; 
32'd25499: dataIn1 = 32'd704
; 
32'd25500: dataIn1 = 32'd730
; 
32'd25501: dataIn1 = 32'd751
; 
32'd25502: dataIn1 = 32'd759
; 
32'd25503: dataIn1 = 32'd762
; 
32'd25504: dataIn1 = 32'd776
; 
32'd25505: dataIn1 = 32'd784
; 
32'd25506: dataIn1 = 32'd567
; 
32'd25507: dataIn1 = 32'd568
; 
32'd25508: dataIn1 = 32'd663
; 
32'd25509: dataIn1 = 32'd667
; 
32'd25510: dataIn1 = 32'd706
; 
32'd25511: dataIn1 = 32'd721
; 
32'd25512: dataIn1 = 32'd737
; 
32'd25513: dataIn1 = 32'd748
; 
32'd25514: dataIn1 = 32'd757
; 
32'd25515: dataIn1 = 32'd758
; 
32'd25516: dataIn1 = 32'd789
; 
32'd25517: dataIn1 = 32'd794
; 
32'd25518: dataIn1 = 32'd586
; 
32'd25519: dataIn1 = 32'd591
; 
32'd25520: dataIn1 = 32'd592
; 
32'd25521: dataIn1 = 32'd597
; 
32'd25522: dataIn1 = 32'd600
; 
32'd25523: dataIn1 = 32'd606
; 
32'd25524: dataIn1 = 32'd638
; 
32'd25525: dataIn1 = 32'd714
; 
32'd25526: dataIn1 = 32'd718
; 
32'd25527: dataIn1 = 32'd724
; 
32'd25528: dataIn1 = 32'd729
; 
32'd25529: dataIn1 = 32'd745
; 
32'd25530: dataIn1 = 32'd765
; 
32'd25531: dataIn1 = 32'd782
; 
32'd25532: dataIn1 = 32'd784
; 
32'd25533: dataIn1 = 32'd800
; 
32'd25534: dataIn1 = 32'd567
; 
32'd25535: dataIn1 = 32'd572
; 
32'd25536: dataIn1 = 32'd611
; 
32'd25537: dataIn1 = 32'd618
; 
32'd25538: dataIn1 = 32'd635
; 
32'd25539: dataIn1 = 32'd640
; 
32'd25540: dataIn1 = 32'd650
; 
32'd25541: dataIn1 = 32'd672
; 
32'd25542: dataIn1 = 32'd700
; 
32'd25543: dataIn1 = 32'd717
; 
32'd25544: dataIn1 = 32'd760
; 
32'd25545: dataIn1 = 32'd769
; 
32'd25546: dataIn1 = 32'd775
; 
32'd25547: dataIn1 = 32'd787
; 
32'd25548: dataIn1 = 32'd592
; 
32'd25549: dataIn1 = 32'd603
; 
32'd25550: dataIn1 = 32'd742
; 
32'd25551: dataIn1 = 32'd745
; 
32'd25552: dataIn1 = 32'd755
; 
32'd25553: dataIn1 = 32'd766
; 
32'd25554: dataIn1 = 32'd767
; 
32'd25555: dataIn1 = 32'd772
; 
32'd25556: dataIn1 = 32'd786
; 
32'd25557: dataIn1 = 32'd573
; 
32'd25558: dataIn1 = 32'd578
; 
32'd25559: dataIn1 = 32'd630
; 
32'd25560: dataIn1 = 32'd634
; 
32'd25561: dataIn1 = 32'd711
; 
32'd25562: dataIn1 = 32'd716
; 
32'd25563: dataIn1 = 32'd726
; 
32'd25564: dataIn1 = 32'd731
; 
32'd25565: dataIn1 = 32'd739
; 
32'd25566: dataIn1 = 32'd771
; 
32'd25567: dataIn1 = 32'd773
; 
32'd25568: dataIn1 = 32'd775
; 
32'd25569: dataIn1 = 32'd793
; 
32'd25570: dataIn1 = 32'd579
; 
32'd25571: dataIn1 = 32'd595
; 
32'd25572: dataIn1 = 32'd627
; 
32'd25573: dataIn1 = 32'd629
; 
32'd25574: dataIn1 = 32'd648
; 
32'd25575: dataIn1 = 32'd670
; 
32'd25576: dataIn1 = 32'd671
; 
32'd25577: dataIn1 = 32'd672
; 
32'd25578: dataIn1 = 32'd684
; 
32'd25579: dataIn1 = 32'd694
; 
32'd25580: dataIn1 = 32'd699
; 
32'd25581: dataIn1 = 32'd710
; 
32'd25582: dataIn1 = 32'd723
; 
32'd25583: dataIn1 = 32'd756
; 
32'd25584: dataIn1 = 32'd796
; 
32'd25585: dataIn1 = 32'd798
; 
32'd25586: dataIn1 = 32'd581
; 
32'd25587: dataIn1 = 32'd590
; 
32'd25588: dataIn1 = 32'd611
; 
32'd25589: dataIn1 = 32'd644
; 
32'd25590: dataIn1 = 32'd645
; 
32'd25591: dataIn1 = 32'd666
; 
32'd25592: dataIn1 = 32'd679
; 
32'd25593: dataIn1 = 32'd682
; 
32'd25594: dataIn1 = 32'd705
; 
32'd25595: dataIn1 = 32'd728
; 
32'd25596: dataIn1 = 32'd748
; 
32'd25597: dataIn1 = 32'd760
; 
32'd25598: dataIn1 = 32'd768
; 
32'd25599: dataIn1 = 32'd772
; 
32'd25600: dataIn1 = 32'd774
; 
32'd25601: dataIn1 = 32'd570
; 
32'd25602: dataIn1 = 32'd577
; 
32'd25603: dataIn1 = 32'd600
; 
32'd25604: dataIn1 = 32'd633
; 
32'd25605: dataIn1 = 32'd637
; 
32'd25606: dataIn1 = 32'd644
; 
32'd25607: dataIn1 = 32'd653
; 
32'd25608: dataIn1 = 32'd671
; 
32'd25609: dataIn1 = 32'd676
; 
32'd25610: dataIn1 = 32'd678
; 
32'd25611: dataIn1 = 32'd697
; 
32'd25612: dataIn1 = 32'd726
; 
32'd25613: dataIn1 = 32'd738
; 
32'd25614: dataIn1 = 32'd784
; 
32'd25615: dataIn1 = 32'd794
; 
32'd25616: dataIn1 = 32'd576
; 
32'd25617: dataIn1 = 32'd577
; 
32'd25618: dataIn1 = 32'd579
; 
32'd25619: dataIn1 = 32'd595
; 
32'd25620: dataIn1 = 32'd597
; 
32'd25621: dataIn1 = 32'd599
; 
32'd25622: dataIn1 = 32'd625
; 
32'd25623: dataIn1 = 32'd644
; 
32'd25624: dataIn1 = 32'd647
; 
32'd25625: dataIn1 = 32'd659
; 
32'd25626: dataIn1 = 32'd660
; 
32'd25627: dataIn1 = 32'd667
; 
32'd25628: dataIn1 = 32'd698
; 
32'd25629: dataIn1 = 32'd702
; 
32'd25630: dataIn1 = 32'd723
; 
32'd25631: dataIn1 = 32'd752
; 
32'd25632: dataIn1 = 32'd763
; 
32'd25633: dataIn1 = 32'd764
; 
32'd25634: dataIn1 = 32'd769
; 
32'd25635: dataIn1 = 32'd772
; 
32'd25636: dataIn1 = 32'd778
; 
32'd25637: dataIn1 = 32'd780
; 
32'd25638: dataIn1 = 32'd784
; 
32'd25639: dataIn1 = 32'd794
; 
32'd25640: dataIn1 = 32'd579
; 
32'd25641: dataIn1 = 32'd587
; 
32'd25642: dataIn1 = 32'd600
; 
32'd25643: dataIn1 = 32'd601
; 
32'd25644: dataIn1 = 32'd644
; 
32'd25645: dataIn1 = 32'd710
; 
32'd25646: dataIn1 = 32'd722
; 
32'd25647: dataIn1 = 32'd753
; 
32'd25648: dataIn1 = 32'd774
; 
32'd25649: dataIn1 = 32'd783
; 
32'd25650: dataIn1 = 32'd796
; 
32'd25651: dataIn1 = 32'd614
; 
32'd25652: dataIn1 = 32'd623
; 
32'd25653: dataIn1 = 32'd684
; 
32'd25654: dataIn1 = 32'd691
; 
32'd25655: dataIn1 = 32'd711
; 
32'd25656: dataIn1 = 32'd727
; 
32'd25657: dataIn1 = 32'd748
; 
32'd25658: dataIn1 = 32'd768
; 
32'd25659: dataIn1 = 32'd769
; 
32'd25660: dataIn1 = 32'd771
; 
32'd25661: dataIn1 = 32'd583
; 
32'd25662: dataIn1 = 32'd614
; 
32'd25663: dataIn1 = 32'd644
; 
32'd25664: dataIn1 = 32'd681
; 
32'd25665: dataIn1 = 32'd709
; 
32'd25666: dataIn1 = 32'd716
; 
32'd25667: dataIn1 = 32'd726
; 
32'd25668: dataIn1 = 32'd748
; 
32'd25669: dataIn1 = 32'd755
; 
32'd25670: dataIn1 = 32'd771
; 
32'd25671: dataIn1 = 32'd774
; 
32'd25672: dataIn1 = 32'd575
; 
32'd25673: dataIn1 = 32'd579
; 
32'd25674: dataIn1 = 32'd586
; 
32'd25675: dataIn1 = 32'd597
; 
32'd25676: dataIn1 = 32'd624
; 
32'd25677: dataIn1 = 32'd637
; 
32'd25678: dataIn1 = 32'd643
; 
32'd25679: dataIn1 = 32'd664
; 
32'd25680: dataIn1 = 32'd674
; 
32'd25681: dataIn1 = 32'd682
; 
32'd25682: dataIn1 = 32'd697
; 
32'd25683: dataIn1 = 32'd701
; 
32'd25684: dataIn1 = 32'd706
; 
32'd25685: dataIn1 = 32'd721
; 
32'd25686: dataIn1 = 32'd726
; 
32'd25687: dataIn1 = 32'd728
; 
32'd25688: dataIn1 = 32'd734
; 
32'd25689: dataIn1 = 32'd744
; 
32'd25690: dataIn1 = 32'd750
; 
32'd25691: dataIn1 = 32'd782
; 
32'd25692: dataIn1 = 32'd798
; 
32'd25693: dataIn1 = 32'd626
; 
32'd25694: dataIn1 = 32'd647
; 
32'd25695: dataIn1 = 32'd649
; 
32'd25696: dataIn1 = 32'd664
; 
32'd25697: dataIn1 = 32'd673
; 
32'd25698: dataIn1 = 32'd698
; 
32'd25699: dataIn1 = 32'd764
; 
32'd25700: dataIn1 = 32'd777
; 
32'd25701: dataIn1 = 32'd784
; 
32'd25702: dataIn1 = 32'd794
; 
32'd25703: dataIn1 = 32'd796
; 
32'd25704: dataIn1 = 32'd797
; 
32'd25705: dataIn1 = 32'd588
; 
32'd25706: dataIn1 = 32'd589
; 
32'd25707: dataIn1 = 32'd596
; 
32'd25708: dataIn1 = 32'd606
; 
32'd25709: dataIn1 = 32'd612
; 
32'd25710: dataIn1 = 32'd647
; 
32'd25711: dataIn1 = 32'd653
; 
32'd25712: dataIn1 = 32'd723
; 
32'd25713: dataIn1 = 32'd746
; 
32'd25714: dataIn1 = 32'd747
; 
32'd25715: dataIn1 = 32'd753
; 
32'd25716: dataIn1 = 32'd757
; 
32'd25717: dataIn1 = 32'd765
; 
32'd25718: dataIn1 = 32'd772
; 
32'd25719: dataIn1 = 32'd780
; 
32'd25720: dataIn1 = 32'd795
; 
32'd25721: dataIn1 = 32'd594
; 
32'd25722: dataIn1 = 32'd611
; 
32'd25723: dataIn1 = 32'd635
; 
32'd25724: dataIn1 = 32'd648
; 
32'd25725: dataIn1 = 32'd657
; 
32'd25726: dataIn1 = 32'd665
; 
32'd25727: dataIn1 = 32'd672
; 
32'd25728: dataIn1 = 32'd684
; 
32'd25729: dataIn1 = 32'd711
; 
32'd25730: dataIn1 = 32'd775
; 
32'd25731: dataIn1 = 32'd778
; 
32'd25732: dataIn1 = 32'd790
; 
32'd25733: dataIn1 = 32'd792
; 
32'd25734: dataIn1 = 32'd594
; 
32'd25735: dataIn1 = 32'd600
; 
32'd25736: dataIn1 = 32'd615
; 
32'd25737: dataIn1 = 32'd648
; 
32'd25738: dataIn1 = 32'd651
; 
32'd25739: dataIn1 = 32'd673
; 
32'd25740: dataIn1 = 32'd706
; 
32'd25741: dataIn1 = 32'd724
; 
32'd25742: dataIn1 = 32'd732
; 
32'd25743: dataIn1 = 32'd757
; 
32'd25744: dataIn1 = 32'd603
; 
32'd25745: dataIn1 = 32'd614
; 
32'd25746: dataIn1 = 32'd615
; 
32'd25747: dataIn1 = 32'd616
; 
32'd25748: dataIn1 = 32'd629
; 
32'd25749: dataIn1 = 32'd633
; 
32'd25750: dataIn1 = 32'd636
; 
32'd25751: dataIn1 = 32'd663
; 
32'd25752: dataIn1 = 32'd703
; 
32'd25753: dataIn1 = 32'd722
; 
32'd25754: dataIn1 = 32'd724
; 
32'd25755: dataIn1 = 32'd727
; 
32'd25756: dataIn1 = 32'd737
; 
32'd25757: dataIn1 = 32'd765
; 
32'd25758: dataIn1 = 32'd775
; 
32'd25759: dataIn1 = 32'd796
; 
32'd25760: dataIn1 = 32'd604
; 
32'd25761: dataIn1 = 32'd647
; 
32'd25762: dataIn1 = 32'd654
; 
32'd25763: dataIn1 = 32'd658
; 
32'd25764: dataIn1 = 32'd668
; 
32'd25765: dataIn1 = 32'd690
; 
32'd25766: dataIn1 = 32'd706
; 
32'd25767: dataIn1 = 32'd739
; 
32'd25768: dataIn1 = 32'd755
; 
32'd25769: dataIn1 = 32'd784
; 
32'd25770: dataIn1 = 32'd785
; 
32'd25771: dataIn1 = 32'd584
; 
32'd25772: dataIn1 = 32'd604
; 
32'd25773: dataIn1 = 32'd620
; 
32'd25774: dataIn1 = 32'd628
; 
32'd25775: dataIn1 = 32'd631
; 
32'd25776: dataIn1 = 32'd636
; 
32'd25777: dataIn1 = 32'd651
; 
32'd25778: dataIn1 = 32'd668
; 
32'd25779: dataIn1 = 32'd673
; 
32'd25780: dataIn1 = 32'd679
; 
32'd25781: dataIn1 = 32'd688
; 
32'd25782: dataIn1 = 32'd711
; 
32'd25783: dataIn1 = 32'd719
; 
32'd25784: dataIn1 = 32'd728
; 
32'd25785: dataIn1 = 32'd736
; 
32'd25786: dataIn1 = 32'd790
; 
32'd25787: dataIn1 = 32'd795
; 
32'd25788: dataIn1 = 32'd586
; 
32'd25789: dataIn1 = 32'd619
; 
32'd25790: dataIn1 = 32'd639
; 
32'd25791: dataIn1 = 32'd650
; 
32'd25792: dataIn1 = 32'd685
; 
32'd25793: dataIn1 = 32'd727
; 
32'd25794: dataIn1 = 32'd739
; 
32'd25795: dataIn1 = 32'd760
; 
32'd25796: dataIn1 = 32'd796
; 
32'd25797: dataIn1 = 32'd612
; 
32'd25798: dataIn1 = 32'd616
; 
32'd25799: dataIn1 = 32'd626
; 
32'd25800: dataIn1 = 32'd634
; 
32'd25801: dataIn1 = 32'd639
; 
32'd25802: dataIn1 = 32'd659
; 
32'd25803: dataIn1 = 32'd672
; 
32'd25804: dataIn1 = 32'd686
; 
32'd25805: dataIn1 = 32'd691
; 
32'd25806: dataIn1 = 32'd716
; 
32'd25807: dataIn1 = 32'd740
; 
32'd25808: dataIn1 = 32'd747
; 
32'd25809: dataIn1 = 32'd758
; 
32'd25810: dataIn1 = 32'd772
; 
32'd25811: dataIn1 = 32'd786
; 
32'd25812: dataIn1 = 32'd791
; 
32'd25813: dataIn1 = 32'd586
; 
32'd25814: dataIn1 = 32'd599
; 
32'd25815: dataIn1 = 32'd619
; 
32'd25816: dataIn1 = 32'd633
; 
32'd25817: dataIn1 = 32'd662
; 
32'd25818: dataIn1 = 32'd672
; 
32'd25819: dataIn1 = 32'd701
; 
32'd25820: dataIn1 = 32'd707
; 
32'd25821: dataIn1 = 32'd711
; 
32'd25822: dataIn1 = 32'd717
; 
32'd25823: dataIn1 = 32'd718
; 
32'd25824: dataIn1 = 32'd720
; 
32'd25825: dataIn1 = 32'd722
; 
32'd25826: dataIn1 = 32'd730
; 
32'd25827: dataIn1 = 32'd762
; 
32'd25828: dataIn1 = 32'd773
; 
32'd25829: dataIn1 = 32'd775
; 
32'd25830: dataIn1 = 32'd779
; 
32'd25831: dataIn1 = 32'd790
; 
32'd25832: dataIn1 = 32'd588
; 
32'd25833: dataIn1 = 32'd592
; 
32'd25834: dataIn1 = 32'd615
; 
32'd25835: dataIn1 = 32'd629
; 
32'd25836: dataIn1 = 32'd641
; 
32'd25837: dataIn1 = 32'd643
; 
32'd25838: dataIn1 = 32'd647
; 
32'd25839: dataIn1 = 32'd654
; 
32'd25840: dataIn1 = 32'd658
; 
32'd25841: dataIn1 = 32'd702
; 
32'd25842: dataIn1 = 32'd755
; 
32'd25843: dataIn1 = 32'd759
; 
32'd25844: dataIn1 = 32'd772
; 
32'd25845: dataIn1 = 32'd778
; 
32'd25846: dataIn1 = 32'd784
; 
32'd25847: dataIn1 = 32'd786
; 
32'd25848: dataIn1 = 32'd789
; 
32'd25849: dataIn1 = 32'd798
; 
32'd25850: dataIn1 = 32'd598
; 
32'd25851: dataIn1 = 32'd612
; 
32'd25852: dataIn1 = 32'd624
; 
32'd25853: dataIn1 = 32'd645
; 
32'd25854: dataIn1 = 32'd651
; 
32'd25855: dataIn1 = 32'd655
; 
32'd25856: dataIn1 = 32'd673
; 
32'd25857: dataIn1 = 32'd675
; 
32'd25858: dataIn1 = 32'd685
; 
32'd25859: dataIn1 = 32'd707
; 
32'd25860: dataIn1 = 32'd712
; 
32'd25861: dataIn1 = 32'd715
; 
32'd25862: dataIn1 = 32'd734
; 
32'd25863: dataIn1 = 32'd735
; 
32'd25864: dataIn1 = 32'd741
; 
32'd25865: dataIn1 = 32'd761
; 
32'd25866: dataIn1 = 32'd777
; 
32'd25867: dataIn1 = 32'd781
; 
32'd25868: dataIn1 = 32'd594
; 
32'd25869: dataIn1 = 32'd609
; 
32'd25870: dataIn1 = 32'd621
; 
32'd25871: dataIn1 = 32'd629
; 
32'd25872: dataIn1 = 32'd630
; 
32'd25873: dataIn1 = 32'd637
; 
32'd25874: dataIn1 = 32'd684
; 
32'd25875: dataIn1 = 32'd695
; 
32'd25876: dataIn1 = 32'd720
; 
32'd25877: dataIn1 = 32'd721
; 
32'd25878: dataIn1 = 32'd589
; 
32'd25879: dataIn1 = 32'd601
; 
32'd25880: dataIn1 = 32'd625
; 
32'd25881: dataIn1 = 32'd705
; 
32'd25882: dataIn1 = 32'd717
; 
32'd25883: dataIn1 = 32'd753
; 
32'd25884: dataIn1 = 32'd760
; 
32'd25885: dataIn1 = 32'd773
; 
32'd25886: dataIn1 = 32'd775
; 
32'd25887: dataIn1 = 32'd792
; 
32'd25888: dataIn1 = 32'd679
; 
32'd25889: dataIn1 = 32'd688
; 
32'd25890: dataIn1 = 32'd692
; 
32'd25891: dataIn1 = 32'd709
; 
32'd25892: dataIn1 = 32'd715
; 
32'd25893: dataIn1 = 32'd719
; 
32'd25894: dataIn1 = 32'd760
; 
32'd25895: dataIn1 = 32'd765
; 
32'd25896: dataIn1 = 32'd772
; 
32'd25897: dataIn1 = 32'd796
; 
32'd25898: dataIn1 = 32'd618
; 
32'd25899: dataIn1 = 32'd621
; 
32'd25900: dataIn1 = 32'd679
; 
32'd25901: dataIn1 = 32'd690
; 
32'd25902: dataIn1 = 32'd704
; 
32'd25903: dataIn1 = 32'd744
; 
32'd25904: dataIn1 = 32'd753
; 
32'd25905: dataIn1 = 32'd756
; 
32'd25906: dataIn1 = 32'd780
; 
32'd25907: dataIn1 = 32'd788
; 
32'd25908: dataIn1 = 32'd600
; 
32'd25909: dataIn1 = 32'd611
; 
32'd25910: dataIn1 = 32'd677
; 
32'd25911: dataIn1 = 32'd688
; 
32'd25912: dataIn1 = 32'd697
; 
32'd25913: dataIn1 = 32'd706
; 
32'd25914: dataIn1 = 32'd708
; 
32'd25915: dataIn1 = 32'd713
; 
32'd25916: dataIn1 = 32'd737
; 
32'd25917: dataIn1 = 32'd760
; 
32'd25918: dataIn1 = 32'd772
; 
32'd25919: dataIn1 = 32'd794
; 
32'd25920: dataIn1 = 32'd596
; 
32'd25921: dataIn1 = 32'd614
; 
32'd25922: dataIn1 = 32'd635
; 
32'd25923: dataIn1 = 32'd650
; 
32'd25924: dataIn1 = 32'd651
; 
32'd25925: dataIn1 = 32'd652
; 
32'd25926: dataIn1 = 32'd685
; 
32'd25927: dataIn1 = 32'd686
; 
32'd25928: dataIn1 = 32'd697
; 
32'd25929: dataIn1 = 32'd713
; 
32'd25930: dataIn1 = 32'd717
; 
32'd25931: dataIn1 = 32'd721
; 
32'd25932: dataIn1 = 32'd722
; 
32'd25933: dataIn1 = 32'd741
; 
32'd25934: dataIn1 = 32'd760
; 
32'd25935: dataIn1 = 32'd781
; 
32'd25936: dataIn1 = 32'd783
; 
32'd25937: dataIn1 = 32'd626
; 
32'd25938: dataIn1 = 32'd629
; 
32'd25939: dataIn1 = 32'd649
; 
32'd25940: dataIn1 = 32'd692
; 
32'd25941: dataIn1 = 32'd734
; 
32'd25942: dataIn1 = 32'd758
; 
32'd25943: dataIn1 = 32'd765
; 
32'd25944: dataIn1 = 32'd604
; 
32'd25945: dataIn1 = 32'd607
; 
32'd25946: dataIn1 = 32'd610
; 
32'd25947: dataIn1 = 32'd616
; 
32'd25948: dataIn1 = 32'd644
; 
32'd25949: dataIn1 = 32'd651
; 
32'd25950: dataIn1 = 32'd658
; 
32'd25951: dataIn1 = 32'd718
; 
32'd25952: dataIn1 = 32'd719
; 
32'd25953: dataIn1 = 32'd725
; 
32'd25954: dataIn1 = 32'd739
; 
32'd25955: dataIn1 = 32'd748
; 
32'd25956: dataIn1 = 32'd754
; 
32'd25957: dataIn1 = 32'd763
; 
32'd25958: dataIn1 = 32'd771
; 
32'd25959: dataIn1 = 32'd778
; 
32'd25960: dataIn1 = 32'd779
; 
32'd25961: dataIn1 = 32'd785
; 
32'd25962: dataIn1 = 32'd619
; 
32'd25963: dataIn1 = 32'd622
; 
32'd25964: dataIn1 = 32'd631
; 
32'd25965: dataIn1 = 32'd636
; 
32'd25966: dataIn1 = 32'd644
; 
32'd25967: dataIn1 = 32'd700
; 
32'd25968: dataIn1 = 32'd738
; 
32'd25969: dataIn1 = 32'd739
; 
32'd25970: dataIn1 = 32'd763
; 
32'd25971: dataIn1 = 32'd769
; 
32'd25972: dataIn1 = 32'd774
; 
32'd25973: dataIn1 = 32'd787
; 
32'd25974: dataIn1 = 32'd790
; 
32'd25975: dataIn1 = 32'd629
; 
32'd25976: dataIn1 = 32'd631
; 
32'd25977: dataIn1 = 32'd647
; 
32'd25978: dataIn1 = 32'd657
; 
32'd25979: dataIn1 = 32'd662
; 
32'd25980: dataIn1 = 32'd669
; 
32'd25981: dataIn1 = 32'd683
; 
32'd25982: dataIn1 = 32'd685
; 
32'd25983: dataIn1 = 32'd690
; 
32'd25984: dataIn1 = 32'd722
; 
32'd25985: dataIn1 = 32'd746
; 
32'd25986: dataIn1 = 32'd788
; 
32'd25987: dataIn1 = 32'd792
; 
32'd25988: dataIn1 = 32'd795
; 
32'd25989: dataIn1 = 32'd600
; 
32'd25990: dataIn1 = 32'd604
; 
32'd25991: dataIn1 = 32'd626
; 
32'd25992: dataIn1 = 32'd633
; 
32'd25993: dataIn1 = 32'd651
; 
32'd25994: dataIn1 = 32'd658
; 
32'd25995: dataIn1 = 32'd666
; 
32'd25996: dataIn1 = 32'd680
; 
32'd25997: dataIn1 = 32'd704
; 
32'd25998: dataIn1 = 32'd706
; 
32'd25999: dataIn1 = 32'd708
; 
32'd26000: dataIn1 = 32'd712
; 
32'd26001: dataIn1 = 32'd738
; 
32'd26002: dataIn1 = 32'd740
; 
32'd26003: dataIn1 = 32'd773
; 
32'd26004: dataIn1 = 32'd607
; 
32'd26005: dataIn1 = 32'd616
; 
32'd26006: dataIn1 = 32'd623
; 
32'd26007: dataIn1 = 32'd682
; 
32'd26008: dataIn1 = 32'd696
; 
32'd26009: dataIn1 = 32'd702
; 
32'd26010: dataIn1 = 32'd709
; 
32'd26011: dataIn1 = 32'd714
; 
32'd26012: dataIn1 = 32'd769
; 
32'd26013: dataIn1 = 32'd779
; 
32'd26014: dataIn1 = 32'd784
; 
32'd26015: dataIn1 = 32'd791
; 
32'd26016: dataIn1 = 32'd800
; 
32'd26017: dataIn1 = 32'd635
; 
32'd26018: dataIn1 = 32'd662
; 
32'd26019: dataIn1 = 32'd664
; 
32'd26020: dataIn1 = 32'd685
; 
32'd26021: dataIn1 = 32'd694
; 
32'd26022: dataIn1 = 32'd695
; 
32'd26023: dataIn1 = 32'd712
; 
32'd26024: dataIn1 = 32'd751
; 
32'd26025: dataIn1 = 32'd756
; 
32'd26026: dataIn1 = 32'd759
; 
32'd26027: dataIn1 = 32'd602
; 
32'd26028: dataIn1 = 32'd604
; 
32'd26029: dataIn1 = 32'd615
; 
32'd26030: dataIn1 = 32'd619
; 
32'd26031: dataIn1 = 32'd645
; 
32'd26032: dataIn1 = 32'd656
; 
32'd26033: dataIn1 = 32'd685
; 
32'd26034: dataIn1 = 32'd688
; 
32'd26035: dataIn1 = 32'd720
; 
32'd26036: dataIn1 = 32'd741
; 
32'd26037: dataIn1 = 32'd746
; 
32'd26038: dataIn1 = 32'd747
; 
32'd26039: dataIn1 = 32'd614
; 
32'd26040: dataIn1 = 32'd618
; 
32'd26041: dataIn1 = 32'd625
; 
32'd26042: dataIn1 = 32'd654
; 
32'd26043: dataIn1 = 32'd665
; 
32'd26044: dataIn1 = 32'd676
; 
32'd26045: dataIn1 = 32'd681
; 
32'd26046: dataIn1 = 32'd702
; 
32'd26047: dataIn1 = 32'd706
; 
32'd26048: dataIn1 = 32'd727
; 
32'd26049: dataIn1 = 32'd743
; 
32'd26050: dataIn1 = 32'd757
; 
32'd26051: dataIn1 = 32'd766
; 
32'd26052: dataIn1 = 32'd771
; 
32'd26053: dataIn1 = 32'd777
; 
32'd26054: dataIn1 = 32'd621
; 
32'd26055: dataIn1 = 32'd642
; 
32'd26056: dataIn1 = 32'd654
; 
32'd26057: dataIn1 = 32'd676
; 
32'd26058: dataIn1 = 32'd678
; 
32'd26059: dataIn1 = 32'd695
; 
32'd26060: dataIn1 = 32'd764
; 
32'd26061: dataIn1 = 32'd798
; 
32'd26062: dataIn1 = 32'd609
; 
32'd26063: dataIn1 = 32'd618
; 
32'd26064: dataIn1 = 32'd634
; 
32'd26065: dataIn1 = 32'd678
; 
32'd26066: dataIn1 = 32'd744
; 
32'd26067: dataIn1 = 32'd757
; 
32'd26068: dataIn1 = 32'd758
; 
32'd26069: dataIn1 = 32'd777
; 
32'd26070: dataIn1 = 32'd791
; 
32'd26071: dataIn1 = 32'd797
; 
32'd26072: dataIn1 = 32'd641
; 
32'd26073: dataIn1 = 32'd642
; 
32'd26074: dataIn1 = 32'd649
; 
32'd26075: dataIn1 = 32'd657
; 
32'd26076: dataIn1 = 32'd666
; 
32'd26077: dataIn1 = 32'd671
; 
32'd26078: dataIn1 = 32'd688
; 
32'd26079: dataIn1 = 32'd696
; 
32'd26080: dataIn1 = 32'd706
; 
32'd26081: dataIn1 = 32'd752
; 
32'd26082: dataIn1 = 32'd761
; 
32'd26083: dataIn1 = 32'd763
; 
32'd26084: dataIn1 = 32'd780
; 
32'd26085: dataIn1 = 32'd783
; 
32'd26086: dataIn1 = 32'd790
; 
32'd26087: dataIn1 = 32'd609
; 
32'd26088: dataIn1 = 32'd632
; 
32'd26089: dataIn1 = 32'd666
; 
32'd26090: dataIn1 = 32'd671
; 
32'd26091: dataIn1 = 32'd696
; 
32'd26092: dataIn1 = 32'd710
; 
32'd26093: dataIn1 = 32'd721
; 
32'd26094: dataIn1 = 32'd731
; 
32'd26095: dataIn1 = 32'd750
; 
32'd26096: dataIn1 = 32'd764
; 
32'd26097: dataIn1 = 32'd777
; 
32'd26098: dataIn1 = 32'd785
; 
32'd26099: dataIn1 = 32'd798
; 
32'd26100: dataIn1 = 32'd800
; 
32'd26101: dataIn1 = 32'd621
; 
32'd26102: dataIn1 = 32'd623
; 
32'd26103: dataIn1 = 32'd654
; 
32'd26104: dataIn1 = 32'd705
; 
32'd26105: dataIn1 = 32'd714
; 
32'd26106: dataIn1 = 32'd723
; 
32'd26107: dataIn1 = 32'd743
; 
32'd26108: dataIn1 = 32'd749
; 
32'd26109: dataIn1 = 32'd617
; 
32'd26110: dataIn1 = 32'd630
; 
32'd26111: dataIn1 = 32'd652
; 
32'd26112: dataIn1 = 32'd654
; 
32'd26113: dataIn1 = 32'd672
; 
32'd26114: dataIn1 = 32'd673
; 
32'd26115: dataIn1 = 32'd692
; 
32'd26116: dataIn1 = 32'd729
; 
32'd26117: dataIn1 = 32'd731
; 
32'd26118: dataIn1 = 32'd742
; 
32'd26119: dataIn1 = 32'd766
; 
32'd26120: dataIn1 = 32'd610
; 
32'd26121: dataIn1 = 32'd616
; 
32'd26122: dataIn1 = 32'd660
; 
32'd26123: dataIn1 = 32'd680
; 
32'd26124: dataIn1 = 32'd713
; 
32'd26125: dataIn1 = 32'd751
; 
32'd26126: dataIn1 = 32'd761
; 
32'd26127: dataIn1 = 32'd780
; 
32'd26128: dataIn1 = 32'd620
; 
32'd26129: dataIn1 = 32'd624
; 
32'd26130: dataIn1 = 32'd697
; 
32'd26131: dataIn1 = 32'd699
; 
32'd26132: dataIn1 = 32'd719
; 
32'd26133: dataIn1 = 32'd721
; 
32'd26134: dataIn1 = 32'd750
; 
32'd26135: dataIn1 = 32'd759
; 
32'd26136: dataIn1 = 32'd764
; 
32'd26137: dataIn1 = 32'd767
; 
32'd26138: dataIn1 = 32'd611
; 
32'd26139: dataIn1 = 32'd627
; 
32'd26140: dataIn1 = 32'd659
; 
32'd26141: dataIn1 = 32'd666
; 
32'd26142: dataIn1 = 32'd723
; 
32'd26143: dataIn1 = 32'd730
; 
32'd26144: dataIn1 = 32'd745
; 
32'd26145: dataIn1 = 32'd752
; 
32'd26146: dataIn1 = 32'd768
; 
32'd26147: dataIn1 = 32'd633
; 
32'd26148: dataIn1 = 32'd637
; 
32'd26149: dataIn1 = 32'd672
; 
32'd26150: dataIn1 = 32'd695
; 
32'd26151: dataIn1 = 32'd726
; 
32'd26152: dataIn1 = 32'd742
; 
32'd26153: dataIn1 = 32'd748
; 
32'd26154: dataIn1 = 32'd755
; 
32'd26155: dataIn1 = 32'd782
; 
32'd26156: dataIn1 = 32'd613
; 
32'd26157: dataIn1 = 32'd659
; 
32'd26158: dataIn1 = 32'd662
; 
32'd26159: dataIn1 = 32'd686
; 
32'd26160: dataIn1 = 32'd689
; 
32'd26161: dataIn1 = 32'd691
; 
32'd26162: dataIn1 = 32'd694
; 
32'd26163: dataIn1 = 32'd711
; 
32'd26164: dataIn1 = 32'd726
; 
32'd26165: dataIn1 = 32'd730
; 
32'd26166: dataIn1 = 32'd757
; 
32'd26167: dataIn1 = 32'd774
; 
32'd26168: dataIn1 = 32'd786
; 
32'd26169: dataIn1 = 32'd639
; 
32'd26170: dataIn1 = 32'd644
; 
32'd26171: dataIn1 = 32'd684
; 
32'd26172: dataIn1 = 32'd690
; 
32'd26173: dataIn1 = 32'd692
; 
32'd26174: dataIn1 = 32'd702
; 
32'd26175: dataIn1 = 32'd730
; 
32'd26176: dataIn1 = 32'd749
; 
32'd26177: dataIn1 = 32'd752
; 
32'd26178: dataIn1 = 32'd756
; 
32'd26179: dataIn1 = 32'd762
; 
32'd26180: dataIn1 = 32'd766
; 
32'd26181: dataIn1 = 32'd777
; 
32'd26182: dataIn1 = 32'd789
; 
32'd26183: dataIn1 = 32'd796
; 
32'd26184: dataIn1 = 32'd652
; 
32'd26185: dataIn1 = 32'd661
; 
32'd26186: dataIn1 = 32'd664
; 
32'd26187: dataIn1 = 32'd685
; 
32'd26188: dataIn1 = 32'd700
; 
32'd26189: dataIn1 = 32'd728
; 
32'd26190: dataIn1 = 32'd747
; 
32'd26191: dataIn1 = 32'd788
; 
32'd26192: dataIn1 = 32'd643
; 
32'd26193: dataIn1 = 32'd646
; 
32'd26194: dataIn1 = 32'd651
; 
32'd26195: dataIn1 = 32'd656
; 
32'd26196: dataIn1 = 32'd673
; 
32'd26197: dataIn1 = 32'd694
; 
32'd26198: dataIn1 = 32'd707
; 
32'd26199: dataIn1 = 32'd709
; 
32'd26200: dataIn1 = 32'd712
; 
32'd26201: dataIn1 = 32'd714
; 
32'd26202: dataIn1 = 32'd719
; 
32'd26203: dataIn1 = 32'd729
; 
32'd26204: dataIn1 = 32'd740
; 
32'd26205: dataIn1 = 32'd763
; 
32'd26206: dataIn1 = 32'd625
; 
32'd26207: dataIn1 = 32'd677
; 
32'd26208: dataIn1 = 32'd678
; 
32'd26209: dataIn1 = 32'd684
; 
32'd26210: dataIn1 = 32'd690
; 
32'd26211: dataIn1 = 32'd691
; 
32'd26212: dataIn1 = 32'd706
; 
32'd26213: dataIn1 = 32'd722
; 
32'd26214: dataIn1 = 32'd747
; 
32'd26215: dataIn1 = 32'd749
; 
32'd26216: dataIn1 = 32'd786
; 
32'd26217: dataIn1 = 32'd619
; 
32'd26218: dataIn1 = 32'd632
; 
32'd26219: dataIn1 = 32'd655
; 
32'd26220: dataIn1 = 32'd682
; 
32'd26221: dataIn1 = 32'd698
; 
32'd26222: dataIn1 = 32'd706
; 
32'd26223: dataIn1 = 32'd707
; 
32'd26224: dataIn1 = 32'd753
; 
32'd26225: dataIn1 = 32'd774
; 
32'd26226: dataIn1 = 32'd799
; 
32'd26227: dataIn1 = 32'd629
; 
32'd26228: dataIn1 = 32'd639
; 
32'd26229: dataIn1 = 32'd674
; 
32'd26230: dataIn1 = 32'd679
; 
32'd26231: dataIn1 = 32'd742
; 
32'd26232: dataIn1 = 32'd757
; 
32'd26233: dataIn1 = 32'd764
; 
32'd26234: dataIn1 = 32'd770
; 
32'd26235: dataIn1 = 32'd783
; 
32'd26236: dataIn1 = 32'd637
; 
32'd26237: dataIn1 = 32'd640
; 
32'd26238: dataIn1 = 32'd652
; 
32'd26239: dataIn1 = 32'd682
; 
32'd26240: dataIn1 = 32'd683
; 
32'd26241: dataIn1 = 32'd687
; 
32'd26242: dataIn1 = 32'd690
; 
32'd26243: dataIn1 = 32'd695
; 
32'd26244: dataIn1 = 32'd697
; 
32'd26245: dataIn1 = 32'd728
; 
32'd26246: dataIn1 = 32'd747
; 
32'd26247: dataIn1 = 32'd793
; 
32'd26248: dataIn1 = 32'd794
; 
32'd26249: dataIn1 = 32'd628
; 
32'd26250: dataIn1 = 32'd657
; 
32'd26251: dataIn1 = 32'd681
; 
32'd26252: dataIn1 = 32'd685
; 
32'd26253: dataIn1 = 32'd687
; 
32'd26254: dataIn1 = 32'd695
; 
32'd26255: dataIn1 = 32'd700
; 
32'd26256: dataIn1 = 32'd702
; 
32'd26257: dataIn1 = 32'd718
; 
32'd26258: dataIn1 = 32'd726
; 
32'd26259: dataIn1 = 32'd734
; 
32'd26260: dataIn1 = 32'd756
; 
32'd26261: dataIn1 = 32'd763
; 
32'd26262: dataIn1 = 32'd782
; 
32'd26263: dataIn1 = 32'd785
; 
32'd26264: dataIn1 = 32'd622
; 
32'd26265: dataIn1 = 32'd641
; 
32'd26266: dataIn1 = 32'd642
; 
32'd26267: dataIn1 = 32'd649
; 
32'd26268: dataIn1 = 32'd681
; 
32'd26269: dataIn1 = 32'd684
; 
32'd26270: dataIn1 = 32'd691
; 
32'd26271: dataIn1 = 32'd697
; 
32'd26272: dataIn1 = 32'd708
; 
32'd26273: dataIn1 = 32'd712
; 
32'd26274: dataIn1 = 32'd746
; 
32'd26275: dataIn1 = 32'd771
; 
32'd26276: dataIn1 = 32'd642
; 
32'd26277: dataIn1 = 32'd652
; 
32'd26278: dataIn1 = 32'd668
; 
32'd26279: dataIn1 = 32'd687
; 
32'd26280: dataIn1 = 32'd725
; 
32'd26281: dataIn1 = 32'd728
; 
32'd26282: dataIn1 = 32'd744
; 
32'd26283: dataIn1 = 32'd797
; 
32'd26284: dataIn1 = 32'd799
; 
32'd26285: dataIn1 = 32'd658
; 
32'd26286: dataIn1 = 32'd668
; 
32'd26287: dataIn1 = 32'd682
; 
32'd26288: dataIn1 = 32'd695
; 
32'd26289: dataIn1 = 32'd718
; 
32'd26290: dataIn1 = 32'd730
; 
32'd26291: dataIn1 = 32'd756
; 
32'd26292: dataIn1 = 32'd797
; 
32'd26293: dataIn1 = 32'd636
; 
32'd26294: dataIn1 = 32'd658
; 
32'd26295: dataIn1 = 32'd665
; 
32'd26296: dataIn1 = 32'd667
; 
32'd26297: dataIn1 = 32'd672
; 
32'd26298: dataIn1 = 32'd697
; 
32'd26299: dataIn1 = 32'd701
; 
32'd26300: dataIn1 = 32'd702
; 
32'd26301: dataIn1 = 32'd718
; 
32'd26302: dataIn1 = 32'd721
; 
32'd26303: dataIn1 = 32'd732
; 
32'd26304: dataIn1 = 32'd735
; 
32'd26305: dataIn1 = 32'd744
; 
32'd26306: dataIn1 = 32'd746
; 
32'd26307: dataIn1 = 32'd778
; 
32'd26308: dataIn1 = 32'd792
; 
32'd26309: dataIn1 = 32'd630
; 
32'd26310: dataIn1 = 32'd637
; 
32'd26311: dataIn1 = 32'd694
; 
32'd26312: dataIn1 = 32'd695
; 
32'd26313: dataIn1 = 32'd699
; 
32'd26314: dataIn1 = 32'd701
; 
32'd26315: dataIn1 = 32'd705
; 
32'd26316: dataIn1 = 32'd722
; 
32'd26317: dataIn1 = 32'd745
; 
32'd26318: dataIn1 = 32'd749
; 
32'd26319: dataIn1 = 32'd755
; 
32'd26320: dataIn1 = 32'd776
; 
32'd26321: dataIn1 = 32'd779
; 
32'd26322: dataIn1 = 32'd787
; 
32'd26323: dataIn1 = 32'd791
; 
32'd26324: dataIn1 = 32'd792
; 
32'd26325: dataIn1 = 32'd793
; 
32'd26326: dataIn1 = 32'd651
; 
32'd26327: dataIn1 = 32'd665
; 
32'd26328: dataIn1 = 32'd680
; 
32'd26329: dataIn1 = 32'd695
; 
32'd26330: dataIn1 = 32'd746
; 
32'd26331: dataIn1 = 32'd759
; 
32'd26332: dataIn1 = 32'd774
; 
32'd26333: dataIn1 = 32'd795
; 
32'd26334: dataIn1 = 32'd796
; 
32'd26335: dataIn1 = 32'd641
; 
32'd26336: dataIn1 = 32'd645
; 
32'd26337: dataIn1 = 32'd667
; 
32'd26338: dataIn1 = 32'd677
; 
32'd26339: dataIn1 = 32'd690
; 
32'd26340: dataIn1 = 32'd701
; 
32'd26341: dataIn1 = 32'd736
; 
32'd26342: dataIn1 = 32'd752
; 
32'd26343: dataIn1 = 32'd757
; 
32'd26344: dataIn1 = 32'd771
; 
32'd26345: dataIn1 = 32'd790
; 
32'd26346: dataIn1 = 32'd795
; 
32'd26347: dataIn1 = 32'd629
; 
32'd26348: dataIn1 = 32'd635
; 
32'd26349: dataIn1 = 32'd638
; 
32'd26350: dataIn1 = 32'd656
; 
32'd26351: dataIn1 = 32'd658
; 
32'd26352: dataIn1 = 32'd703
; 
32'd26353: dataIn1 = 32'd704
; 
32'd26354: dataIn1 = 32'd709
; 
32'd26355: dataIn1 = 32'd762
; 
32'd26356: dataIn1 = 32'd640
; 
32'd26357: dataIn1 = 32'd654
; 
32'd26358: dataIn1 = 32'd660
; 
32'd26359: dataIn1 = 32'd721
; 
32'd26360: dataIn1 = 32'd775
; 
32'd26361: dataIn1 = 32'd643
; 
32'd26362: dataIn1 = 32'd670
; 
32'd26363: dataIn1 = 32'd680
; 
32'd26364: dataIn1 = 32'd690
; 
32'd26365: dataIn1 = 32'd694
; 
32'd26366: dataIn1 = 32'd710
; 
32'd26367: dataIn1 = 32'd754
; 
32'd26368: dataIn1 = 32'd770
; 
32'd26369: dataIn1 = 32'd780
; 
32'd26370: dataIn1 = 32'd794
; 
32'd26371: dataIn1 = 32'd796
; 
32'd26372: dataIn1 = 32'd797
; 
32'd26373: dataIn1 = 32'd638
; 
32'd26374: dataIn1 = 32'd667
; 
32'd26375: dataIn1 = 32'd668
; 
32'd26376: dataIn1 = 32'd675
; 
32'd26377: dataIn1 = 32'd758
; 
32'd26378: dataIn1 = 32'd760
; 
32'd26379: dataIn1 = 32'd634
; 
32'd26380: dataIn1 = 32'd645
; 
32'd26381: dataIn1 = 32'd663
; 
32'd26382: dataIn1 = 32'd684
; 
32'd26383: dataIn1 = 32'd685
; 
32'd26384: dataIn1 = 32'd712
; 
32'd26385: dataIn1 = 32'd743
; 
32'd26386: dataIn1 = 32'd750
; 
32'd26387: dataIn1 = 32'd752
; 
32'd26388: dataIn1 = 32'd767
; 
32'd26389: dataIn1 = 32'd773
; 
32'd26390: dataIn1 = 32'd796
; 
32'd26391: dataIn1 = 32'd638
; 
32'd26392: dataIn1 = 32'd644
; 
32'd26393: dataIn1 = 32'd646
; 
32'd26394: dataIn1 = 32'd666
; 
32'd26395: dataIn1 = 32'd668
; 
32'd26396: dataIn1 = 32'd677
; 
32'd26397: dataIn1 = 32'd689
; 
32'd26398: dataIn1 = 32'd716
; 
32'd26399: dataIn1 = 32'd732
; 
32'd26400: dataIn1 = 32'd736
; 
32'd26401: dataIn1 = 32'd753
; 
32'd26402: dataIn1 = 32'd775
; 
32'd26403: dataIn1 = 32'd782
; 
32'd26404: dataIn1 = 32'd788
; 
32'd26405: dataIn1 = 32'd789
; 
32'd26406: dataIn1 = 32'd791
; 
32'd26407: dataIn1 = 32'd661
; 
32'd26408: dataIn1 = 32'd667
; 
32'd26409: dataIn1 = 32'd676
; 
32'd26410: dataIn1 = 32'd725
; 
32'd26411: dataIn1 = 32'd730
; 
32'd26412: dataIn1 = 32'd735
; 
32'd26413: dataIn1 = 32'd757
; 
32'd26414: dataIn1 = 32'd767
; 
32'd26415: dataIn1 = 32'd639
; 
32'd26416: dataIn1 = 32'd643
; 
32'd26417: dataIn1 = 32'd644
; 
32'd26418: dataIn1 = 32'd669
; 
32'd26419: dataIn1 = 32'd692
; 
32'd26420: dataIn1 = 32'd729
; 
32'd26421: dataIn1 = 32'd734
; 
32'd26422: dataIn1 = 32'd756
; 
32'd26423: dataIn1 = 32'd791
; 
32'd26424: dataIn1 = 32'd642
; 
32'd26425: dataIn1 = 32'd644
; 
32'd26426: dataIn1 = 32'd662
; 
32'd26427: dataIn1 = 32'd702
; 
32'd26428: dataIn1 = 32'd747
; 
32'd26429: dataIn1 = 32'd642
; 
32'd26430: dataIn1 = 32'd652
; 
32'd26431: dataIn1 = 32'd659
; 
32'd26432: dataIn1 = 32'd660
; 
32'd26433: dataIn1 = 32'd665
; 
32'd26434: dataIn1 = 32'd686
; 
32'd26435: dataIn1 = 32'd692
; 
32'd26436: dataIn1 = 32'd709
; 
32'd26437: dataIn1 = 32'd717
; 
32'd26438: dataIn1 = 32'd722
; 
32'd26439: dataIn1 = 32'd723
; 
32'd26440: dataIn1 = 32'd736
; 
32'd26441: dataIn1 = 32'd764
; 
32'd26442: dataIn1 = 32'd788
; 
32'd26443: dataIn1 = 32'd793
; 
32'd26444: dataIn1 = 32'd794
; 
32'd26445: dataIn1 = 32'd799
; 
32'd26446: dataIn1 = 32'd644
; 
32'd26447: dataIn1 = 32'd658
; 
32'd26448: dataIn1 = 32'd683
; 
32'd26449: dataIn1 = 32'd689
; 
32'd26450: dataIn1 = 32'd732
; 
32'd26451: dataIn1 = 32'd738
; 
32'd26452: dataIn1 = 32'd756
; 
32'd26453: dataIn1 = 32'd780
; 
32'd26454: dataIn1 = 32'd641
; 
32'd26455: dataIn1 = 32'd671
; 
32'd26456: dataIn1 = 32'd686
; 
32'd26457: dataIn1 = 32'd701
; 
32'd26458: dataIn1 = 32'd712
; 
32'd26459: dataIn1 = 32'd736
; 
32'd26460: dataIn1 = 32'd748
; 
32'd26461: dataIn1 = 32'd766
; 
32'd26462: dataIn1 = 32'd776
; 
32'd26463: dataIn1 = 32'd795
; 
32'd26464: dataIn1 = 32'd798
; 
32'd26465: dataIn1 = 32'd655
; 
32'd26466: dataIn1 = 32'd669
; 
32'd26467: dataIn1 = 32'd673
; 
32'd26468: dataIn1 = 32'd680
; 
32'd26469: dataIn1 = 32'd681
; 
32'd26470: dataIn1 = 32'd689
; 
32'd26471: dataIn1 = 32'd695
; 
32'd26472: dataIn1 = 32'd700
; 
32'd26473: dataIn1 = 32'd713
; 
32'd26474: dataIn1 = 32'd715
; 
32'd26475: dataIn1 = 32'd742
; 
32'd26476: dataIn1 = 32'd743
; 
32'd26477: dataIn1 = 32'd800
; 
32'd26478: dataIn1 = 32'd649
; 
32'd26479: dataIn1 = 32'd657
; 
32'd26480: dataIn1 = 32'd720
; 
32'd26481: dataIn1 = 32'd723
; 
32'd26482: dataIn1 = 32'd776
; 
32'd26483: dataIn1 = 32'd668
; 
32'd26484: dataIn1 = 32'd670
; 
32'd26485: dataIn1 = 32'd723
; 
32'd26486: dataIn1 = 32'd743
; 
32'd26487: dataIn1 = 32'd759
; 
32'd26488: dataIn1 = 32'd762
; 
32'd26489: dataIn1 = 32'd768
; 
32'd26490: dataIn1 = 32'd798
; 
32'd26491: dataIn1 = 32'd656
; 
32'd26492: dataIn1 = 32'd672
; 
32'd26493: dataIn1 = 32'd678
; 
32'd26494: dataIn1 = 32'd681
; 
32'd26495: dataIn1 = 32'd708
; 
32'd26496: dataIn1 = 32'd715
; 
32'd26497: dataIn1 = 32'd726
; 
32'd26498: dataIn1 = 32'd744
; 
32'd26499: dataIn1 = 32'd777
; 
32'd26500: dataIn1 = 32'd778
; 
32'd26501: dataIn1 = 32'd656
; 
32'd26502: dataIn1 = 32'd658
; 
32'd26503: dataIn1 = 32'd667
; 
32'd26504: dataIn1 = 32'd672
; 
32'd26505: dataIn1 = 32'd675
; 
32'd26506: dataIn1 = 32'd685
; 
32'd26507: dataIn1 = 32'd694
; 
32'd26508: dataIn1 = 32'd697
; 
32'd26509: dataIn1 = 32'd712
; 
32'd26510: dataIn1 = 32'd735
; 
32'd26511: dataIn1 = 32'd759
; 
32'd26512: dataIn1 = 32'd799
; 
32'd26513: dataIn1 = 32'd670
; 
32'd26514: dataIn1 = 32'd672
; 
32'd26515: dataIn1 = 32'd711
; 
32'd26516: dataIn1 = 32'd743
; 
32'd26517: dataIn1 = 32'd749
; 
32'd26518: dataIn1 = 32'd752
; 
32'd26519: dataIn1 = 32'd669
; 
32'd26520: dataIn1 = 32'd683
; 
32'd26521: dataIn1 = 32'd693
; 
32'd26522: dataIn1 = 32'd714
; 
32'd26523: dataIn1 = 32'd744
; 
32'd26524: dataIn1 = 32'd765
; 
32'd26525: dataIn1 = 32'd797
; 
32'd26526: dataIn1 = 32'd649
; 
32'd26527: dataIn1 = 32'd651
; 
32'd26528: dataIn1 = 32'd671
; 
32'd26529: dataIn1 = 32'd672
; 
32'd26530: dataIn1 = 32'd709
; 
32'd26531: dataIn1 = 32'd723
; 
32'd26532: dataIn1 = 32'd732
; 
32'd26533: dataIn1 = 32'd783
; 
32'd26534: dataIn1 = 32'd785
; 
32'd26535: dataIn1 = 32'd786
; 
32'd26536: dataIn1 = 32'd796
; 
32'd26537: dataIn1 = 32'd652
; 
32'd26538: dataIn1 = 32'd682
; 
32'd26539: dataIn1 = 32'd687
; 
32'd26540: dataIn1 = 32'd690
; 
32'd26541: dataIn1 = 32'd698
; 
32'd26542: dataIn1 = 32'd725
; 
32'd26543: dataIn1 = 32'd789
; 
32'd26544: dataIn1 = 32'd794
; 
32'd26545: dataIn1 = 32'd797
; 
32'd26546: dataIn1 = 32'd650
; 
32'd26547: dataIn1 = 32'd753
; 
32'd26548: dataIn1 = 32'd771
; 
32'd26549: dataIn1 = 32'd777
; 
32'd26550: dataIn1 = 32'd656
; 
32'd26551: dataIn1 = 32'd657
; 
32'd26552: dataIn1 = 32'd704
; 
32'd26553: dataIn1 = 32'd731
; 
32'd26554: dataIn1 = 32'd733
; 
32'd26555: dataIn1 = 32'd752
; 
32'd26556: dataIn1 = 32'd754
; 
32'd26557: dataIn1 = 32'd787
; 
32'd26558: dataIn1 = 32'd652
; 
32'd26559: dataIn1 = 32'd681
; 
32'd26560: dataIn1 = 32'd694
; 
32'd26561: dataIn1 = 32'd700
; 
32'd26562: dataIn1 = 32'd709
; 
32'd26563: dataIn1 = 32'd712
; 
32'd26564: dataIn1 = 32'd714
; 
32'd26565: dataIn1 = 32'd724
; 
32'd26566: dataIn1 = 32'd763
; 
32'd26567: dataIn1 = 32'd665
; 
32'd26568: dataIn1 = 32'd673
; 
32'd26569: dataIn1 = 32'd681
; 
32'd26570: dataIn1 = 32'd692
; 
32'd26571: dataIn1 = 32'd730
; 
32'd26572: dataIn1 = 32'd746
; 
32'd26573: dataIn1 = 32'd772
; 
32'd26574: dataIn1 = 32'd688
; 
32'd26575: dataIn1 = 32'd696
; 
32'd26576: dataIn1 = 32'd701
; 
32'd26577: dataIn1 = 32'd705
; 
32'd26578: dataIn1 = 32'd708
; 
32'd26579: dataIn1 = 32'd713
; 
32'd26580: dataIn1 = 32'd714
; 
32'd26581: dataIn1 = 32'd730
; 
32'd26582: dataIn1 = 32'd755
; 
32'd26583: dataIn1 = 32'd768
; 
32'd26584: dataIn1 = 32'd778
; 
32'd26585: dataIn1 = 32'd662
; 
32'd26586: dataIn1 = 32'd675
; 
32'd26587: dataIn1 = 32'd720
; 
32'd26588: dataIn1 = 32'd745
; 
32'd26589: dataIn1 = 32'd767
; 
32'd26590: dataIn1 = 32'd776
; 
32'd26591: dataIn1 = 32'd665
; 
32'd26592: dataIn1 = 32'd668
; 
32'd26593: dataIn1 = 32'd698
; 
32'd26594: dataIn1 = 32'd730
; 
32'd26595: dataIn1 = 32'd757
; 
32'd26596: dataIn1 = 32'd793
; 
32'd26597: dataIn1 = 32'd795
; 
32'd26598: dataIn1 = 32'd799
; 
32'd26599: dataIn1 = 32'd689
; 
32'd26600: dataIn1 = 32'd691
; 
32'd26601: dataIn1 = 32'd693
; 
32'd26602: dataIn1 = 32'd696
; 
32'd26603: dataIn1 = 32'd699
; 
32'd26604: dataIn1 = 32'd705
; 
32'd26605: dataIn1 = 32'd715
; 
32'd26606: dataIn1 = 32'd749
; 
32'd26607: dataIn1 = 32'd759
; 
32'd26608: dataIn1 = 32'd782
; 
32'd26609: dataIn1 = 32'd788
; 
32'd26610: dataIn1 = 32'd799
; 
32'd26611: dataIn1 = 32'd675
; 
32'd26612: dataIn1 = 32'd702
; 
32'd26613: dataIn1 = 32'd715
; 
32'd26614: dataIn1 = 32'd717
; 
32'd26615: dataIn1 = 32'd720
; 
32'd26616: dataIn1 = 32'd724
; 
32'd26617: dataIn1 = 32'd745
; 
32'd26618: dataIn1 = 32'd756
; 
32'd26619: dataIn1 = 32'd778
; 
32'd26620: dataIn1 = 32'd665
; 
32'd26621: dataIn1 = 32'd666
; 
32'd26622: dataIn1 = 32'd682
; 
32'd26623: dataIn1 = 32'd697
; 
32'd26624: dataIn1 = 32'd698
; 
32'd26625: dataIn1 = 32'd710
; 
32'd26626: dataIn1 = 32'd717
; 
32'd26627: dataIn1 = 32'd724
; 
32'd26628: dataIn1 = 32'd762
; 
32'd26629: dataIn1 = 32'd790
; 
32'd26630: dataIn1 = 32'd671
; 
32'd26631: dataIn1 = 32'd674
; 
32'd26632: dataIn1 = 32'd686
; 
32'd26633: dataIn1 = 32'd687
; 
32'd26634: dataIn1 = 32'd726
; 
32'd26635: dataIn1 = 32'd735
; 
32'd26636: dataIn1 = 32'd744
; 
32'd26637: dataIn1 = 32'd752
; 
32'd26638: dataIn1 = 32'd797
; 
32'd26639: dataIn1 = 32'd675
; 
32'd26640: dataIn1 = 32'd681
; 
32'd26641: dataIn1 = 32'd712
; 
32'd26642: dataIn1 = 32'd739
; 
32'd26643: dataIn1 = 32'd780
; 
32'd26644: dataIn1 = 32'd786
; 
32'd26645: dataIn1 = 32'd794
; 
32'd26646: dataIn1 = 32'd673
; 
32'd26647: dataIn1 = 32'd678
; 
32'd26648: dataIn1 = 32'd703
; 
32'd26649: dataIn1 = 32'd706
; 
32'd26650: dataIn1 = 32'd743
; 
32'd26651: dataIn1 = 32'd754
; 
32'd26652: dataIn1 = 32'd796
; 
32'd26653: dataIn1 = 32'd686
; 
32'd26654: dataIn1 = 32'd699
; 
32'd26655: dataIn1 = 32'd707
; 
32'd26656: dataIn1 = 32'd708
; 
32'd26657: dataIn1 = 32'd745
; 
32'd26658: dataIn1 = 32'd791
; 
32'd26659: dataIn1 = 32'd669
; 
32'd26660: dataIn1 = 32'd693
; 
32'd26661: dataIn1 = 32'd700
; 
32'd26662: dataIn1 = 32'd724
; 
32'd26663: dataIn1 = 32'd733
; 
32'd26664: dataIn1 = 32'd752
; 
32'd26665: dataIn1 = 32'd756
; 
32'd26666: dataIn1 = 32'd794
; 
32'd26667: dataIn1 = 32'd796
; 
32'd26668: dataIn1 = 32'd665
; 
32'd26669: dataIn1 = 32'd669
; 
32'd26670: dataIn1 = 32'd674
; 
32'd26671: dataIn1 = 32'd699
; 
32'd26672: dataIn1 = 32'd703
; 
32'd26673: dataIn1 = 32'd709
; 
32'd26674: dataIn1 = 32'd757
; 
32'd26675: dataIn1 = 32'd791
; 
32'd26676: dataIn1 = 32'd680
; 
32'd26677: dataIn1 = 32'd702
; 
32'd26678: dataIn1 = 32'd703
; 
32'd26679: dataIn1 = 32'd706
; 
32'd26680: dataIn1 = 32'd724
; 
32'd26681: dataIn1 = 32'd799
; 
32'd26682: dataIn1 = 32'd686
; 
32'd26683: dataIn1 = 32'd713
; 
32'd26684: dataIn1 = 32'd723
; 
32'd26685: dataIn1 = 32'd738
; 
32'd26686: dataIn1 = 32'd742
; 
32'd26687: dataIn1 = 32'd744
; 
32'd26688: dataIn1 = 32'd781
; 
32'd26689: dataIn1 = 32'd687
; 
32'd26690: dataIn1 = 32'd689
; 
32'd26691: dataIn1 = 32'd702
; 
32'd26692: dataIn1 = 32'd717
; 
32'd26693: dataIn1 = 32'd725
; 
32'd26694: dataIn1 = 32'd731
; 
32'd26695: dataIn1 = 32'd753
; 
32'd26696: dataIn1 = 32'd787
; 
32'd26697: dataIn1 = 32'd788
; 
32'd26698: dataIn1 = 32'd793
; 
32'd26699: dataIn1 = 32'd707
; 
32'd26700: dataIn1 = 32'd710
; 
32'd26701: dataIn1 = 32'd736
; 
32'd26702: dataIn1 = 32'd753
; 
32'd26703: dataIn1 = 32'd754
; 
32'd26704: dataIn1 = 32'd764
; 
32'd26705: dataIn1 = 32'd770
; 
32'd26706: dataIn1 = 32'd771
; 
32'd26707: dataIn1 = 32'd772
; 
32'd26708: dataIn1 = 32'd777
; 
32'd26709: dataIn1 = 32'd780
; 
32'd26710: dataIn1 = 32'd785
; 
32'd26711: dataIn1 = 32'd685
; 
32'd26712: dataIn1 = 32'd700
; 
32'd26713: dataIn1 = 32'd737
; 
32'd26714: dataIn1 = 32'd767
; 
32'd26715: dataIn1 = 32'd790
; 
32'd26716: dataIn1 = 32'd673
; 
32'd26717: dataIn1 = 32'd675
; 
32'd26718: dataIn1 = 32'd687
; 
32'd26719: dataIn1 = 32'd693
; 
32'd26720: dataIn1 = 32'd697
; 
32'd26721: dataIn1 = 32'd746
; 
32'd26722: dataIn1 = 32'd764
; 
32'd26723: dataIn1 = 32'd767
; 
32'd26724: dataIn1 = 32'd677
; 
32'd26725: dataIn1 = 32'd706
; 
32'd26726: dataIn1 = 32'd735
; 
32'd26727: dataIn1 = 32'd743
; 
32'd26728: dataIn1 = 32'd751
; 
32'd26729: dataIn1 = 32'd773
; 
32'd26730: dataIn1 = 32'd779
; 
32'd26731: dataIn1 = 32'd679
; 
32'd26732: dataIn1 = 32'd716
; 
32'd26733: dataIn1 = 32'd733
; 
32'd26734: dataIn1 = 32'd758
; 
32'd26735: dataIn1 = 32'd769
; 
32'd26736: dataIn1 = 32'd696
; 
32'd26737: dataIn1 = 32'd727
; 
32'd26738: dataIn1 = 32'd748
; 
32'd26739: dataIn1 = 32'd753
; 
32'd26740: dataIn1 = 32'd759
; 
32'd26741: dataIn1 = 32'd764
; 
32'd26742: dataIn1 = 32'd767
; 
32'd26743: dataIn1 = 32'd774
; 
32'd26744: dataIn1 = 32'd782
; 
32'd26745: dataIn1 = 32'd795
; 
32'd26746: dataIn1 = 32'd798
; 
32'd26747: dataIn1 = 32'd683
; 
32'd26748: dataIn1 = 32'd700
; 
32'd26749: dataIn1 = 32'd721
; 
32'd26750: dataIn1 = 32'd724
; 
32'd26751: dataIn1 = 32'd729
; 
32'd26752: dataIn1 = 32'd770
; 
32'd26753: dataIn1 = 32'd788
; 
32'd26754: dataIn1 = 32'd687
; 
32'd26755: dataIn1 = 32'd748
; 
32'd26756: dataIn1 = 32'd777
; 
32'd26757: dataIn1 = 32'd789
; 
32'd26758: dataIn1 = 32'd798
; 
32'd26759: dataIn1 = 32'd685
; 
32'd26760: dataIn1 = 32'd696
; 
32'd26761: dataIn1 = 32'd707
; 
32'd26762: dataIn1 = 32'd708
; 
32'd26763: dataIn1 = 32'd738
; 
32'd26764: dataIn1 = 32'd747
; 
32'd26765: dataIn1 = 32'd756
; 
32'd26766: dataIn1 = 32'd680
; 
32'd26767: dataIn1 = 32'd686
; 
32'd26768: dataIn1 = 32'd703
; 
32'd26769: dataIn1 = 32'd727
; 
32'd26770: dataIn1 = 32'd763
; 
32'd26771: dataIn1 = 32'd779
; 
32'd26772: dataIn1 = 32'd692
; 
32'd26773: dataIn1 = 32'd755
; 
32'd26774: dataIn1 = 32'd798
; 
32'd26775: dataIn1 = 32'd717
; 
32'd26776: dataIn1 = 32'd723
; 
32'd26777: dataIn1 = 32'd730
; 
32'd26778: dataIn1 = 32'd734
; 
32'd26779: dataIn1 = 32'd735
; 
32'd26780: dataIn1 = 32'd743
; 
32'd26781: dataIn1 = 32'd784
; 
32'd26782: dataIn1 = 32'd786
; 
32'd26783: dataIn1 = 32'd725
; 
32'd26784: dataIn1 = 32'd754
; 
32'd26785: dataIn1 = 32'd760
; 
32'd26786: dataIn1 = 32'd775
; 
32'd26787: dataIn1 = 32'd780
; 
32'd26788: dataIn1 = 32'd798
; 
32'd26789: dataIn1 = 32'd684
; 
32'd26790: dataIn1 = 32'd687
; 
32'd26791: dataIn1 = 32'd695
; 
32'd26792: dataIn1 = 32'd748
; 
32'd26793: dataIn1 = 32'd751
; 
32'd26794: dataIn1 = 32'd758
; 
32'd26795: dataIn1 = 32'd759
; 
32'd26796: dataIn1 = 32'd782
; 
32'd26797: dataIn1 = 32'd688
; 
32'd26798: dataIn1 = 32'd698
; 
32'd26799: dataIn1 = 32'd717
; 
32'd26800: dataIn1 = 32'd733
; 
32'd26801: dataIn1 = 32'd736
; 
32'd26802: dataIn1 = 32'd771
; 
32'd26803: dataIn1 = 32'd698
; 
32'd26804: dataIn1 = 32'd710
; 
32'd26805: dataIn1 = 32'd711
; 
32'd26806: dataIn1 = 32'd712
; 
32'd26807: dataIn1 = 32'd737
; 
32'd26808: dataIn1 = 32'd740
; 
32'd26809: dataIn1 = 32'd779
; 
32'd26810: dataIn1 = 32'd784
; 
32'd26811: dataIn1 = 32'd798
; 
32'd26812: dataIn1 = 32'd692
; 
32'd26813: dataIn1 = 32'd698
; 
32'd26814: dataIn1 = 32'd729
; 
32'd26815: dataIn1 = 32'd735
; 
32'd26816: dataIn1 = 32'd744
; 
32'd26817: dataIn1 = 32'd763
; 
32'd26818: dataIn1 = 32'd778
; 
32'd26819: dataIn1 = 32'd798
; 
32'd26820: dataIn1 = 32'd690
; 
32'd26821: dataIn1 = 32'd701
; 
32'd26822: dataIn1 = 32'd717
; 
32'd26823: dataIn1 = 32'd718
; 
32'd26824: dataIn1 = 32'd773
; 
32'd26825: dataIn1 = 32'd782
; 
32'd26826: dataIn1 = 32'd716
; 
32'd26827: dataIn1 = 32'd743
; 
32'd26828: dataIn1 = 32'd745
; 
32'd26829: dataIn1 = 32'd753
; 
32'd26830: dataIn1 = 32'd754
; 
32'd26831: dataIn1 = 32'd761
; 
32'd26832: dataIn1 = 32'd768
; 
32'd26833: dataIn1 = 32'd784
; 
32'd26834: dataIn1 = 32'd703
; 
32'd26835: dataIn1 = 32'd742
; 
32'd26836: dataIn1 = 32'd748
; 
32'd26837: dataIn1 = 32'd757
; 
32'd26838: dataIn1 = 32'd759
; 
32'd26839: dataIn1 = 32'd770
; 
32'd26840: dataIn1 = 32'd780
; 
32'd26841: dataIn1 = 32'd784
; 
32'd26842: dataIn1 = 32'd796
; 
32'd26843: dataIn1 = 32'd797
; 
32'd26844: dataIn1 = 32'd713
; 
32'd26845: dataIn1 = 32'd722
; 
32'd26846: dataIn1 = 32'd731
; 
32'd26847: dataIn1 = 32'd732
; 
32'd26848: dataIn1 = 32'd740
; 
32'd26849: dataIn1 = 32'd742
; 
32'd26850: dataIn1 = 32'd758
; 
32'd26851: dataIn1 = 32'd761
; 
32'd26852: dataIn1 = 32'd699
; 
32'd26853: dataIn1 = 32'd707
; 
32'd26854: dataIn1 = 32'd727
; 
32'd26855: dataIn1 = 32'd733
; 
32'd26856: dataIn1 = 32'd752
; 
32'd26857: dataIn1 = 32'd709
; 
32'd26858: dataIn1 = 32'd730
; 
32'd26859: dataIn1 = 32'd740
; 
32'd26860: dataIn1 = 32'd756
; 
32'd26861: dataIn1 = 32'd764
; 
32'd26862: dataIn1 = 32'd771
; 
32'd26863: dataIn1 = 32'd784
; 
32'd26864: dataIn1 = 32'd708
; 
32'd26865: dataIn1 = 32'd756
; 
32'd26866: dataIn1 = 32'd764
; 
32'd26867: dataIn1 = 32'd693
; 
32'd26868: dataIn1 = 32'd695
; 
32'd26869: dataIn1 = 32'd696
; 
32'd26870: dataIn1 = 32'd753
; 
32'd26871: dataIn1 = 32'd728
; 
32'd26872: dataIn1 = 32'd746
; 
32'd26873: dataIn1 = 32'd776
; 
32'd26874: dataIn1 = 32'd781
; 
32'd26875: dataIn1 = 32'd749
; 
32'd26876: dataIn1 = 32'd778
; 
32'd26877: dataIn1 = 32'd780
; 
32'd26878: dataIn1 = 32'd798
; 
32'd26879: dataIn1 = 32'd721
; 
32'd26880: dataIn1 = 32'd769
; 
32'd26881: dataIn1 = 32'd773
; 
32'd26882: dataIn1 = 32'd775
; 
32'd26883: dataIn1 = 32'd786
; 
32'd26884: dataIn1 = 32'd703
; 
32'd26885: dataIn1 = 32'd710
; 
32'd26886: dataIn1 = 32'd724
; 
32'd26887: dataIn1 = 32'd725
; 
32'd26888: dataIn1 = 32'd790
; 
32'd26889: dataIn1 = 32'd791
; 
32'd26890: dataIn1 = 32'd795
; 
32'd26891: dataIn1 = 32'd704
; 
32'd26892: dataIn1 = 32'd706
; 
32'd26893: dataIn1 = 32'd707
; 
32'd26894: dataIn1 = 32'd710
; 
32'd26895: dataIn1 = 32'd717
; 
32'd26896: dataIn1 = 32'd746
; 
32'd26897: dataIn1 = 32'd763
; 
32'd26898: dataIn1 = 32'd797
; 
32'd26899: dataIn1 = 32'd707
; 
32'd26900: dataIn1 = 32'd713
; 
32'd26901: dataIn1 = 32'd727
; 
32'd26902: dataIn1 = 32'd762
; 
32'd26903: dataIn1 = 32'd771
; 
32'd26904: dataIn1 = 32'd749
; 
32'd26905: dataIn1 = 32'd780
; 
32'd26906: dataIn1 = 32'd781
; 
32'd26907: dataIn1 = 32'd787
; 
32'd26908: dataIn1 = 32'd800
; 
32'd26909: dataIn1 = 32'd704
; 
32'd26910: dataIn1 = 32'd706
; 
32'd26911: dataIn1 = 32'd711
; 
32'd26912: dataIn1 = 32'd725
; 
32'd26913: dataIn1 = 32'd745
; 
32'd26914: dataIn1 = 32'd757
; 
32'd26915: dataIn1 = 32'd762
; 
32'd26916: dataIn1 = 32'd771
; 
32'd26917: dataIn1 = 32'd777
; 
32'd26918: dataIn1 = 32'd787
; 
32'd26919: dataIn1 = 32'd797
; 
32'd26920: dataIn1 = 32'd742
; 
32'd26921: dataIn1 = 32'd768
; 
32'd26922: dataIn1 = 32'd780
; 
32'd26923: dataIn1 = 32'd794
; 
32'd26924: dataIn1 = 32'd800
; 
32'd26925: dataIn1 = 32'd728
; 
32'd26926: dataIn1 = 32'd739
; 
32'd26927: dataIn1 = 32'd752
; 
32'd26928: dataIn1 = 32'd755
; 
32'd26929: dataIn1 = 32'd773
; 
32'd26930: dataIn1 = 32'd774
; 
32'd26931: dataIn1 = 32'd712
; 
32'd26932: dataIn1 = 32'd724
; 
32'd26933: dataIn1 = 32'd726
; 
32'd26934: dataIn1 = 32'd750
; 
32'd26935: dataIn1 = 32'd751
; 
32'd26936: dataIn1 = 32'd726
; 
32'd26937: dataIn1 = 32'd740
; 
32'd26938: dataIn1 = 32'd756
; 
32'd26939: dataIn1 = 32'd768
; 
32'd26940: dataIn1 = 32'd775
; 
32'd26941: dataIn1 = 32'd778
; 
32'd26942: dataIn1 = 32'd708
; 
32'd26943: dataIn1 = 32'd726
; 
32'd26944: dataIn1 = 32'd736
; 
32'd26945: dataIn1 = 32'd768
; 
32'd26946: dataIn1 = 32'd773
; 
32'd26947: dataIn1 = 32'd777
; 
32'd26948: dataIn1 = 32'd787
; 
32'd26949: dataIn1 = 32'd726
; 
32'd26950: dataIn1 = 32'd718
; 
32'd26951: dataIn1 = 32'd727
; 
32'd26952: dataIn1 = 32'd764
; 
32'd26953: dataIn1 = 32'd779
; 
32'd26954: dataIn1 = 32'd784
; 
32'd26955: dataIn1 = 32'd797
; 
32'd26956: dataIn1 = 32'd800
; 
32'd26957: dataIn1 = 32'd758
; 
32'd26958: dataIn1 = 32'd765
; 
32'd26959: dataIn1 = 32'd767
; 
32'd26960: dataIn1 = 32'd769
; 
32'd26961: dataIn1 = 32'd770
; 
32'd26962: dataIn1 = 32'd718
; 
32'd26963: dataIn1 = 32'd769
; 
32'd26964: dataIn1 = 32'd771
; 
32'd26965: dataIn1 = 32'd782
; 
32'd26966: dataIn1 = 32'd785
; 
32'd26967: dataIn1 = 32'd751
; 
32'd26968: dataIn1 = 32'd759
; 
32'd26969: dataIn1 = 32'd772
; 
32'd26970: dataIn1 = 32'd717
; 
32'd26971: dataIn1 = 32'd750
; 
32'd26972: dataIn1 = 32'd782
; 
32'd26973: dataIn1 = 32'd789
; 
32'd26974: dataIn1 = 32'd791
; 
32'd26975: dataIn1 = 32'd713
; 
32'd26976: dataIn1 = 32'd719
; 
32'd26977: dataIn1 = 32'd720
; 
32'd26978: dataIn1 = 32'd726
; 
32'd26979: dataIn1 = 32'd735
; 
32'd26980: dataIn1 = 32'd769
; 
32'd26981: dataIn1 = 32'd787
; 
32'd26982: dataIn1 = 32'd800
; 
32'd26983: dataIn1 = 32'd718
; 
32'd26984: dataIn1 = 32'd738
; 
32'd26985: dataIn1 = 32'd752
; 
32'd26986: dataIn1 = 32'd765
; 
32'd26987: dataIn1 = 32'd768
; 
32'd26988: dataIn1 = 32'd773
; 
32'd26989: dataIn1 = 32'd777
; 
32'd26990: dataIn1 = 32'd718
; 
32'd26991: dataIn1 = 32'd721
; 
32'd26992: dataIn1 = 32'd735
; 
32'd26993: dataIn1 = 32'd742
; 
32'd26994: dataIn1 = 32'd745
; 
32'd26995: dataIn1 = 32'd753
; 
32'd26996: dataIn1 = 32'd755
; 
32'd26997: dataIn1 = 32'd776
; 
32'd26998: dataIn1 = 32'd784
; 
32'd26999: dataIn1 = 32'd729
; 
32'd27000: dataIn1 = 32'd736
; 
32'd27001: dataIn1 = 32'd744
; 
32'd27002: dataIn1 = 32'd763
; 
32'd27003: dataIn1 = 32'd794
; 
32'd27004: dataIn1 = 32'd767
; 
32'd27005: dataIn1 = 32'd789
; 
32'd27006: dataIn1 = 32'd729
; 
32'd27007: dataIn1 = 32'd732
; 
32'd27008: dataIn1 = 32'd751
; 
32'd27009: dataIn1 = 32'd787
; 
32'd27010: dataIn1 = 32'd736
; 
32'd27011: dataIn1 = 32'd754
; 
32'd27012: dataIn1 = 32'd758
; 
32'd27013: dataIn1 = 32'd775
; 
32'd27014: dataIn1 = 32'd781
; 
32'd27015: dataIn1 = 32'd783
; 
32'd27016: dataIn1 = 32'd748
; 
32'd27017: dataIn1 = 32'd773
; 
32'd27018: dataIn1 = 32'd785
; 
32'd27019: dataIn1 = 32'd792
; 
32'd27020: dataIn1 = 32'd722
; 
32'd27021: dataIn1 = 32'd732
; 
32'd27022: dataIn1 = 32'd750
; 
32'd27023: dataIn1 = 32'd795
; 
32'd27024: dataIn1 = 32'd749
; 
32'd27025: dataIn1 = 32'd766
; 
32'd27026: dataIn1 = 32'd771
; 
32'd27027: dataIn1 = 32'd794
; 
32'd27028: dataIn1 = 32'd784
; 
32'd27029: dataIn1 = 32'd793
; 
32'd27030: dataIn1 = 32'd725
; 
32'd27031: dataIn1 = 32'd743
; 
32'd27032: dataIn1 = 32'd775
; 
32'd27033: dataIn1 = 32'd788
; 
32'd27034: dataIn1 = 32'd791
; 
32'd27035: dataIn1 = 32'd800
; 
32'd27036: dataIn1 = 32'd728
; 
32'd27037: dataIn1 = 32'd783
; 
32'd27038: dataIn1 = 32'd738
; 
32'd27039: dataIn1 = 32'd759
; 
32'd27040: dataIn1 = 32'd761
; 
32'd27041: dataIn1 = 32'd770
; 
32'd27042: dataIn1 = 32'd777
; 
32'd27043: dataIn1 = 32'd783
; 
32'd27044: dataIn1 = 32'd788
; 
32'd27045: dataIn1 = 32'd747
; 
32'd27046: dataIn1 = 32'd769
; 
32'd27047: dataIn1 = 32'd771
; 
32'd27048: dataIn1 = 32'd780
; 
32'd27049: dataIn1 = 32'd784
; 
32'd27050: dataIn1 = 32'd742
; 
32'd27051: dataIn1 = 32'd746
; 
32'd27052: dataIn1 = 32'd770
; 
32'd27053: dataIn1 = 32'd793
; 
32'd27054: dataIn1 = 32'd795
; 
32'd27055: dataIn1 = 32'd755
; 
32'd27056: dataIn1 = 32'd757
; 
32'd27057: dataIn1 = 32'd758
; 
32'd27058: dataIn1 = 32'd762
; 
32'd27059: dataIn1 = 32'd800
; 
32'd27060: dataIn1 = 32'd748
; 
32'd27061: dataIn1 = 32'd761
; 
32'd27062: dataIn1 = 32'd765
; 
32'd27063: dataIn1 = 32'd788
; 
32'd27064: dataIn1 = 32'd740
; 
32'd27065: dataIn1 = 32'd756
; 
32'd27066: dataIn1 = 32'd768
; 
32'd27067: dataIn1 = 32'd764
; 
32'd27068: dataIn1 = 32'd780
; 
32'd27069: dataIn1 = 32'd786
; 
32'd27070: dataIn1 = 32'd790
; 
32'd27071: dataIn1 = 32'd798
; 
32'd27072: dataIn1 = 32'd791
; 
32'd27073: dataIn1 = 32'd797
; 
32'd27074: dataIn1 = 32'd764
; 
32'd27075: dataIn1 = 32'd788
; 
32'd27076: dataIn1 = 32'd745
; 
32'd27077: dataIn1 = 32'd750
; 
32'd27078: dataIn1 = 32'd773
; 
32'd27079: dataIn1 = 32'd776
; 
32'd27080: dataIn1 = 32'd797
; 
32'd27081: dataIn1 = 32'd800
; 
32'd27082: dataIn1 = 32'd741
; 
32'd27083: dataIn1 = 32'd748
; 
32'd27084: dataIn1 = 32'd750
; 
32'd27085: dataIn1 = 32'd753
; 
32'd27086: dataIn1 = 32'd790
; 
32'd27087: dataIn1 = 32'd798
; 
32'd27088: dataIn1 = 32'd759
; 
32'd27089: dataIn1 = 32'd761
; 
32'd27090: dataIn1 = 32'd764
; 
32'd27091: dataIn1 = 32'd784
; 
32'd27092: dataIn1 = 32'd790
; 
32'd27093: dataIn1 = 32'd794
; 
32'd27094: dataIn1 = 32'd798
; 
32'd27095: dataIn1 = 32'd744
; 
32'd27096: dataIn1 = 32'd795
; 
32'd27097: dataIn1 = 32'd778
; 
32'd27098: dataIn1 = 32'd743
; 
32'd27099: dataIn1 = 32'd758
; 
32'd27100: dataIn1 = 32'd767
; 
32'd27101: dataIn1 = 32'd794
; 
32'd27102: dataIn1 = 32'd743
; 
32'd27103: dataIn1 = 32'd776
; 
32'd27104: dataIn1 = 32'd786
; 
32'd27105: dataIn1 = 32'd795
; 
32'd27106: dataIn1 = 32'd751
; 
32'd27107: dataIn1 = 32'd780
; 
32'd27108: dataIn1 = 32'd786
; 
32'd27109: dataIn1 = 32'd797
; 
32'd27110: dataIn1 = 32'd749
; 
32'd27111: dataIn1 = 32'd751
; 
32'd27112: dataIn1 = 32'd755
; 
32'd27113: dataIn1 = 32'd757
; 
32'd27114: dataIn1 = 32'd765
; 
32'd27115: dataIn1 = 32'd795
; 
32'd27116: dataIn1 = 32'd753
; 
32'd27117: dataIn1 = 32'd784
; 
32'd27118: dataIn1 = 32'd748
; 
32'd27119: dataIn1 = 32'd763
; 
32'd27120: dataIn1 = 32'd768
; 
32'd27121: dataIn1 = 32'd772
; 
32'd27122: dataIn1 = 32'd782
; 
32'd27123: dataIn1 = 32'd759
; 
32'd27124: dataIn1 = 32'd772
; 
32'd27125: dataIn1 = 32'd756
; 
32'd27126: dataIn1 = 32'd757
; 
32'd27127: dataIn1 = 32'd762
; 
32'd27128: dataIn1 = 32'd768
; 
32'd27129: dataIn1 = 32'd793
; 
32'd27130: dataIn1 = 32'd759
; 
32'd27131: dataIn1 = 32'd765
; 
32'd27132: dataIn1 = 32'd777
; 
32'd27133: dataIn1 = 32'd756
; 
32'd27134: dataIn1 = 32'd764
; 
32'd27135: dataIn1 = 32'd777
; 
32'd27136: dataIn1 = 32'd789
; 
32'd27137: dataIn1 = 32'd754
; 
32'd27138: dataIn1 = 32'd755
; 
32'd27139: dataIn1 = 32'd783
; 
32'd27140: dataIn1 = 32'd789
; 
32'd27141: dataIn1 = 32'd792
; 
32'd27142: dataIn1 = 32'd799
; 
32'd27143: dataIn1 = 32'd790
; 
32'd27144: dataIn1 = 32'd791
; 
32'd27145: dataIn1 = 32'd762
; 
32'd27146: dataIn1 = 32'd783
; 
32'd27147: dataIn1 = 32'd762
; 
32'd27148: dataIn1 = 32'd788
; 
32'd27149: dataIn1 = 32'd797
; 
32'd27150: dataIn1 = 32'd775
; 
32'd27151: dataIn1 = 32'd789
; 
32'd27152: dataIn1 = 32'd800
; 
32'd27153: dataIn1 = 32'd770
; 
32'd27154: dataIn1 = 32'd781
; 
32'd27155: dataIn1 = 32'd784
; 
32'd27156: dataIn1 = 32'd772
; 
32'd27157: dataIn1 = 32'd774
; 
32'd27158: dataIn1 = 32'd784
; 
32'd27159: dataIn1 = 32'd786
; 
32'd27160: dataIn1 = 32'd791
; 
32'd27161: dataIn1 = 32'd776
; 
32'd27162: dataIn1 = 32'd785
; 
32'd27163: dataIn1 = 32'd799
; 
32'd27164: dataIn1 = 32'd776
; 
32'd27165: dataIn1 = 32'd800
; 
32'd27166: dataIn1 = 32'd779
; 
32'd27167: dataIn1 = 32'd783
; 
32'd27168: dataIn1 = 32'd796
; 
32'd27169: dataIn1 = 32'd778
; 
32'd27170: dataIn1 = 32'd788
; 
32'd27171: dataIn1 = 32'd776
; 
32'd27172: dataIn1 = 32'd798
; 
32'd27173: dataIn1 = 32'd798
; 
32'd27174: dataIn1 = 32'd787
; 
32'd27175: dataIn1 = 32'd788
; 
32'd27176: dataIn1 = 32'd795
; 
32'd27177: dataIn1 = 32'd795
; 
32'd27178: dataIn1 = 32'd800
; 
32'd27179: dataIn1 = 32'd782
; 
32'd27180: dataIn1 = 32'd786
; 
32'd27181: dataIn1 = 32'd800
; 
32'd27182: dataIn1 = 32'd786
; 
32'd27183: dataIn1 = 32'd797
; 
32'd27184: dataIn1 = 32'd785
; 
32'd27185: dataIn1 = 32'd788
; 
32'd27186: dataIn1 = 32'd788
; 
32'd27187: dataIn1 = 32'd793
; 
32'd27188: dataIn1 = 32'd795
; 
32'd27189: dataIn1 = 32'd800
; 
32'd27190: dataIn1 = 32'd792
; 
32'd27191: dataIn1 = 32'd798
; 
32'd27192: dataIn1 = 32'd796
; 
32'd27193: dataIn1 = 32'd799
; 
32'd27194: dataIn1 = 32'd798
; 
32'd27195: dataIn1 = 32'd800
; 
default:  
	dataIn1 = 32'd99999; 
endcase 
case(addr2) 
32'd2: dataIn2 = 32'd1; 
32'd3: dataIn2 = 32'd1; 
32'd4: dataIn2 = 32'd0; 
32'd5: dataIn2 = 32'd1; 
32'd6: dataIn2 = 32'd1; 
32'd7: dataIn2 = 32'd1; 
32'd8: dataIn2 = 32'd1; 
32'd9: dataIn2 = 32'd0; 
32'd10: dataIn2 = 32'd0; 
32'd11: dataIn2 = 32'd1; 
32'd12: dataIn2 = 32'd0; 
32'd13: dataIn2 = 32'd1; 
32'd14: dataIn2 = 32'd1; 
32'd15: dataIn2 = 32'd0; 
32'd16: dataIn2 = 32'd1; 
32'd17: dataIn2 = 32'd1; 
32'd18: dataIn2 = 32'd0; 
32'd19: dataIn2 = 32'd1; 
32'd20: dataIn2 = 32'd1; 
32'd21: dataIn2 = 32'd0; 
32'd22: dataIn2 = 32'd0; 
32'd23: dataIn2 = 32'd0; 
32'd24: dataIn2 = 32'd0; 
32'd25: dataIn2 = 32'd0; 
32'd26: dataIn2 = 32'd1; 
32'd27: dataIn2 = 32'd1; 
32'd28: dataIn2 = 32'd1; 
32'd29: dataIn2 = 32'd0; 
32'd30: dataIn2 = 32'd0; 
32'd31: dataIn2 = 32'd1; 
32'd32: dataIn2 = 32'd0; 
32'd33: dataIn2 = 32'd0; 
32'd34: dataIn2 = 32'd1; 
32'd35: dataIn2 = 32'd0; 
32'd36: dataIn2 = 32'd1; 
32'd37: dataIn2 = 32'd0; 
32'd38: dataIn2 = 32'd0; 
32'd39: dataIn2 = 32'd1; 
32'd40: dataIn2 = 32'd1; 
32'd41: dataIn2 = 32'd0; 
32'd42: dataIn2 = 32'd1; 
32'd43: dataIn2 = 32'd1; 
32'd44: dataIn2 = 32'd0; 
32'd45: dataIn2 = 32'd1; 
32'd46: dataIn2 = 32'd1; 
32'd47: dataIn2 = 32'd1; 
32'd48: dataIn2 = 32'd0; 
32'd49: dataIn2 = 32'd1; 
32'd50: dataIn2 = 32'd0; 
32'd51: dataIn2 = 32'd0; 
32'd52: dataIn2 = 32'd0; 
32'd53: dataIn2 = 32'd1; 
32'd54: dataIn2 = 32'd0; 
32'd55: dataIn2 = 32'd1; 
32'd56: dataIn2 = 32'd1; 
32'd57: dataIn2 = 32'd1; 
32'd58: dataIn2 = 32'd0; 
32'd59: dataIn2 = 32'd1; 
32'd60: dataIn2 = 32'd1; 
32'd61: dataIn2 = 32'd1; 
32'd62: dataIn2 = 32'd0; 
32'd63: dataIn2 = 32'd0; 
32'd64: dataIn2 = 32'd1; 
32'd65: dataIn2 = 32'd0; 
32'd66: dataIn2 = 32'd1; 
32'd67: dataIn2 = 32'd1; 
32'd68: dataIn2 = 32'd1; 
32'd69: dataIn2 = 32'd1; 
32'd70: dataIn2 = 32'd1; 
32'd71: dataIn2 = 32'd1; 
32'd72: dataIn2 = 32'd1; 
32'd73: dataIn2 = 32'd1; 
32'd74: dataIn2 = 32'd1; 
32'd75: dataIn2 = 32'd0; 
32'd76: dataIn2 = 32'd0; 
32'd77: dataIn2 = 32'd1; 
32'd78: dataIn2 = 32'd1; 
32'd79: dataIn2 = 32'd1; 
32'd80: dataIn2 = 32'd1; 
32'd81: dataIn2 = 32'd1; 
32'd82: dataIn2 = 32'd0; 
32'd83: dataIn2 = 32'd1; 
32'd84: dataIn2 = 32'd1; 
32'd85: dataIn2 = 32'd0; 
32'd86: dataIn2 = 32'd0; 
32'd87: dataIn2 = 32'd0; 
32'd88: dataIn2 = 32'd0; 
32'd89: dataIn2 = 32'd1; 
32'd90: dataIn2 = 32'd0; 
32'd91: dataIn2 = 32'd1; 
32'd92: dataIn2 = 32'd0; 
32'd93: dataIn2 = 32'd1; 
32'd94: dataIn2 = 32'd1; 
32'd95: dataIn2 = 32'd1; 
32'd96: dataIn2 = 32'd1; 
32'd97: dataIn2 = 32'd1; 
32'd98: dataIn2 = 32'd0; 
32'd99: dataIn2 = 32'd1; 
32'd100: dataIn2 = 32'd1; 
32'd101: dataIn2 = 32'd1; 
32'd102: dataIn2 = 32'd1; 
32'd103: dataIn2 = 32'd0; 
32'd104: dataIn2 = 32'd1; 
32'd105: dataIn2 = 32'd1; 
32'd106: dataIn2 = 32'd0; 
32'd107: dataIn2 = 32'd1; 
32'd108: dataIn2 = 32'd1; 
32'd109: dataIn2 = 32'd0; 
32'd110: dataIn2 = 32'd1; 
32'd111: dataIn2 = 32'd1; 
32'd112: dataIn2 = 32'd1; 
32'd113: dataIn2 = 32'd0; 
32'd114: dataIn2 = 32'd0; 
32'd115: dataIn2 = 32'd0; 
32'd116: dataIn2 = 32'd1; 
32'd117: dataIn2 = 32'd0; 
32'd118: dataIn2 = 32'd1; 
32'd119: dataIn2 = 32'd0; 
32'd120: dataIn2 = 32'd1; 
32'd121: dataIn2 = 32'd1; 
32'd122: dataIn2 = 32'd0; 
32'd123: dataIn2 = 32'd1; 
32'd124: dataIn2 = 32'd0; 
32'd125: dataIn2 = 32'd1; 
32'd126: dataIn2 = 32'd0; 
32'd127: dataIn2 = 32'd1; 
32'd128: dataIn2 = 32'd0; 
32'd129: dataIn2 = 32'd0; 
32'd130: dataIn2 = 32'd0; 
32'd131: dataIn2 = 32'd1; 
32'd132: dataIn2 = 32'd0; 
32'd133: dataIn2 = 32'd1; 
32'd134: dataIn2 = 32'd1; 
32'd135: dataIn2 = 32'd0; 
32'd136: dataIn2 = 32'd0; 
32'd137: dataIn2 = 32'd0; 
32'd138: dataIn2 = 32'd0; 
32'd139: dataIn2 = 32'd0; 
32'd140: dataIn2 = 32'd1; 
32'd141: dataIn2 = 32'd0; 
32'd142: dataIn2 = 32'd0; 
32'd143: dataIn2 = 32'd1; 
32'd144: dataIn2 = 32'd1; 
32'd145: dataIn2 = 32'd0; 
32'd146: dataIn2 = 32'd1; 
32'd147: dataIn2 = 32'd1; 
32'd148: dataIn2 = 32'd1; 
32'd149: dataIn2 = 32'd0; 
32'd150: dataIn2 = 32'd0; 
32'd151: dataIn2 = 32'd1; 
32'd152: dataIn2 = 32'd1; 
32'd153: dataIn2 = 32'd0; 
32'd154: dataIn2 = 32'd0; 
32'd155: dataIn2 = 32'd1; 
32'd156: dataIn2 = 32'd1; 
32'd157: dataIn2 = 32'd1; 
32'd158: dataIn2 = 32'd1; 
32'd159: dataIn2 = 32'd0; 
32'd160: dataIn2 = 32'd1; 
32'd161: dataIn2 = 32'd0; 
32'd162: dataIn2 = 32'd0; 
32'd163: dataIn2 = 32'd1; 
32'd164: dataIn2 = 32'd0; 
32'd165: dataIn2 = 32'd0; 
32'd166: dataIn2 = 32'd0; 
32'd167: dataIn2 = 32'd1; 
32'd168: dataIn2 = 32'd1; 
32'd169: dataIn2 = 32'd1; 
32'd170: dataIn2 = 32'd0; 
32'd171: dataIn2 = 32'd0; 
32'd172: dataIn2 = 32'd0; 
32'd173: dataIn2 = 32'd0; 
32'd174: dataIn2 = 32'd1; 
32'd175: dataIn2 = 32'd1; 
32'd176: dataIn2 = 32'd0; 
32'd177: dataIn2 = 32'd1; 
32'd178: dataIn2 = 32'd1; 
32'd179: dataIn2 = 32'd0; 
32'd180: dataIn2 = 32'd1; 
32'd181: dataIn2 = 32'd1; 
32'd182: dataIn2 = 32'd0; 
32'd183: dataIn2 = 32'd1; 
32'd184: dataIn2 = 32'd1; 
32'd185: dataIn2 = 32'd1; 
32'd186: dataIn2 = 32'd1; 
32'd187: dataIn2 = 32'd0; 
32'd188: dataIn2 = 32'd0; 
32'd189: dataIn2 = 32'd1; 
32'd190: dataIn2 = 32'd0; 
32'd191: dataIn2 = 32'd0; 
32'd192: dataIn2 = 32'd1; 
32'd193: dataIn2 = 32'd0; 
32'd194: dataIn2 = 32'd0; 
32'd195: dataIn2 = 32'd1; 
32'd196: dataIn2 = 32'd1; 
32'd197: dataIn2 = 32'd0; 
32'd198: dataIn2 = 32'd1; 
32'd199: dataIn2 = 32'd0; 
32'd200: dataIn2 = 32'd0; 
32'd201: dataIn2 = 32'd1; 
32'd202: dataIn2 = 32'd1; 
32'd203: dataIn2 = 32'd0; 
32'd204: dataIn2 = 32'd0; 
32'd205: dataIn2 = 32'd0; 
32'd206: dataIn2 = 32'd1; 
32'd207: dataIn2 = 32'd0; 
32'd208: dataIn2 = 32'd1; 
32'd209: dataIn2 = 32'd0; 
32'd210: dataIn2 = 32'd0; 
32'd211: dataIn2 = 32'd1; 
32'd212: dataIn2 = 32'd0; 
32'd213: dataIn2 = 32'd0; 
32'd214: dataIn2 = 32'd0; 
32'd215: dataIn2 = 32'd1; 
32'd216: dataIn2 = 32'd1; 
32'd217: dataIn2 = 32'd1; 
32'd218: dataIn2 = 32'd0; 
32'd219: dataIn2 = 32'd1; 
32'd220: dataIn2 = 32'd0; 
32'd221: dataIn2 = 32'd1; 
32'd222: dataIn2 = 32'd0; 
32'd223: dataIn2 = 32'd1; 
32'd224: dataIn2 = 32'd1; 
32'd225: dataIn2 = 32'd0; 
32'd226: dataIn2 = 32'd1; 
32'd227: dataIn2 = 32'd0; 
32'd228: dataIn2 = 32'd0; 
32'd229: dataIn2 = 32'd0; 
32'd230: dataIn2 = 32'd0; 
32'd231: dataIn2 = 32'd0; 
32'd232: dataIn2 = 32'd0; 
32'd233: dataIn2 = 32'd0; 
32'd234: dataIn2 = 32'd1; 
32'd235: dataIn2 = 32'd1; 
32'd236: dataIn2 = 32'd1; 
32'd237: dataIn2 = 32'd0; 
32'd238: dataIn2 = 32'd0; 
32'd239: dataIn2 = 32'd0; 
32'd240: dataIn2 = 32'd0; 
32'd241: dataIn2 = 32'd0; 
32'd242: dataIn2 = 32'd0; 
32'd243: dataIn2 = 32'd1; 
32'd244: dataIn2 = 32'd1; 
32'd245: dataIn2 = 32'd1; 
32'd246: dataIn2 = 32'd0; 
32'd247: dataIn2 = 32'd1; 
32'd248: dataIn2 = 32'd1; 
32'd249: dataIn2 = 32'd1; 
32'd250: dataIn2 = 32'd1; 
32'd251: dataIn2 = 32'd1; 
32'd252: dataIn2 = 32'd0; 
32'd253: dataIn2 = 32'd1; 
32'd254: dataIn2 = 32'd0; 
32'd255: dataIn2 = 32'd1; 
32'd256: dataIn2 = 32'd0; 
32'd257: dataIn2 = 32'd1; 
32'd258: dataIn2 = 32'd1; 
32'd259: dataIn2 = 32'd1; 
32'd260: dataIn2 = 32'd0; 
32'd261: dataIn2 = 32'd1; 
32'd262: dataIn2 = 32'd1; 
32'd263: dataIn2 = 32'd0; 
32'd264: dataIn2 = 32'd1; 
32'd265: dataIn2 = 32'd0; 
32'd266: dataIn2 = 32'd1; 
32'd267: dataIn2 = 32'd1; 
32'd268: dataIn2 = 32'd1; 
32'd269: dataIn2 = 32'd0; 
32'd270: dataIn2 = 32'd1; 
32'd271: dataIn2 = 32'd0; 
32'd272: dataIn2 = 32'd1; 
32'd273: dataIn2 = 32'd1; 
32'd274: dataIn2 = 32'd0; 
32'd275: dataIn2 = 32'd0; 
32'd276: dataIn2 = 32'd1; 
32'd277: dataIn2 = 32'd1; 
32'd278: dataIn2 = 32'd1; 
32'd279: dataIn2 = 32'd1; 
32'd280: dataIn2 = 32'd0; 
32'd281: dataIn2 = 32'd0; 
32'd282: dataIn2 = 32'd1; 
32'd283: dataIn2 = 32'd1; 
32'd284: dataIn2 = 32'd1; 
32'd285: dataIn2 = 32'd0; 
32'd286: dataIn2 = 32'd1; 
32'd287: dataIn2 = 32'd0; 
32'd288: dataIn2 = 32'd1; 
32'd289: dataIn2 = 32'd1; 
32'd290: dataIn2 = 32'd1; 
32'd291: dataIn2 = 32'd1; 
32'd292: dataIn2 = 32'd1; 
32'd293: dataIn2 = 32'd0; 
32'd294: dataIn2 = 32'd0; 
32'd295: dataIn2 = 32'd0; 
32'd296: dataIn2 = 32'd0; 
32'd297: dataIn2 = 32'd0; 
32'd298: dataIn2 = 32'd1; 
32'd299: dataIn2 = 32'd0; 
32'd300: dataIn2 = 32'd1; 
32'd301: dataIn2 = 32'd0; 
32'd302: dataIn2 = 32'd0; 
32'd303: dataIn2 = 32'd1; 
32'd304: dataIn2 = 32'd1; 
32'd305: dataIn2 = 32'd1; 
32'd306: dataIn2 = 32'd0; 
32'd307: dataIn2 = 32'd1; 
32'd308: dataIn2 = 32'd0; 
32'd309: dataIn2 = 32'd1; 
32'd310: dataIn2 = 32'd0; 
32'd311: dataIn2 = 32'd1; 
32'd312: dataIn2 = 32'd1; 
32'd313: dataIn2 = 32'd0; 
32'd314: dataIn2 = 32'd0; 
32'd315: dataIn2 = 32'd1; 
32'd316: dataIn2 = 32'd1; 
32'd317: dataIn2 = 32'd1; 
32'd318: dataIn2 = 32'd1; 
32'd319: dataIn2 = 32'd1; 
32'd320: dataIn2 = 32'd1; 
32'd321: dataIn2 = 32'd1; 
32'd322: dataIn2 = 32'd1; 
32'd323: dataIn2 = 32'd0; 
32'd324: dataIn2 = 32'd0; 
32'd325: dataIn2 = 32'd0; 
32'd326: dataIn2 = 32'd0; 
32'd327: dataIn2 = 32'd0; 
32'd328: dataIn2 = 32'd0; 
32'd329: dataIn2 = 32'd0; 
32'd330: dataIn2 = 32'd0; 
32'd331: dataIn2 = 32'd0; 
32'd332: dataIn2 = 32'd1; 
32'd333: dataIn2 = 32'd0; 
32'd334: dataIn2 = 32'd1; 
32'd335: dataIn2 = 32'd1; 
32'd336: dataIn2 = 32'd1; 
32'd337: dataIn2 = 32'd1; 
32'd338: dataIn2 = 32'd1; 
32'd339: dataIn2 = 32'd0; 
32'd340: dataIn2 = 32'd0; 
32'd341: dataIn2 = 32'd0; 
32'd342: dataIn2 = 32'd1; 
32'd343: dataIn2 = 32'd0; 
32'd344: dataIn2 = 32'd1; 
32'd345: dataIn2 = 32'd0; 
32'd346: dataIn2 = 32'd0; 
32'd347: dataIn2 = 32'd1; 
32'd348: dataIn2 = 32'd1; 
32'd349: dataIn2 = 32'd1; 
32'd350: dataIn2 = 32'd0; 
32'd351: dataIn2 = 32'd0; 
32'd352: dataIn2 = 32'd1; 
32'd353: dataIn2 = 32'd1; 
32'd354: dataIn2 = 32'd1; 
32'd355: dataIn2 = 32'd1; 
32'd356: dataIn2 = 32'd0; 
32'd357: dataIn2 = 32'd1; 
32'd358: dataIn2 = 32'd0; 
32'd359: dataIn2 = 32'd1; 
32'd360: dataIn2 = 32'd0; 
32'd361: dataIn2 = 32'd0; 
32'd362: dataIn2 = 32'd0; 
32'd363: dataIn2 = 32'd1; 
32'd364: dataIn2 = 32'd0; 
32'd365: dataIn2 = 32'd1; 
32'd366: dataIn2 = 32'd0; 
32'd367: dataIn2 = 32'd1; 
32'd368: dataIn2 = 32'd1; 
32'd369: dataIn2 = 32'd0; 
32'd370: dataIn2 = 32'd1; 
32'd371: dataIn2 = 32'd1; 
32'd372: dataIn2 = 32'd0; 
32'd373: dataIn2 = 32'd1; 
32'd374: dataIn2 = 32'd1; 
32'd375: dataIn2 = 32'd0; 
32'd376: dataIn2 = 32'd1; 
32'd377: dataIn2 = 32'd0; 
32'd378: dataIn2 = 32'd0; 
32'd379: dataIn2 = 32'd0; 
32'd380: dataIn2 = 32'd0; 
32'd381: dataIn2 = 32'd0; 
32'd382: dataIn2 = 32'd0; 
32'd383: dataIn2 = 32'd1; 
32'd384: dataIn2 = 32'd0; 
32'd385: dataIn2 = 32'd1; 
32'd386: dataIn2 = 32'd1; 
32'd387: dataIn2 = 32'd0; 
32'd388: dataIn2 = 32'd0; 
32'd389: dataIn2 = 32'd0; 
32'd390: dataIn2 = 32'd1; 
32'd391: dataIn2 = 32'd1; 
32'd392: dataIn2 = 32'd1; 
32'd393: dataIn2 = 32'd1; 
32'd394: dataIn2 = 32'd0; 
32'd395: dataIn2 = 32'd0; 
32'd396: dataIn2 = 32'd0; 
32'd397: dataIn2 = 32'd1; 
32'd398: dataIn2 = 32'd1; 
32'd399: dataIn2 = 32'd1; 
32'd400: dataIn2 = 32'd0; 
32'd401: dataIn2 = 32'd1; 
32'd402: dataIn2 = 32'd0; 
32'd403: dataIn2 = 32'd0; 
32'd404: dataIn2 = 32'd1; 
32'd405: dataIn2 = 32'd1; 
32'd406: dataIn2 = 32'd0; 
32'd407: dataIn2 = 32'd0; 
32'd408: dataIn2 = 32'd0; 
32'd409: dataIn2 = 32'd0; 
32'd410: dataIn2 = 32'd1; 
32'd411: dataIn2 = 32'd1; 
32'd412: dataIn2 = 32'd1; 
32'd413: dataIn2 = 32'd1; 
32'd414: dataIn2 = 32'd1; 
32'd415: dataIn2 = 32'd0; 
32'd416: dataIn2 = 32'd0; 
32'd417: dataIn2 = 32'd1; 
32'd418: dataIn2 = 32'd0; 
32'd419: dataIn2 = 32'd1; 
32'd420: dataIn2 = 32'd1; 
32'd421: dataIn2 = 32'd1; 
32'd422: dataIn2 = 32'd1; 
32'd423: dataIn2 = 32'd1; 
32'd424: dataIn2 = 32'd0; 
32'd425: dataIn2 = 32'd1; 
32'd426: dataIn2 = 32'd0; 
32'd427: dataIn2 = 32'd0; 
32'd428: dataIn2 = 32'd0; 
32'd429: dataIn2 = 32'd0; 
32'd430: dataIn2 = 32'd0; 
32'd431: dataIn2 = 32'd1; 
32'd432: dataIn2 = 32'd0; 
32'd433: dataIn2 = 32'd0; 
32'd434: dataIn2 = 32'd0; 
32'd435: dataIn2 = 32'd1; 
32'd436: dataIn2 = 32'd1; 
32'd437: dataIn2 = 32'd0; 
32'd438: dataIn2 = 32'd1; 
32'd439: dataIn2 = 32'd1; 
32'd440: dataIn2 = 32'd0; 
32'd441: dataIn2 = 32'd1; 
32'd442: dataIn2 = 32'd0; 
32'd443: dataIn2 = 32'd0; 
32'd444: dataIn2 = 32'd1; 
32'd445: dataIn2 = 32'd1; 
32'd446: dataIn2 = 32'd0; 
32'd447: dataIn2 = 32'd0; 
32'd448: dataIn2 = 32'd1; 
32'd449: dataIn2 = 32'd0; 
32'd450: dataIn2 = 32'd0; 
32'd451: dataIn2 = 32'd0; 
32'd452: dataIn2 = 32'd0; 
32'd453: dataIn2 = 32'd1; 
32'd454: dataIn2 = 32'd1; 
32'd455: dataIn2 = 32'd0; 
32'd456: dataIn2 = 32'd1; 
32'd457: dataIn2 = 32'd1; 
32'd458: dataIn2 = 32'd1; 
32'd459: dataIn2 = 32'd0; 
32'd460: dataIn2 = 32'd0; 
32'd461: dataIn2 = 32'd1; 
32'd462: dataIn2 = 32'd1; 
32'd463: dataIn2 = 32'd1; 
32'd464: dataIn2 = 32'd1; 
32'd465: dataIn2 = 32'd0; 
32'd466: dataIn2 = 32'd0; 
32'd467: dataIn2 = 32'd0; 
32'd468: dataIn2 = 32'd1; 
32'd469: dataIn2 = 32'd1; 
32'd470: dataIn2 = 32'd1; 
32'd471: dataIn2 = 32'd0; 
32'd472: dataIn2 = 32'd1; 
32'd473: dataIn2 = 32'd1; 
32'd474: dataIn2 = 32'd0; 
32'd475: dataIn2 = 32'd1; 
32'd476: dataIn2 = 32'd1; 
32'd477: dataIn2 = 32'd0; 
32'd478: dataIn2 = 32'd0; 
32'd479: dataIn2 = 32'd1; 
32'd480: dataIn2 = 32'd1; 
32'd481: dataIn2 = 32'd1; 
32'd482: dataIn2 = 32'd0; 
32'd483: dataIn2 = 32'd0; 
32'd484: dataIn2 = 32'd0; 
32'd485: dataIn2 = 32'd1; 
32'd486: dataIn2 = 32'd0; 
32'd487: dataIn2 = 32'd0; 
32'd488: dataIn2 = 32'd1; 
32'd489: dataIn2 = 32'd0; 
32'd490: dataIn2 = 32'd1; 
32'd491: dataIn2 = 32'd0; 
32'd492: dataIn2 = 32'd0; 
32'd493: dataIn2 = 32'd0; 
32'd494: dataIn2 = 32'd0; 
32'd495: dataIn2 = 32'd0; 
32'd496: dataIn2 = 32'd0; 
32'd497: dataIn2 = 32'd1; 
32'd498: dataIn2 = 32'd0; 
32'd499: dataIn2 = 32'd0; 
32'd500: dataIn2 = 32'd0; 
32'd501: dataIn2 = 32'd0; 
32'd502: dataIn2 = 32'd0; 
32'd503: dataIn2 = 32'd1; 
32'd504: dataIn2 = 32'd1; 
32'd505: dataIn2 = 32'd1; 
32'd506: dataIn2 = 32'd1; 
32'd507: dataIn2 = 32'd0; 
32'd508: dataIn2 = 32'd0; 
32'd509: dataIn2 = 32'd1; 
32'd510: dataIn2 = 32'd0; 
32'd511: dataIn2 = 32'd0; 
32'd512: dataIn2 = 32'd0; 
32'd513: dataIn2 = 32'd0; 
32'd514: dataIn2 = 32'd0; 
32'd515: dataIn2 = 32'd1; 
32'd516: dataIn2 = 32'd0; 
32'd517: dataIn2 = 32'd0; 
32'd518: dataIn2 = 32'd0; 
32'd519: dataIn2 = 32'd0; 
32'd520: dataIn2 = 32'd1; 
32'd521: dataIn2 = 32'd0; 
32'd522: dataIn2 = 32'd1; 
32'd523: dataIn2 = 32'd0; 
32'd524: dataIn2 = 32'd1; 
32'd525: dataIn2 = 32'd0; 
32'd526: dataIn2 = 32'd0; 
32'd527: dataIn2 = 32'd1; 
32'd528: dataIn2 = 32'd0; 
32'd529: dataIn2 = 32'd1; 
32'd530: dataIn2 = 32'd0; 
32'd531: dataIn2 = 32'd0; 
32'd532: dataIn2 = 32'd1; 
32'd533: dataIn2 = 32'd0; 
32'd534: dataIn2 = 32'd1; 
32'd535: dataIn2 = 32'd1; 
32'd536: dataIn2 = 32'd0; 
32'd537: dataIn2 = 32'd0; 
32'd538: dataIn2 = 32'd0; 
32'd539: dataIn2 = 32'd0; 
32'd540: dataIn2 = 32'd0; 
32'd541: dataIn2 = 32'd1; 
32'd542: dataIn2 = 32'd1; 
32'd543: dataIn2 = 32'd0; 
32'd544: dataIn2 = 32'd1; 
32'd545: dataIn2 = 32'd1; 
32'd546: dataIn2 = 32'd1; 
32'd547: dataIn2 = 32'd0; 
32'd548: dataIn2 = 32'd0; 
32'd549: dataIn2 = 32'd1; 
32'd550: dataIn2 = 32'd1; 
32'd551: dataIn2 = 32'd1; 
32'd552: dataIn2 = 32'd0; 
32'd553: dataIn2 = 32'd0; 
32'd554: dataIn2 = 32'd1; 
32'd555: dataIn2 = 32'd1; 
32'd556: dataIn2 = 32'd0; 
32'd557: dataIn2 = 32'd1; 
32'd558: dataIn2 = 32'd1; 
32'd559: dataIn2 = 32'd0; 
32'd560: dataIn2 = 32'd0; 
32'd561: dataIn2 = 32'd0; 
32'd562: dataIn2 = 32'd1; 
32'd563: dataIn2 = 32'd0; 
32'd564: dataIn2 = 32'd0; 
32'd565: dataIn2 = 32'd0; 
32'd566: dataIn2 = 32'd1; 
32'd567: dataIn2 = 32'd1; 
32'd568: dataIn2 = 32'd1; 
32'd569: dataIn2 = 32'd1; 
32'd570: dataIn2 = 32'd1; 
32'd571: dataIn2 = 32'd1; 
32'd572: dataIn2 = 32'd0; 
32'd573: dataIn2 = 32'd1; 
32'd574: dataIn2 = 32'd1; 
32'd575: dataIn2 = 32'd1; 
32'd576: dataIn2 = 32'd0; 
32'd577: dataIn2 = 32'd1; 
32'd578: dataIn2 = 32'd0; 
32'd579: dataIn2 = 32'd0; 
32'd580: dataIn2 = 32'd0; 
32'd581: dataIn2 = 32'd1; 
32'd582: dataIn2 = 32'd0; 
32'd583: dataIn2 = 32'd0; 
32'd584: dataIn2 = 32'd1; 
32'd585: dataIn2 = 32'd0; 
32'd586: dataIn2 = 32'd1; 
32'd587: dataIn2 = 32'd1; 
32'd588: dataIn2 = 32'd0; 
32'd589: dataIn2 = 32'd0; 
32'd590: dataIn2 = 32'd0; 
32'd591: dataIn2 = 32'd0; 
32'd592: dataIn2 = 32'd1; 
32'd593: dataIn2 = 32'd1; 
32'd594: dataIn2 = 32'd1; 
32'd595: dataIn2 = 32'd1; 
32'd596: dataIn2 = 32'd0; 
32'd597: dataIn2 = 32'd0; 
32'd598: dataIn2 = 32'd0; 
32'd599: dataIn2 = 32'd0; 
32'd600: dataIn2 = 32'd0; 
32'd601: dataIn2 = 32'd0; 
32'd602: dataIn2 = 32'd0; 
32'd603: dataIn2 = 32'd0; 
32'd604: dataIn2 = 32'd0; 
32'd605: dataIn2 = 32'd0; 
32'd606: dataIn2 = 32'd1; 
32'd607: dataIn2 = 32'd0; 
32'd608: dataIn2 = 32'd0; 
32'd609: dataIn2 = 32'd0; 
32'd610: dataIn2 = 32'd0; 
32'd611: dataIn2 = 32'd1; 
32'd612: dataIn2 = 32'd1; 
32'd613: dataIn2 = 32'd0; 
32'd614: dataIn2 = 32'd1; 
32'd615: dataIn2 = 32'd0; 
32'd616: dataIn2 = 32'd0; 
32'd617: dataIn2 = 32'd0; 
32'd618: dataIn2 = 32'd1; 
32'd619: dataIn2 = 32'd0; 
32'd620: dataIn2 = 32'd0; 
32'd621: dataIn2 = 32'd1; 
32'd622: dataIn2 = 32'd0; 
32'd623: dataIn2 = 32'd0; 
32'd624: dataIn2 = 32'd0; 
32'd625: dataIn2 = 32'd1; 
32'd626: dataIn2 = 32'd0; 
32'd627: dataIn2 = 32'd0; 
32'd628: dataIn2 = 32'd0; 
32'd629: dataIn2 = 32'd1; 
32'd630: dataIn2 = 32'd1; 
32'd631: dataIn2 = 32'd1; 
32'd632: dataIn2 = 32'd1; 
32'd633: dataIn2 = 32'd0; 
32'd634: dataIn2 = 32'd1; 
32'd635: dataIn2 = 32'd1; 
32'd636: dataIn2 = 32'd1; 
32'd637: dataIn2 = 32'd1; 
32'd638: dataIn2 = 32'd0; 
32'd639: dataIn2 = 32'd1; 
32'd640: dataIn2 = 32'd1; 
32'd641: dataIn2 = 32'd1; 
32'd642: dataIn2 = 32'd0; 
32'd643: dataIn2 = 32'd1; 
32'd644: dataIn2 = 32'd0; 
32'd645: dataIn2 = 32'd0; 
32'd646: dataIn2 = 32'd1; 
32'd647: dataIn2 = 32'd1; 
32'd648: dataIn2 = 32'd0; 
32'd649: dataIn2 = 32'd1; 
32'd650: dataIn2 = 32'd0; 
32'd651: dataIn2 = 32'd0; 
32'd652: dataIn2 = 32'd0; 
32'd653: dataIn2 = 32'd0; 
32'd654: dataIn2 = 32'd1; 
32'd655: dataIn2 = 32'd0; 
32'd656: dataIn2 = 32'd1; 
32'd657: dataIn2 = 32'd0; 
32'd658: dataIn2 = 32'd0; 
32'd659: dataIn2 = 32'd1; 
32'd660: dataIn2 = 32'd0; 
32'd661: dataIn2 = 32'd0; 
32'd662: dataIn2 = 32'd0; 
32'd663: dataIn2 = 32'd0; 
32'd664: dataIn2 = 32'd1; 
32'd665: dataIn2 = 32'd0; 
32'd666: dataIn2 = 32'd0; 
32'd667: dataIn2 = 32'd0; 
32'd668: dataIn2 = 32'd1; 
32'd669: dataIn2 = 32'd1; 
32'd670: dataIn2 = 32'd1; 
32'd671: dataIn2 = 32'd1; 
32'd672: dataIn2 = 32'd0; 
32'd673: dataIn2 = 32'd0; 
32'd674: dataIn2 = 32'd0; 
32'd675: dataIn2 = 32'd0; 
32'd676: dataIn2 = 32'd1; 
32'd677: dataIn2 = 32'd0; 
32'd678: dataIn2 = 32'd0; 
32'd679: dataIn2 = 32'd1; 
32'd680: dataIn2 = 32'd1; 
32'd681: dataIn2 = 32'd0; 
32'd682: dataIn2 = 32'd1; 
32'd683: dataIn2 = 32'd1; 
32'd684: dataIn2 = 32'd0; 
32'd685: dataIn2 = 32'd1; 
32'd686: dataIn2 = 32'd0; 
32'd687: dataIn2 = 32'd1; 
32'd688: dataIn2 = 32'd1; 
32'd689: dataIn2 = 32'd0; 
32'd690: dataIn2 = 32'd0; 
32'd691: dataIn2 = 32'd0; 
32'd692: dataIn2 = 32'd1; 
32'd693: dataIn2 = 32'd0; 
32'd694: dataIn2 = 32'd0; 
32'd695: dataIn2 = 32'd0; 
32'd696: dataIn2 = 32'd0; 
32'd697: dataIn2 = 32'd0; 
32'd698: dataIn2 = 32'd1; 
32'd699: dataIn2 = 32'd1; 
32'd700: dataIn2 = 32'd1; 
32'd701: dataIn2 = 32'd0; 
32'd702: dataIn2 = 32'd1; 
32'd703: dataIn2 = 32'd0; 
32'd704: dataIn2 = 32'd0; 
32'd705: dataIn2 = 32'd0; 
32'd706: dataIn2 = 32'd0; 
32'd707: dataIn2 = 32'd1; 
32'd708: dataIn2 = 32'd0; 
32'd709: dataIn2 = 32'd1; 
32'd710: dataIn2 = 32'd1; 
32'd711: dataIn2 = 32'd0; 
32'd712: dataIn2 = 32'd1; 
32'd713: dataIn2 = 32'd0; 
32'd714: dataIn2 = 32'd0; 
32'd715: dataIn2 = 32'd1; 
32'd716: dataIn2 = 32'd0; 
32'd717: dataIn2 = 32'd1; 
32'd718: dataIn2 = 32'd1; 
32'd719: dataIn2 = 32'd0; 
32'd720: dataIn2 = 32'd1; 
32'd721: dataIn2 = 32'd1; 
32'd722: dataIn2 = 32'd1; 
32'd723: dataIn2 = 32'd0; 
32'd724: dataIn2 = 32'd1; 
32'd725: dataIn2 = 32'd1; 
32'd726: dataIn2 = 32'd0; 
32'd727: dataIn2 = 32'd1; 
32'd728: dataIn2 = 32'd0; 
32'd729: dataIn2 = 32'd0; 
32'd730: dataIn2 = 32'd1; 
32'd731: dataIn2 = 32'd0; 
32'd732: dataIn2 = 32'd0; 
32'd733: dataIn2 = 32'd0; 
32'd734: dataIn2 = 32'd0; 
32'd735: dataIn2 = 32'd1; 
32'd736: dataIn2 = 32'd1; 
32'd737: dataIn2 = 32'd1; 
32'd738: dataIn2 = 32'd1; 
32'd739: dataIn2 = 32'd0; 
32'd740: dataIn2 = 32'd0; 
32'd741: dataIn2 = 32'd0; 
32'd742: dataIn2 = 32'd1; 
32'd743: dataIn2 = 32'd0; 
32'd744: dataIn2 = 32'd0; 
32'd745: dataIn2 = 32'd1; 
32'd746: dataIn2 = 32'd1; 
32'd747: dataIn2 = 32'd0; 
32'd748: dataIn2 = 32'd0; 
32'd749: dataIn2 = 32'd0; 
32'd750: dataIn2 = 32'd1; 
32'd751: dataIn2 = 32'd1; 
32'd752: dataIn2 = 32'd1; 
32'd753: dataIn2 = 32'd1; 
32'd754: dataIn2 = 32'd1; 
32'd755: dataIn2 = 32'd0; 
32'd756: dataIn2 = 32'd0; 
32'd757: dataIn2 = 32'd0; 
32'd758: dataIn2 = 32'd1; 
32'd759: dataIn2 = 32'd0; 
32'd760: dataIn2 = 32'd1; 
32'd761: dataIn2 = 32'd1; 
32'd762: dataIn2 = 32'd1; 
32'd763: dataIn2 = 32'd1; 
32'd764: dataIn2 = 32'd1; 
32'd765: dataIn2 = 32'd1; 
32'd766: dataIn2 = 32'd0; 
32'd767: dataIn2 = 32'd0; 
32'd768: dataIn2 = 32'd1; 
32'd769: dataIn2 = 32'd1; 
32'd770: dataIn2 = 32'd0; 
32'd771: dataIn2 = 32'd0; 
32'd772: dataIn2 = 32'd0; 
32'd773: dataIn2 = 32'd1; 
32'd774: dataIn2 = 32'd1; 
32'd775: dataIn2 = 32'd0; 
32'd776: dataIn2 = 32'd0; 
32'd777: dataIn2 = 32'd1; 
32'd778: dataIn2 = 32'd0; 
32'd779: dataIn2 = 32'd0; 
32'd780: dataIn2 = 32'd0; 
32'd781: dataIn2 = 32'd1; 
32'd782: dataIn2 = 32'd1; 
32'd783: dataIn2 = 32'd0; 
32'd784: dataIn2 = 32'd0; 
32'd785: dataIn2 = 32'd0; 
32'd786: dataIn2 = 32'd1; 
32'd787: dataIn2 = 32'd1; 
32'd788: dataIn2 = 32'd1; 
32'd789: dataIn2 = 32'd0; 
32'd790: dataIn2 = 32'd1; 
32'd791: dataIn2 = 32'd1; 
32'd792: dataIn2 = 32'd1; 
32'd793: dataIn2 = 32'd0; 
32'd794: dataIn2 = 32'd0; 
32'd795: dataIn2 = 32'd1; 
32'd796: dataIn2 = 32'd1; 
32'd797: dataIn2 = 32'd0; 
32'd798: dataIn2 = 32'd1; 
32'd799: dataIn2 = 32'd0; 
32'd800: dataIn2 = 32'd1; 
32'd801: dataIn2 = 32'd0; 
default: 
	dataIn2 = 32'd99999; 
endcase 
end 
always begin 
#10 Clk = ~Clk; 
end 
//========== VCD ============ 
`ifdef VCD 
initial 
begin 
	$dumpfile("g10.vcd");  
	$dumpvars; 
end 
`endif 
//===========RTLVCD ========== 
`ifdef RTLVCD 
initial 
begin 
	$dumpfile("hht_rtl.vcd"); 
	$dumpvars; 
end 
`endif 
endmodule 
