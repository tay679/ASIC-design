//991x991 
// Code your testbench here 
// or browse Examples 
// Verilog test bench for HHT with buffer 
`timescale 1ns/1ps 
module testbench; 
  parameter V_SIZE = 9; 
  parameter COL_SIZE = 6027 ; 
reg Clk,Rst,WR,mem_init; 
reg [31:0] dataIn1,dataIn2,csize; 
reg [31:0]v_values_base; 
wire [31:0]addr1,addr2; 
wire [4:0] regaddr1,regaddr2; 
reg[31:0] cpu_addr;
wire hht;
wire [31:0]val[0:8]; 
reg [31:0]wdata_col_base; 
wire [31:0] dataOut; 
reg fe_init; 
reg wn,rn,RD; 
wire [4:0]adata; 
wire [31:0] rdata; 
 // Instantiate memory module 
//  memmodel m1 (addr,dataIn,dataOut,WR,Clk,Rst); 
//  mem_buffer m1 (dataOut, full, empty, Clk, Rst, wn, rn, dataIn); 
control t1 (Clk,wdata_col_base,v_values_base,addr1,addr2,dataIn1,dataIn2,Rst,RD,csize,cpu_addr,hht,regaddr1,regaddr2,rdata,adata); ;  
//frontend t1 (Clk,Rst,fe_init,wdata_col_base,data_req,dataIn,init, 
//{m_cols[0],m_cols[1],m_cols[2],m_cols[3],m_cols[4]}, 
//done,wn); 
initial begin 
Clk = 1'b0; 
  RD = 1'b1; 
 #15; 
Rst = 1'b0; 
cpu_addr = 32'd126;
  v_values_base = 32'd2; 
  wdata_col_base = 32'd9930 ; 
  csize = COL_SIZE; 
 fe_init = 1'b1; 
#15 Rst = 1'b1; 
// RD = 1'b0; 
// RD = 1'b1; 
 #1320000; 
$finish; 
end 
always @(*) begin 
//$display("%b,%b",t1.fe1.count,t1.fe1.vdata_req); 
case(addr1)  
32'd9930: dataIn1 = 32'd1
; 
32'd9931: dataIn1 = 32'd84
; 
32'd9932: dataIn1 = 32'd2
; 
32'd9933: dataIn1 = 32'd85
; 
32'd9934: dataIn1 = 32'd122
; 
32'd9935: dataIn1 = 32'd147
; 
32'd9936: dataIn1 = 32'd165
; 
32'd9937: dataIn1 = 32'd3
; 
32'd9938: dataIn1 = 32'd122
; 
32'd9939: dataIn1 = 32'd4
; 
32'd9940: dataIn1 = 32'd122
; 
32'd9941: dataIn1 = 32'd123
; 
32'd9942: dataIn1 = 32'd141
; 
32'd9943: dataIn1 = 32'd5
; 
32'd9944: dataIn1 = 32'd85
; 
32'd9945: dataIn1 = 32'd123
; 
32'd9946: dataIn1 = 32'd6
; 
32'd9947: dataIn1 = 32'd7
; 
32'd9948: dataIn1 = 32'd101
; 
32'd9949: dataIn1 = 32'd124
; 
32'd9950: dataIn1 = 32'd8
; 
32'd9951: dataIn1 = 32'd107
; 
32'd9952: dataIn1 = 32'd124
; 
32'd9953: dataIn1 = 32'd125
; 
32'd9954: dataIn1 = 32'd9
; 
32'd9955: dataIn1 = 32'd107
; 
32'd9956: dataIn1 = 32'd112
; 
32'd9957: dataIn1 = 32'd124
; 
32'd9958: dataIn1 = 32'd10
; 
32'd9959: dataIn1 = 32'd11
; 
32'd9960: dataIn1 = 32'd96
; 
32'd9961: dataIn1 = 32'd12
; 
32'd9962: dataIn1 = 32'd107
; 
32'd9963: dataIn1 = 32'd126
; 
32'd9964: dataIn1 = 32'd139
; 
32'd9965: dataIn1 = 32'd153
; 
32'd9966: dataIn1 = 32'd13
; 
32'd9967: dataIn1 = 32'd86
; 
32'd9968: dataIn1 = 32'd96
; 
32'd9969: dataIn1 = 32'd126
; 
32'd9970: dataIn1 = 32'd14
; 
32'd9971: dataIn1 = 32'd120
; 
32'd9972: dataIn1 = 32'd15
; 
32'd9973: dataIn1 = 32'd120
; 
32'd9974: dataIn1 = 32'd127
; 
32'd9975: dataIn1 = 32'd16
; 
32'd9976: dataIn1 = 32'd120
; 
32'd9977: dataIn1 = 32'd159
; 
32'd9978: dataIn1 = 32'd17
; 
32'd9979: dataIn1 = 32'd94
; 
32'd9980: dataIn1 = 32'd127
; 
32'd9981: dataIn1 = 32'd18
; 
32'd9982: dataIn1 = 32'd94
; 
32'd9983: dataIn1 = 32'd19
; 
32'd9984: dataIn1 = 32'd94
; 
32'd9985: dataIn1 = 32'd20
; 
32'd9986: dataIn1 = 32'd102
; 
32'd9987: dataIn1 = 32'd114
; 
32'd9988: dataIn1 = 32'd21
; 
32'd9989: dataIn1 = 32'd102
; 
32'd9990: dataIn1 = 32'd140
; 
32'd9991: dataIn1 = 32'd22
; 
32'd9992: dataIn1 = 32'd83
; 
32'd9993: dataIn1 = 32'd99
; 
32'd9994: dataIn1 = 32'd102
; 
32'd9995: dataIn1 = 32'd23
; 
32'd9996: dataIn1 = 32'd99
; 
32'd9997: dataIn1 = 32'd24
; 
32'd9998: dataIn1 = 32'd99
; 
32'd9999: dataIn1 = 32'd25
; 
32'd10000: dataIn1 = 32'd26
; 
32'd10001: dataIn1 = 32'd115
; 
32'd10002: dataIn1 = 32'd140
; 
32'd10003: dataIn1 = 32'd142
; 
32'd10004: dataIn1 = 32'd154
; 
32'd10005: dataIn1 = 32'd164
; 
32'd10006: dataIn1 = 32'd27
; 
32'd10007: dataIn1 = 32'd128
; 
32'd10008: dataIn1 = 32'd140
; 
32'd10009: dataIn1 = 32'd142
; 
32'd10010: dataIn1 = 32'd28
; 
32'd10011: dataIn1 = 32'd115
; 
32'd10012: dataIn1 = 32'd29
; 
32'd10013: dataIn1 = 32'd116
; 
32'd10014: dataIn1 = 32'd144
; 
32'd10015: dataIn1 = 32'd156
; 
32'd10016: dataIn1 = 32'd166
; 
32'd10017: dataIn1 = 32'd195
; 
32'd10018: dataIn1 = 32'd30
; 
32'd10019: dataIn1 = 32'd115
; 
32'd10020: dataIn1 = 32'd144
; 
32'd10021: dataIn1 = 32'd31
; 
32'd10022: dataIn1 = 32'd129
; 
32'd10023: dataIn1 = 32'd144
; 
32'd10024: dataIn1 = 32'd32
; 
32'd10025: dataIn1 = 32'd106
; 
32'd10026: dataIn1 = 32'd118
; 
32'd10027: dataIn1 = 32'd130
; 
32'd10028: dataIn1 = 32'd167
; 
32'd10029: dataIn1 = 32'd33
; 
32'd10030: dataIn1 = 32'd106
; 
32'd10031: dataIn1 = 32'd34
; 
32'd10032: dataIn1 = 32'd84
; 
32'd10033: dataIn1 = 32'd106
; 
32'd10034: dataIn1 = 32'd35
; 
32'd10035: dataIn1 = 32'd84
; 
32'd10036: dataIn1 = 32'd95
; 
32'd10037: dataIn1 = 32'd36
; 
32'd10038: dataIn1 = 32'd95
; 
32'd10039: dataIn1 = 32'd103
; 
32'd10040: dataIn1 = 32'd37
; 
32'd10041: dataIn1 = 32'd95
; 
32'd10042: dataIn1 = 32'd38
; 
32'd10043: dataIn1 = 32'd92
; 
32'd10044: dataIn1 = 32'd129
; 
32'd10045: dataIn1 = 32'd39
; 
32'd10046: dataIn1 = 32'd40
; 
32'd10047: dataIn1 = 32'd104
; 
32'd10048: dataIn1 = 32'd113
; 
32'd10049: dataIn1 = 32'd117
; 
32'd10050: dataIn1 = 32'd129
; 
32'd10051: dataIn1 = 32'd155
; 
32'd10052: dataIn1 = 32'd157
; 
32'd10053: dataIn1 = 32'd160
; 
32'd10054: dataIn1 = 32'd168
; 
32'd10055: dataIn1 = 32'd41
; 
32'd10056: dataIn1 = 32'd92
; 
32'd10057: dataIn1 = 32'd105
; 
32'd10058: dataIn1 = 32'd42
; 
32'd10059: dataIn1 = 32'd93
; 
32'd10060: dataIn1 = 32'd104
; 
32'd10061: dataIn1 = 32'd43
; 
32'd10062: dataIn1 = 32'd105
; 
32'd10063: dataIn1 = 32'd44
; 
32'd10064: dataIn1 = 32'd45
; 
32'd10065: dataIn1 = 32'd93
; 
32'd10066: dataIn1 = 32'd109
; 
32'd10067: dataIn1 = 32'd131
; 
32'd10068: dataIn1 = 32'd46
; 
32'd10069: dataIn1 = 32'd93
; 
32'd10070: dataIn1 = 32'd131
; 
32'd10071: dataIn1 = 32'd47
; 
32'd10072: dataIn1 = 32'd48
; 
32'd10073: dataIn1 = 32'd103
; 
32'd10074: dataIn1 = 32'd132
; 
32'd10075: dataIn1 = 32'd49
; 
32'd10076: dataIn1 = 32'd103
; 
32'd10077: dataIn1 = 32'd108
; 
32'd10078: dataIn1 = 32'd133
; 
32'd10079: dataIn1 = 32'd50
; 
32'd10080: dataIn1 = 32'd109
; 
32'd10081: dataIn1 = 32'd133
; 
32'd10082: dataIn1 = 32'd51
; 
32'd10083: dataIn1 = 32'd108
; 
32'd10084: dataIn1 = 32'd52
; 
32'd10085: dataIn1 = 32'd112
; 
32'd10086: dataIn1 = 32'd162
; 
32'd10087: dataIn1 = 32'd169
; 
32'd10088: dataIn1 = 32'd181
; 
32'd10089: dataIn1 = 32'd53
; 
32'd10090: dataIn1 = 32'd108
; 
32'd10091: dataIn1 = 32'd54
; 
32'd10092: dataIn1 = 32'd55
; 
32'd10093: dataIn1 = 32'd101
; 
32'd10094: dataIn1 = 32'd111
; 
32'd10095: dataIn1 = 32'd112
; 
32'd10096: dataIn1 = 32'd56
; 
32'd10097: dataIn1 = 32'd83
; 
32'd10098: dataIn1 = 32'd57
; 
32'd10099: dataIn1 = 32'd85
; 
32'd10100: dataIn1 = 32'd101
; 
32'd10101: dataIn1 = 32'd111
; 
32'd10102: dataIn1 = 32'd58
; 
32'd10103: dataIn1 = 32'd96
; 
32'd10104: dataIn1 = 32'd59
; 
32'd10105: dataIn1 = 32'd86
; 
32'd10106: dataIn1 = 32'd109
; 
32'd10107: dataIn1 = 32'd60
; 
32'd10108: dataIn1 = 32'd86
; 
32'd10109: dataIn1 = 32'd110
; 
32'd10110: dataIn1 = 32'd61
; 
32'd10111: dataIn1 = 32'd92
; 
32'd10112: dataIn1 = 32'd110
; 
32'd10113: dataIn1 = 32'd62
; 
32'd10114: dataIn1 = 32'd100
; 
32'd10115: dataIn1 = 32'd132
; 
32'd10116: dataIn1 = 32'd134
; 
32'd10117: dataIn1 = 32'd63
; 
32'd10118: dataIn1 = 32'd132
; 
32'd10119: dataIn1 = 32'd64
; 
32'd10120: dataIn1 = 32'd104
; 
32'd10121: dataIn1 = 32'd65
; 
32'd10122: dataIn1 = 32'd100
; 
32'd10123: dataIn1 = 32'd66
; 
32'd10124: dataIn1 = 32'd128
; 
32'd10125: dataIn1 = 32'd67
; 
32'd10126: dataIn1 = 32'd110
; 
32'd10127: dataIn1 = 32'd127
; 
32'd10128: dataIn1 = 32'd68
; 
32'd10129: dataIn1 = 32'd116
; 
32'd10130: dataIn1 = 32'd69
; 
32'd10131: dataIn1 = 32'd83
; 
32'd10132: dataIn1 = 32'd114
; 
32'd10133: dataIn1 = 32'd119
; 
32'd10134: dataIn1 = 32'd70
; 
32'd10135: dataIn1 = 32'd114
; 
32'd10136: dataIn1 = 32'd135
; 
32'd10137: dataIn1 = 32'd159
; 
32'd10138: dataIn1 = 32'd170
; 
32'd10139: dataIn1 = 32'd179
; 
32'd10140: dataIn1 = 32'd189
; 
32'd10141: dataIn1 = 32'd213
; 
32'd10142: dataIn1 = 32'd71
; 
32'd10143: dataIn1 = 32'd135
; 
32'd10144: dataIn1 = 32'd72
; 
32'd10145: dataIn1 = 32'd135
; 
32'd10146: dataIn1 = 32'd73
; 
32'd10147: dataIn1 = 32'd74
; 
32'd10148: dataIn1 = 32'd136
; 
32'd10149: dataIn1 = 32'd75
; 
32'd10150: dataIn1 = 32'd118
; 
32'd10151: dataIn1 = 32'd76
; 
32'd10152: dataIn1 = 32'd118
; 
32'd10153: dataIn1 = 32'd137
; 
32'd10154: dataIn1 = 32'd77
; 
32'd10155: dataIn1 = 32'd137
; 
32'd10156: dataIn1 = 32'd78
; 
32'd10157: dataIn1 = 32'd117
; 
32'd10158: dataIn1 = 32'd137
; 
32'd10159: dataIn1 = 32'd145
; 
32'd10160: dataIn1 = 32'd148
; 
32'd10161: dataIn1 = 32'd79
; 
32'd10162: dataIn1 = 32'd97
; 
32'd10163: dataIn1 = 32'd80
; 
32'd10164: dataIn1 = 32'd113
; 
32'd10165: dataIn1 = 32'd117
; 
32'd10166: dataIn1 = 32'd145
; 
32'd10167: dataIn1 = 32'd146
; 
32'd10168: dataIn1 = 32'd188
; 
32'd10169: dataIn1 = 32'd81
; 
32'd10170: dataIn1 = 32'd97
; 
32'd10171: dataIn1 = 32'd125
; 
32'd10172: dataIn1 = 32'd82
; 
32'd10173: dataIn1 = 32'd113
; 
32'd10174: dataIn1 = 32'd125
; 
32'd10175: dataIn1 = 32'd141
; 
32'd10176: dataIn1 = 32'd146
; 
32'd10177: dataIn1 = 32'd171
; 
32'd10178: dataIn1 = 32'd83
; 
32'd10179: dataIn1 = 32'd119
; 
32'd10180: dataIn1 = 32'd169
; 
32'd10181: dataIn1 = 32'd182
; 
32'd10182: dataIn1 = 32'd196
; 
32'd10183: dataIn1 = 32'd84
; 
32'd10184: dataIn1 = 32'd172
; 
32'd10185: dataIn1 = 32'd183
; 
32'd10186: dataIn1 = 32'd191
; 
32'd10187: dataIn1 = 32'd85
; 
32'd10188: dataIn1 = 32'd147
; 
32'd10189: dataIn1 = 32'd152
; 
32'd10190: dataIn1 = 32'd173
; 
32'd10191: dataIn1 = 32'd214
; 
32'd10192: dataIn1 = 32'd86
; 
32'd10193: dataIn1 = 32'd121
; 
32'd10194: dataIn1 = 32'd161
; 
32'd10195: dataIn1 = 32'd174
; 
32'd10196: dataIn1 = 32'd198
; 
32'd10197: dataIn1 = 32'd87
; 
32'd10198: dataIn1 = 32'd100
; 
32'd10199: dataIn1 = 32'd160
; 
32'd10200: dataIn1 = 32'd83
; 
32'd10201: dataIn1 = 32'd88
; 
32'd10202: dataIn1 = 32'd119
; 
32'd10203: dataIn1 = 32'd89
; 
32'd10204: dataIn1 = 32'd165
; 
32'd10205: dataIn1 = 32'd175
; 
32'd10206: dataIn1 = 32'd90
; 
32'd10207: dataIn1 = 32'd130
; 
32'd10208: dataIn1 = 32'd91
; 
32'd10209: dataIn1 = 32'd97
; 
32'd10210: dataIn1 = 32'd139
; 
32'd10211: dataIn1 = 32'd159
; 
32'd10212: dataIn1 = 32'd176
; 
32'd10213: dataIn1 = 32'd92
; 
32'd10214: dataIn1 = 32'd105
; 
32'd10215: dataIn1 = 32'd116
; 
32'd10216: dataIn1 = 32'd155
; 
32'd10217: dataIn1 = 32'd156
; 
32'd10218: dataIn1 = 32'd177
; 
32'd10219: dataIn1 = 32'd93
; 
32'd10220: dataIn1 = 32'd134
; 
32'd10221: dataIn1 = 32'd178
; 
32'd10222: dataIn1 = 32'd94
; 
32'd10223: dataIn1 = 32'd128
; 
32'd10224: dataIn1 = 32'd179
; 
32'd10225: dataIn1 = 32'd194
; 
32'd10226: dataIn1 = 32'd221
; 
32'd10227: dataIn1 = 32'd95
; 
32'd10228: dataIn1 = 32'd180
; 
32'd10229: dataIn1 = 32'd190
; 
32'd10230: dataIn1 = 32'd96
; 
32'd10231: dataIn1 = 32'd126
; 
32'd10232: dataIn1 = 32'd174
; 
32'd10233: dataIn1 = 32'd181
; 
32'd10234: dataIn1 = 32'd184
; 
32'd10235: dataIn1 = 32'd97
; 
32'd10236: dataIn1 = 32'd145
; 
32'd10237: dataIn1 = 32'd153
; 
32'd10238: dataIn1 = 32'd176
; 
32'd10239: dataIn1 = 32'd204
; 
32'd10240: dataIn1 = 32'd98
; 
32'd10241: dataIn1 = 32'd123
; 
32'd10242: dataIn1 = 32'd141
; 
32'd10243: dataIn1 = 32'd99
; 
32'd10244: dataIn1 = 32'd154
; 
32'd10245: dataIn1 = 32'd185
; 
32'd10246: dataIn1 = 32'd196
; 
32'd10247: dataIn1 = 32'd100
; 
32'd10248: dataIn1 = 32'd151
; 
32'd10249: dataIn1 = 32'd171
; 
32'd10250: dataIn1 = 32'd222
; 
32'd10251: dataIn1 = 32'd101
; 
32'd10252: dataIn1 = 32'd111
; 
32'd10253: dataIn1 = 32'd173
; 
32'd10254: dataIn1 = 32'd187
; 
32'd10255: dataIn1 = 32'd102
; 
32'd10256: dataIn1 = 32'd182
; 
32'd10257: dataIn1 = 32'd210
; 
32'd10258: dataIn1 = 32'd265
; 
32'd10259: dataIn1 = 32'd103
; 
32'd10260: dataIn1 = 32'd149
; 
32'd10261: dataIn1 = 32'd158
; 
32'd10262: dataIn1 = 32'd164
; 
32'd10263: dataIn1 = 32'd180
; 
32'd10264: dataIn1 = 32'd199
; 
32'd10265: dataIn1 = 32'd215
; 
32'd10266: dataIn1 = 32'd104
; 
32'd10267: dataIn1 = 32'd134
; 
32'd10268: dataIn1 = 32'd160
; 
32'd10269: dataIn1 = 32'd163
; 
32'd10270: dataIn1 = 32'd201
; 
32'd10271: dataIn1 = 32'd92
; 
32'd10272: dataIn1 = 32'd105
; 
32'd10273: dataIn1 = 32'd121
; 
32'd10274: dataIn1 = 32'd155
; 
32'd10275: dataIn1 = 32'd163
; 
32'd10276: dataIn1 = 32'd177
; 
32'd10277: dataIn1 = 32'd106
; 
32'd10278: dataIn1 = 32'd130
; 
32'd10279: dataIn1 = 32'd150
; 
32'd10280: dataIn1 = 32'd183
; 
32'd10281: dataIn1 = 32'd107
; 
32'd10282: dataIn1 = 32'd184
; 
32'd10283: dataIn1 = 32'd193
; 
32'd10284: dataIn1 = 32'd108
; 
32'd10285: dataIn1 = 32'd158
; 
32'd10286: dataIn1 = 32'd185
; 
32'd10287: dataIn1 = 32'd109
; 
32'd10288: dataIn1 = 32'd121
; 
32'd10289: dataIn1 = 32'd131
; 
32'd10290: dataIn1 = 32'd162
; 
32'd10291: dataIn1 = 32'd174
; 
32'd10292: dataIn1 = 32'd178
; 
32'd10293: dataIn1 = 32'd223
; 
32'd10294: dataIn1 = 32'd110
; 
32'd10295: dataIn1 = 32'd177
; 
32'd10296: dataIn1 = 32'd101
; 
32'd10297: dataIn1 = 32'd111
; 
32'd10298: dataIn1 = 32'd173
; 
32'd10299: dataIn1 = 32'd186
; 
32'd10300: dataIn1 = 32'd112
; 
32'd10301: dataIn1 = 32'd169
; 
32'd10302: dataIn1 = 32'd181
; 
32'd10303: dataIn1 = 32'd184
; 
32'd10304: dataIn1 = 32'd187
; 
32'd10305: dataIn1 = 32'd224
; 
32'd10306: dataIn1 = 32'd248
; 
32'd10307: dataIn1 = 32'd113
; 
32'd10308: dataIn1 = 32'd146
; 
32'd10309: dataIn1 = 32'd168
; 
32'd10310: dataIn1 = 32'd171
; 
32'd10311: dataIn1 = 32'd188
; 
32'd10312: dataIn1 = 32'd114
; 
32'd10313: dataIn1 = 32'd179
; 
32'd10314: dataIn1 = 32'd182
; 
32'd10315: dataIn1 = 32'd189
; 
32'd10316: dataIn1 = 32'd115
; 
32'd10317: dataIn1 = 32'd142
; 
32'd10318: dataIn1 = 32'd150
; 
32'd10319: dataIn1 = 32'd190
; 
32'd10320: dataIn1 = 32'd92
; 
32'd10321: dataIn1 = 32'd116
; 
32'd10322: dataIn1 = 32'd143
; 
32'd10323: dataIn1 = 32'd117
; 
32'd10324: dataIn1 = 32'd148
; 
32'd10325: dataIn1 = 32'd188
; 
32'd10326: dataIn1 = 32'd208
; 
32'd10327: dataIn1 = 32'd118
; 
32'd10328: dataIn1 = 32'd136
; 
32'd10329: dataIn1 = 32'd148
; 
32'd10330: dataIn1 = 32'd170
; 
32'd10331: dataIn1 = 32'd225
; 
32'd10332: dataIn1 = 32'd83
; 
32'd10333: dataIn1 = 32'd119
; 
32'd10334: dataIn1 = 32'd152
; 
32'd10335: dataIn1 = 32'd189
; 
32'd10336: dataIn1 = 32'd226
; 
32'd10337: dataIn1 = 32'd120
; 
32'd10338: dataIn1 = 32'd139
; 
32'd10339: dataIn1 = 32'd161
; 
32'd10340: dataIn1 = 32'd227
; 
32'd10341: dataIn1 = 32'd86
; 
32'd10342: dataIn1 = 32'd105
; 
32'd10343: dataIn1 = 32'd109
; 
32'd10344: dataIn1 = 32'd121
; 
32'd10345: dataIn1 = 32'd198
; 
32'd10346: dataIn1 = 32'd200
; 
32'd10347: dataIn1 = 32'd122
; 
32'd10348: dataIn1 = 32'd151
; 
32'd10349: dataIn1 = 32'd172
; 
32'd10350: dataIn1 = 32'd191
; 
32'd10351: dataIn1 = 32'd192
; 
32'd10352: dataIn1 = 32'd228
; 
32'd10353: dataIn1 = 32'd123
; 
32'd10354: dataIn1 = 32'd147
; 
32'd10355: dataIn1 = 32'd187
; 
32'd10356: dataIn1 = 32'd192
; 
32'd10357: dataIn1 = 32'd211
; 
32'd10358: dataIn1 = 32'd220
; 
32'd10359: dataIn1 = 32'd228
; 
32'd10360: dataIn1 = 32'd124
; 
32'd10361: dataIn1 = 32'd193
; 
32'd10362: dataIn1 = 32'd125
; 
32'd10363: dataIn1 = 32'd153
; 
32'd10364: dataIn1 = 32'd193
; 
32'd10365: dataIn1 = 32'd204
; 
32'd10366: dataIn1 = 32'd220
; 
32'd10367: dataIn1 = 32'd229
; 
32'd10368: dataIn1 = 32'd96
; 
32'd10369: dataIn1 = 32'd126
; 
32'd10370: dataIn1 = 32'd197
; 
32'd10371: dataIn1 = 32'd218
; 
32'd10372: dataIn1 = 32'd230
; 
32'd10373: dataIn1 = 32'd127
; 
32'd10374: dataIn1 = 32'd143
; 
32'd10375: dataIn1 = 32'd161
; 
32'd10376: dataIn1 = 32'd194
; 
32'd10377: dataIn1 = 32'd94
; 
32'd10378: dataIn1 = 32'd128
; 
32'd10379: dataIn1 = 32'd143
; 
32'd10380: dataIn1 = 32'd195
; 
32'd10381: dataIn1 = 32'd210
; 
32'd10382: dataIn1 = 32'd219
; 
32'd10383: dataIn1 = 32'd221
; 
32'd10384: dataIn1 = 32'd231
; 
32'd10385: dataIn1 = 32'd129
; 
32'd10386: dataIn1 = 32'd156
; 
32'd10387: dataIn1 = 32'd157
; 
32'd10388: dataIn1 = 32'd209
; 
32'd10389: dataIn1 = 32'd212
; 
32'd10390: dataIn1 = 32'd106
; 
32'd10391: dataIn1 = 32'd130
; 
32'd10392: dataIn1 = 32'd167
; 
32'd10393: dataIn1 = 32'd175
; 
32'd10394: dataIn1 = 32'd225
; 
32'd10395: dataIn1 = 32'd232
; 
32'd10396: dataIn1 = 32'd109
; 
32'd10397: dataIn1 = 32'd131
; 
32'd10398: dataIn1 = 32'd133
; 
32'd10399: dataIn1 = 32'd149
; 
32'd10400: dataIn1 = 32'd178
; 
32'd10401: dataIn1 = 32'd233
; 
32'd10402: dataIn1 = 32'd132
; 
32'd10403: dataIn1 = 32'd172
; 
32'd10404: dataIn1 = 32'd216
; 
32'd10405: dataIn1 = 32'd233
; 
32'd10406: dataIn1 = 32'd234
; 
32'd10407: dataIn1 = 32'd131
; 
32'd10408: dataIn1 = 32'd133
; 
32'd10409: dataIn1 = 32'd149
; 
32'd10410: dataIn1 = 32'd162
; 
32'd10411: dataIn1 = 32'd93
; 
32'd10412: dataIn1 = 32'd104
; 
32'd10413: dataIn1 = 32'd134
; 
32'd10414: dataIn1 = 32'd201
; 
32'd10415: dataIn1 = 32'd222
; 
32'd10416: dataIn1 = 32'd235
; 
32'd10417: dataIn1 = 32'd135
; 
32'd10418: dataIn1 = 32'd136
; 
32'd10419: dataIn1 = 32'd152
; 
32'd10420: dataIn1 = 32'd236
; 
32'd10421: dataIn1 = 32'd118
; 
32'd10422: dataIn1 = 32'd135
; 
32'd10423: dataIn1 = 32'd136
; 
32'd10424: dataIn1 = 32'd170
; 
32'd10425: dataIn1 = 32'd175
; 
32'd10426: dataIn1 = 32'd236
; 
32'd10427: dataIn1 = 32'd137
; 
32'd10428: dataIn1 = 32'd176
; 
32'd10429: dataIn1 = 32'd213
; 
32'd10430: dataIn1 = 32'd122
; 
32'd10431: dataIn1 = 32'd138
; 
32'd10432: dataIn1 = 32'd151
; 
32'd10433: dataIn1 = 32'd120
; 
32'd10434: dataIn1 = 32'd139
; 
32'd10435: dataIn1 = 32'd197
; 
32'd10436: dataIn1 = 32'd140
; 
32'd10437: dataIn1 = 32'd154
; 
32'd10438: dataIn1 = 32'd141
; 
32'd10439: dataIn1 = 32'd192
; 
32'd10440: dataIn1 = 32'd115
; 
32'd10441: dataIn1 = 32'd142
; 
32'd10442: dataIn1 = 32'd166
; 
32'd10443: dataIn1 = 32'd219
; 
32'd10444: dataIn1 = 32'd116
; 
32'd10445: dataIn1 = 32'd127
; 
32'd10446: dataIn1 = 32'd128
; 
32'd10447: dataIn1 = 32'd143
; 
32'd10448: dataIn1 = 32'd195
; 
32'd10449: dataIn1 = 32'd207
; 
32'd10450: dataIn1 = 32'd284
; 
32'd10451: dataIn1 = 32'd144
; 
32'd10452: dataIn1 = 32'd150
; 
32'd10453: dataIn1 = 32'd166
; 
32'd10454: dataIn1 = 32'd202
; 
32'd10455: dataIn1 = 32'd212
; 
32'd10456: dataIn1 = 32'd97
; 
32'd10457: dataIn1 = 32'd145
; 
32'd10458: dataIn1 = 32'd208
; 
32'd10459: dataIn1 = 32'd237
; 
32'd10460: dataIn1 = 32'd113
; 
32'd10461: dataIn1 = 32'd146
; 
32'd10462: dataIn1 = 32'd204
; 
32'd10463: dataIn1 = 32'd85
; 
32'd10464: dataIn1 = 32'd123
; 
32'd10465: dataIn1 = 32'd147
; 
32'd10466: dataIn1 = 32'd165
; 
32'd10467: dataIn1 = 32'd228
; 
32'd10468: dataIn1 = 32'd117
; 
32'd10469: dataIn1 = 32'd118
; 
32'd10470: dataIn1 = 32'd148
; 
32'd10471: dataIn1 = 32'd237
; 
32'd10472: dataIn1 = 32'd238
; 
32'd10473: dataIn1 = 32'd245
; 
32'd10474: dataIn1 = 32'd266
; 
32'd10475: dataIn1 = 32'd103
; 
32'd10476: dataIn1 = 32'd131
; 
32'd10477: dataIn1 = 32'd133
; 
32'd10478: dataIn1 = 32'd149
; 
32'd10479: dataIn1 = 32'd158
; 
32'd10480: dataIn1 = 32'd239
; 
32'd10481: dataIn1 = 32'd106
; 
32'd10482: dataIn1 = 32'd115
; 
32'd10483: dataIn1 = 32'd144
; 
32'd10484: dataIn1 = 32'd150
; 
32'd10485: dataIn1 = 32'd167
; 
32'd10486: dataIn1 = 32'd100
; 
32'd10487: dataIn1 = 32'd122
; 
32'd10488: dataIn1 = 32'd151
; 
32'd10489: dataIn1 = 32'd216
; 
32'd10490: dataIn1 = 32'd85
; 
32'd10491: dataIn1 = 32'd119
; 
32'd10492: dataIn1 = 32'd135
; 
32'd10493: dataIn1 = 32'd152
; 
32'd10494: dataIn1 = 32'd186
; 
32'd10495: dataIn1 = 32'd214
; 
32'd10496: dataIn1 = 32'd226
; 
32'd10497: dataIn1 = 32'd267
; 
32'd10498: dataIn1 = 32'd97
; 
32'd10499: dataIn1 = 32'd125
; 
32'd10500: dataIn1 = 32'd153
; 
32'd10501: dataIn1 = 32'd197
; 
32'd10502: dataIn1 = 32'd99
; 
32'd10503: dataIn1 = 32'd140
; 
32'd10504: dataIn1 = 32'd154
; 
32'd10505: dataIn1 = 32'd164
; 
32'd10506: dataIn1 = 32'd206
; 
32'd10507: dataIn1 = 32'd210
; 
32'd10508: dataIn1 = 32'd252
; 
32'd10509: dataIn1 = 32'd268
; 
32'd10510: dataIn1 = 32'd92
; 
32'd10511: dataIn1 = 32'd105
; 
32'd10512: dataIn1 = 32'd155
; 
32'd10513: dataIn1 = 32'd157
; 
32'd10514: dataIn1 = 32'd163
; 
32'd10515: dataIn1 = 32'd92
; 
32'd10516: dataIn1 = 32'd129
; 
32'd10517: dataIn1 = 32'd156
; 
32'd10518: dataIn1 = 32'd205
; 
32'd10519: dataIn1 = 32'd212
; 
32'd10520: dataIn1 = 32'd240
; 
32'd10521: dataIn1 = 32'd257
; 
32'd10522: dataIn1 = 32'd264
; 
32'd10523: dataIn1 = 32'd274
; 
32'd10524: dataIn1 = 32'd129
; 
32'd10525: dataIn1 = 32'd155
; 
32'd10526: dataIn1 = 32'd157
; 
32'd10527: dataIn1 = 32'd209
; 
32'd10528: dataIn1 = 32'd251
; 
32'd10529: dataIn1 = 32'd257
; 
32'd10530: dataIn1 = 32'd258
; 
32'd10531: dataIn1 = 32'd103
; 
32'd10532: dataIn1 = 32'd108
; 
32'd10533: dataIn1 = 32'd149
; 
32'd10534: dataIn1 = 32'd158
; 
32'd10535: dataIn1 = 32'd185
; 
32'd10536: dataIn1 = 32'd159
; 
32'd10537: dataIn1 = 32'd253
; 
32'd10538: dataIn1 = 32'd269
; 
32'd10539: dataIn1 = 32'd104
; 
32'd10540: dataIn1 = 32'd160
; 
32'd10541: dataIn1 = 32'd168
; 
32'd10542: dataIn1 = 32'd251
; 
32'd10543: dataIn1 = 32'd86
; 
32'd10544: dataIn1 = 32'd120
; 
32'd10545: dataIn1 = 32'd127
; 
32'd10546: dataIn1 = 32'd161
; 
32'd10547: dataIn1 = 32'd194
; 
32'd10548: dataIn1 = 32'd207
; 
32'd10549: dataIn1 = 32'd218
; 
32'd10550: dataIn1 = 32'd243
; 
32'd10551: dataIn1 = 32'd109
; 
32'd10552: dataIn1 = 32'd133
; 
32'd10553: dataIn1 = 32'd162
; 
32'd10554: dataIn1 = 32'd223
; 
32'd10555: dataIn1 = 32'd242
; 
32'd10556: dataIn1 = 32'd246
; 
32'd10557: dataIn1 = 32'd270
; 
32'd10558: dataIn1 = 32'd104
; 
32'd10559: dataIn1 = 32'd105
; 
32'd10560: dataIn1 = 32'd155
; 
32'd10561: dataIn1 = 32'd163
; 
32'd10562: dataIn1 = 32'd201
; 
32'd10563: dataIn1 = 32'd103
; 
32'd10564: dataIn1 = 32'd154
; 
32'd10565: dataIn1 = 32'd164
; 
32'd10566: dataIn1 = 32'd180
; 
32'd10567: dataIn1 = 32'd190
; 
32'd10568: dataIn1 = 32'd199
; 
32'd10569: dataIn1 = 32'd215
; 
32'd10570: dataIn1 = 32'd252
; 
32'd10571: dataIn1 = 32'd147
; 
32'd10572: dataIn1 = 32'd165
; 
32'd10573: dataIn1 = 32'd191
; 
32'd10574: dataIn1 = 32'd214
; 
32'd10575: dataIn1 = 32'd142
; 
32'd10576: dataIn1 = 32'd144
; 
32'd10577: dataIn1 = 32'd166
; 
32'd10578: dataIn1 = 32'd219
; 
32'd10579: dataIn1 = 32'd240
; 
32'd10580: dataIn1 = 32'd241
; 
32'd10581: dataIn1 = 32'd130
; 
32'd10582: dataIn1 = 32'd150
; 
32'd10583: dataIn1 = 32'd167
; 
32'd10584: dataIn1 = 32'd202
; 
32'd10585: dataIn1 = 32'd238
; 
32'd10586: dataIn1 = 32'd259
; 
32'd10587: dataIn1 = 32'd271
; 
32'd10588: dataIn1 = 32'd289
; 
32'd10589: dataIn1 = 32'd113
; 
32'd10590: dataIn1 = 32'd160
; 
32'd10591: dataIn1 = 32'd168
; 
32'd10592: dataIn1 = 32'd209
; 
32'd10593: dataIn1 = 32'd217
; 
32'd10594: dataIn1 = 32'd83
; 
32'd10595: dataIn1 = 32'd112
; 
32'd10596: dataIn1 = 32'd169
; 
32'd10597: dataIn1 = 32'd203
; 
32'd10598: dataIn1 = 32'd248
; 
32'd10599: dataIn1 = 32'd270
; 
32'd10600: dataIn1 = 32'd272
; 
32'd10601: dataIn1 = 32'd118
; 
32'd10602: dataIn1 = 32'd136
; 
32'd10603: dataIn1 = 32'd170
; 
32'd10604: dataIn1 = 32'd213
; 
32'd10605: dataIn1 = 32'd100
; 
32'd10606: dataIn1 = 32'd113
; 
32'd10607: dataIn1 = 32'd171
; 
32'd10608: dataIn1 = 32'd217
; 
32'd10609: dataIn1 = 32'd260
; 
32'd10610: dataIn1 = 32'd263
; 
32'd10611: dataIn1 = 32'd84
; 
32'd10612: dataIn1 = 32'd122
; 
32'd10613: dataIn1 = 32'd132
; 
32'd10614: dataIn1 = 32'd172
; 
32'd10615: dataIn1 = 32'd216
; 
32'd10616: dataIn1 = 32'd85
; 
32'd10617: dataIn1 = 32'd101
; 
32'd10618: dataIn1 = 32'd111
; 
32'd10619: dataIn1 = 32'd173
; 
32'd10620: dataIn1 = 32'd186
; 
32'd10621: dataIn1 = 32'd203
; 
32'd10622: dataIn1 = 32'd211
; 
32'd10623: dataIn1 = 32'd86
; 
32'd10624: dataIn1 = 32'd96
; 
32'd10625: dataIn1 = 32'd109
; 
32'd10626: dataIn1 = 32'd174
; 
32'd10627: dataIn1 = 32'd198
; 
32'd10628: dataIn1 = 32'd218
; 
32'd10629: dataIn1 = 32'd242
; 
32'd10630: dataIn1 = 32'd130
; 
32'd10631: dataIn1 = 32'd136
; 
32'd10632: dataIn1 = 32'd175
; 
32'd10633: dataIn1 = 32'd225
; 
32'd10634: dataIn1 = 32'd232
; 
32'd10635: dataIn1 = 32'd273
; 
32'd10636: dataIn1 = 32'd97
; 
32'd10637: dataIn1 = 32'd137
; 
32'd10638: dataIn1 = 32'd176
; 
32'd10639: dataIn1 = 32'd237
; 
32'd10640: dataIn1 = 32'd253
; 
32'd10641: dataIn1 = 32'd92
; 
32'd10642: dataIn1 = 32'd105
; 
32'd10643: dataIn1 = 32'd110
; 
32'd10644: dataIn1 = 32'd177
; 
32'd10645: dataIn1 = 32'd200
; 
32'd10646: dataIn1 = 32'd205
; 
32'd10647: dataIn1 = 32'd207
; 
32'd10648: dataIn1 = 32'd264
; 
32'd10649: dataIn1 = 32'd274
; 
32'd10650: dataIn1 = 32'd298
; 
32'd10651: dataIn1 = 32'd311
; 
32'd10652: dataIn1 = 32'd93
; 
32'd10653: dataIn1 = 32'd109
; 
32'd10654: dataIn1 = 32'd131
; 
32'd10655: dataIn1 = 32'd178
; 
32'd10656: dataIn1 = 32'd200
; 
32'd10657: dataIn1 = 32'd223
; 
32'd10658: dataIn1 = 32'd94
; 
32'd10659: dataIn1 = 32'd114
; 
32'd10660: dataIn1 = 32'd179
; 
32'd10661: dataIn1 = 32'd265
; 
32'd10662: dataIn1 = 32'd269
; 
32'd10663: dataIn1 = 32'd275
; 
32'd10664: dataIn1 = 32'd286
; 
32'd10665: dataIn1 = 32'd95
; 
32'd10666: dataIn1 = 32'd103
; 
32'd10667: dataIn1 = 32'd164
; 
32'd10668: dataIn1 = 32'd180
; 
32'd10669: dataIn1 = 32'd183
; 
32'd10670: dataIn1 = 32'd199
; 
32'd10671: dataIn1 = 32'd96
; 
32'd10672: dataIn1 = 32'd112
; 
32'd10673: dataIn1 = 32'd181
; 
32'd10674: dataIn1 = 32'd224
; 
32'd10675: dataIn1 = 32'd242
; 
32'd10676: dataIn1 = 32'd83
; 
32'd10677: dataIn1 = 32'd102
; 
32'd10678: dataIn1 = 32'd114
; 
32'd10679: dataIn1 = 32'd182
; 
32'd10680: dataIn1 = 32'd196
; 
32'd10681: dataIn1 = 32'd262
; 
32'd10682: dataIn1 = 32'd265
; 
32'd10683: dataIn1 = 32'd276
; 
32'd10684: dataIn1 = 32'd84
; 
32'd10685: dataIn1 = 32'd106
; 
32'd10686: dataIn1 = 32'd180
; 
32'd10687: dataIn1 = 32'd183
; 
32'd10688: dataIn1 = 32'd234
; 
32'd10689: dataIn1 = 32'd250
; 
32'd10690: dataIn1 = 32'd277
; 
32'd10691: dataIn1 = 32'd96
; 
32'd10692: dataIn1 = 32'd107
; 
32'd10693: dataIn1 = 32'd112
; 
32'd10694: dataIn1 = 32'd184
; 
32'd10695: dataIn1 = 32'd224
; 
32'd10696: dataIn1 = 32'd230
; 
32'd10697: dataIn1 = 32'd99
; 
32'd10698: dataIn1 = 32'd108
; 
32'd10699: dataIn1 = 32'd158
; 
32'd10700: dataIn1 = 32'd185
; 
32'd10701: dataIn1 = 32'd206
; 
32'd10702: dataIn1 = 32'd111
; 
32'd10703: dataIn1 = 32'd152
; 
32'd10704: dataIn1 = 32'd173
; 
32'd10705: dataIn1 = 32'd186
; 
32'd10706: dataIn1 = 32'd203
; 
32'd10707: dataIn1 = 32'd101
; 
32'd10708: dataIn1 = 32'd112
; 
32'd10709: dataIn1 = 32'd123
; 
32'd10710: dataIn1 = 32'd187
; 
32'd10711: dataIn1 = 32'd211
; 
32'd10712: dataIn1 = 32'd113
; 
32'd10713: dataIn1 = 32'd117
; 
32'd10714: dataIn1 = 32'd188
; 
32'd10715: dataIn1 = 32'd208
; 
32'd10716: dataIn1 = 32'd217
; 
32'd10717: dataIn1 = 32'd114
; 
32'd10718: dataIn1 = 32'd119
; 
32'd10719: dataIn1 = 32'd189
; 
32'd10720: dataIn1 = 32'd226
; 
32'd10721: dataIn1 = 32'd261
; 
32'd10722: dataIn1 = 32'd95
; 
32'd10723: dataIn1 = 32'd115
; 
32'd10724: dataIn1 = 32'd164
; 
32'd10725: dataIn1 = 32'd190
; 
32'd10726: dataIn1 = 32'd202
; 
32'd10727: dataIn1 = 32'd250
; 
32'd10728: dataIn1 = 32'd84
; 
32'd10729: dataIn1 = 32'd122
; 
32'd10730: dataIn1 = 32'd165
; 
32'd10731: dataIn1 = 32'd191
; 
32'd10732: dataIn1 = 32'd255
; 
32'd10733: dataIn1 = 32'd278
; 
32'd10734: dataIn1 = 32'd122
; 
32'd10735: dataIn1 = 32'd123
; 
32'd10736: dataIn1 = 32'd141
; 
32'd10737: dataIn1 = 32'd192
; 
32'd10738: dataIn1 = 32'd220
; 
32'd10739: dataIn1 = 32'd279
; 
32'd10740: dataIn1 = 32'd107
; 
32'd10741: dataIn1 = 32'd124
; 
32'd10742: dataIn1 = 32'd125
; 
32'd10743: dataIn1 = 32'd193
; 
32'd10744: dataIn1 = 32'd229
; 
32'd10745: dataIn1 = 32'd244
; 
32'd10746: dataIn1 = 32'd94
; 
32'd10747: dataIn1 = 32'd127
; 
32'd10748: dataIn1 = 32'd161
; 
32'd10749: dataIn1 = 32'd194
; 
32'd10750: dataIn1 = 32'd221
; 
32'd10751: dataIn1 = 32'd243
; 
32'd10752: dataIn1 = 32'd128
; 
32'd10753: dataIn1 = 32'd143
; 
32'd10754: dataIn1 = 32'd195
; 
32'd10755: dataIn1 = 32'd205
; 
32'd10756: dataIn1 = 32'd231
; 
32'd10757: dataIn1 = 32'd83
; 
32'd10758: dataIn1 = 32'd99
; 
32'd10759: dataIn1 = 32'd182
; 
32'd10760: dataIn1 = 32'd196
; 
32'd10761: dataIn1 = 32'd206
; 
32'd10762: dataIn1 = 32'd276
; 
32'd10763: dataIn1 = 32'd126
; 
32'd10764: dataIn1 = 32'd139
; 
32'd10765: dataIn1 = 32'd153
; 
32'd10766: dataIn1 = 32'd197
; 
32'd10767: dataIn1 = 32'd227
; 
32'd10768: dataIn1 = 32'd229
; 
32'd10769: dataIn1 = 32'd253
; 
32'd10770: dataIn1 = 32'd256
; 
32'd10771: dataIn1 = 32'd280
; 
32'd10772: dataIn1 = 32'd86
; 
32'd10773: dataIn1 = 32'd121
; 
32'd10774: dataIn1 = 32'd174
; 
32'd10775: dataIn1 = 32'd198
; 
32'd10776: dataIn1 = 32'd249
; 
32'd10777: dataIn1 = 32'd281
; 
32'd10778: dataIn1 = 32'd312
; 
32'd10779: dataIn1 = 32'd327
; 
32'd10780: dataIn1 = 32'd103
; 
32'd10781: dataIn1 = 32'd164
; 
32'd10782: dataIn1 = 32'd180
; 
32'd10783: dataIn1 = 32'd199
; 
32'd10784: dataIn1 = 32'd215
; 
32'd10785: dataIn1 = 32'd234
; 
32'd10786: dataIn1 = 32'd282
; 
32'd10787: dataIn1 = 32'd295
; 
32'd10788: dataIn1 = 32'd303
; 
32'd10789: dataIn1 = 32'd121
; 
32'd10790: dataIn1 = 32'd177
; 
32'd10791: dataIn1 = 32'd178
; 
32'd10792: dataIn1 = 32'd200
; 
32'd10793: dataIn1 = 32'd235
; 
32'd10794: dataIn1 = 32'd249
; 
32'd10795: dataIn1 = 32'd311
; 
32'd10796: dataIn1 = 32'd104
; 
32'd10797: dataIn1 = 32'd134
; 
32'd10798: dataIn1 = 32'd163
; 
32'd10799: dataIn1 = 32'd201
; 
32'd10800: dataIn1 = 32'd235
; 
32'd10801: dataIn1 = 32'd144
; 
32'd10802: dataIn1 = 32'd167
; 
32'd10803: dataIn1 = 32'd190
; 
32'd10804: dataIn1 = 32'd202
; 
32'd10805: dataIn1 = 32'd250
; 
32'd10806: dataIn1 = 32'd259
; 
32'd10807: dataIn1 = 32'd271
; 
32'd10808: dataIn1 = 32'd301
; 
32'd10809: dataIn1 = 32'd304
; 
32'd10810: dataIn1 = 32'd332
; 
32'd10811: dataIn1 = 32'd169
; 
32'd10812: dataIn1 = 32'd173
; 
32'd10813: dataIn1 = 32'd186
; 
32'd10814: dataIn1 = 32'd203
; 
32'd10815: dataIn1 = 32'd248
; 
32'd10816: dataIn1 = 32'd262
; 
32'd10817: dataIn1 = 32'd305
; 
32'd10818: dataIn1 = 32'd334
; 
32'd10819: dataIn1 = 32'd97
; 
32'd10820: dataIn1 = 32'd125
; 
32'd10821: dataIn1 = 32'd146
; 
32'd10822: dataIn1 = 32'd204
; 
32'd10823: dataIn1 = 32'd260
; 
32'd10824: dataIn1 = 32'd280
; 
32'd10825: dataIn1 = 32'd283
; 
32'd10826: dataIn1 = 32'd156
; 
32'd10827: dataIn1 = 32'd177
; 
32'd10828: dataIn1 = 32'd195
; 
32'd10829: dataIn1 = 32'd205
; 
32'd10830: dataIn1 = 32'd240
; 
32'd10831: dataIn1 = 32'd284
; 
32'd10832: dataIn1 = 32'd154
; 
32'd10833: dataIn1 = 32'd185
; 
32'd10834: dataIn1 = 32'd196
; 
32'd10835: dataIn1 = 32'd206
; 
32'd10836: dataIn1 = 32'd239
; 
32'd10837: dataIn1 = 32'd268
; 
32'd10838: dataIn1 = 32'd272
; 
32'd10839: dataIn1 = 32'd295
; 
32'd10840: dataIn1 = 32'd308
; 
32'd10841: dataIn1 = 32'd143
; 
32'd10842: dataIn1 = 32'd161
; 
32'd10843: dataIn1 = 32'd177
; 
32'd10844: dataIn1 = 32'd207
; 
32'd10845: dataIn1 = 32'd281
; 
32'd10846: dataIn1 = 32'd298
; 
32'd10847: dataIn1 = 32'd117
; 
32'd10848: dataIn1 = 32'd145
; 
32'd10849: dataIn1 = 32'd188
; 
32'd10850: dataIn1 = 32'd208
; 
32'd10851: dataIn1 = 32'd258
; 
32'd10852: dataIn1 = 32'd283
; 
32'd10853: dataIn1 = 32'd129
; 
32'd10854: dataIn1 = 32'd157
; 
32'd10855: dataIn1 = 32'd168
; 
32'd10856: dataIn1 = 32'd209
; 
32'd10857: dataIn1 = 32'd102
; 
32'd10858: dataIn1 = 32'd128
; 
32'd10859: dataIn1 = 32'd154
; 
32'd10860: dataIn1 = 32'd210
; 
32'd10861: dataIn1 = 32'd268
; 
32'd10862: dataIn1 = 32'd123
; 
32'd10863: dataIn1 = 32'd173
; 
32'd10864: dataIn1 = 32'd187
; 
32'd10865: dataIn1 = 32'd211
; 
32'd10866: dataIn1 = 32'd285
; 
32'd10867: dataIn1 = 32'd290
; 
32'd10868: dataIn1 = 32'd309
; 
32'd10869: dataIn1 = 32'd129
; 
32'd10870: dataIn1 = 32'd144
; 
32'd10871: dataIn1 = 32'd156
; 
32'd10872: dataIn1 = 32'd212
; 
32'd10873: dataIn1 = 32'd257
; 
32'd10874: dataIn1 = 32'd271
; 
32'd10875: dataIn1 = 32'd137
; 
32'd10876: dataIn1 = 32'd170
; 
32'd10877: dataIn1 = 32'd213
; 
32'd10878: dataIn1 = 32'd245
; 
32'd10879: dataIn1 = 32'd286
; 
32'd10880: dataIn1 = 32'd294
; 
32'd10881: dataIn1 = 32'd299
; 
32'd10882: dataIn1 = 32'd313
; 
32'd10883: dataIn1 = 32'd85
; 
32'd10884: dataIn1 = 32'd152
; 
32'd10885: dataIn1 = 32'd165
; 
32'd10886: dataIn1 = 32'd214
; 
32'd10887: dataIn1 = 32'd255
; 
32'd10888: dataIn1 = 32'd267
; 
32'd10889: dataIn1 = 32'd103
; 
32'd10890: dataIn1 = 32'd164
; 
32'd10891: dataIn1 = 32'd199
; 
32'd10892: dataIn1 = 32'd215
; 
32'd10893: dataIn1 = 32'd239
; 
32'd10894: dataIn1 = 32'd132
; 
32'd10895: dataIn1 = 32'd151
; 
32'd10896: dataIn1 = 32'd172
; 
32'd10897: dataIn1 = 32'd216
; 
32'd10898: dataIn1 = 32'd222
; 
32'd10899: dataIn1 = 32'd287
; 
32'd10900: dataIn1 = 32'd168
; 
32'd10901: dataIn1 = 32'd171
; 
32'd10902: dataIn1 = 32'd188
; 
32'd10903: dataIn1 = 32'd217
; 
32'd10904: dataIn1 = 32'd258
; 
32'd10905: dataIn1 = 32'd126
; 
32'd10906: dataIn1 = 32'd161
; 
32'd10907: dataIn1 = 32'd174
; 
32'd10908: dataIn1 = 32'd218
; 
32'd10909: dataIn1 = 32'd227
; 
32'd10910: dataIn1 = 32'd247
; 
32'd10911: dataIn1 = 32'd281
; 
32'd10912: dataIn1 = 32'd314
; 
32'd10913: dataIn1 = 32'd128
; 
32'd10914: dataIn1 = 32'd142
; 
32'd10915: dataIn1 = 32'd166
; 
32'd10916: dataIn1 = 32'd219
; 
32'd10917: dataIn1 = 32'd231
; 
32'd10918: dataIn1 = 32'd241
; 
32'd10919: dataIn1 = 32'd123
; 
32'd10920: dataIn1 = 32'd125
; 
32'd10921: dataIn1 = 32'd192
; 
32'd10922: dataIn1 = 32'd220
; 
32'd10923: dataIn1 = 32'd244
; 
32'd10924: dataIn1 = 32'd260
; 
32'd10925: dataIn1 = 32'd288
; 
32'd10926: dataIn1 = 32'd94
; 
32'd10927: dataIn1 = 32'd128
; 
32'd10928: dataIn1 = 32'd194
; 
32'd10929: dataIn1 = 32'd221
; 
32'd10930: dataIn1 = 32'd269
; 
32'd10931: dataIn1 = 32'd315
; 
32'd10932: dataIn1 = 32'd323
; 
32'd10933: dataIn1 = 32'd335
; 
32'd10934: dataIn1 = 32'd100
; 
32'd10935: dataIn1 = 32'd134
; 
32'd10936: dataIn1 = 32'd216
; 
32'd10937: dataIn1 = 32'd222
; 
32'd10938: dataIn1 = 32'd233
; 
32'd10939: dataIn1 = 32'd263
; 
32'd10940: dataIn1 = 32'd316
; 
32'd10941: dataIn1 = 32'd109
; 
32'd10942: dataIn1 = 32'd162
; 
32'd10943: dataIn1 = 32'd178
; 
32'd10944: dataIn1 = 32'd223
; 
32'd10945: dataIn1 = 32'd246
; 
32'd10946: dataIn1 = 32'd249
; 
32'd10947: dataIn1 = 32'd292
; 
32'd10948: dataIn1 = 32'd317
; 
32'd10949: dataIn1 = 32'd112
; 
32'd10950: dataIn1 = 32'd181
; 
32'd10951: dataIn1 = 32'd184
; 
32'd10952: dataIn1 = 32'd224
; 
32'd10953: dataIn1 = 32'd118
; 
32'd10954: dataIn1 = 32'd130
; 
32'd10955: dataIn1 = 32'd175
; 
32'd10956: dataIn1 = 32'd225
; 
32'd10957: dataIn1 = 32'd232
; 
32'd10958: dataIn1 = 32'd238
; 
32'd10959: dataIn1 = 32'd254
; 
32'd10960: dataIn1 = 32'd289
; 
32'd10961: dataIn1 = 32'd119
; 
32'd10962: dataIn1 = 32'd152
; 
32'd10963: dataIn1 = 32'd189
; 
32'd10964: dataIn1 = 32'd226
; 
32'd10965: dataIn1 = 32'd236
; 
32'd10966: dataIn1 = 32'd261
; 
32'd10967: dataIn1 = 32'd262
; 
32'd10968: dataIn1 = 32'd120
; 
32'd10969: dataIn1 = 32'd197
; 
32'd10970: dataIn1 = 32'd218
; 
32'd10971: dataIn1 = 32'd227
; 
32'd10972: dataIn1 = 32'd243
; 
32'd10973: dataIn1 = 32'd256
; 
32'd10974: dataIn1 = 32'd122
; 
32'd10975: dataIn1 = 32'd123
; 
32'd10976: dataIn1 = 32'd147
; 
32'd10977: dataIn1 = 32'd228
; 
32'd10978: dataIn1 = 32'd255
; 
32'd10979: dataIn1 = 32'd278
; 
32'd10980: dataIn1 = 32'd285
; 
32'd10981: dataIn1 = 32'd290
; 
32'd10982: dataIn1 = 32'd125
; 
32'd10983: dataIn1 = 32'd193
; 
32'd10984: dataIn1 = 32'd197
; 
32'd10985: dataIn1 = 32'd229
; 
32'd10986: dataIn1 = 32'd230
; 
32'd10987: dataIn1 = 32'd244
; 
32'd10988: dataIn1 = 32'd291
; 
32'd10989: dataIn1 = 32'd297
; 
32'd10990: dataIn1 = 32'd318
; 
32'd10991: dataIn1 = 32'd126
; 
32'd10992: dataIn1 = 32'd184
; 
32'd10993: dataIn1 = 32'd229
; 
32'd10994: dataIn1 = 32'd230
; 
32'd10995: dataIn1 = 32'd247
; 
32'd10996: dataIn1 = 32'd291
; 
32'd10997: dataIn1 = 32'd326
; 
32'd10998: dataIn1 = 32'd128
; 
32'd10999: dataIn1 = 32'd195
; 
32'd11000: dataIn1 = 32'd219
; 
32'd11001: dataIn1 = 32'd231
; 
32'd11002: dataIn1 = 32'd241
; 
32'd11003: dataIn1 = 32'd284
; 
32'd11004: dataIn1 = 32'd315
; 
32'd11005: dataIn1 = 32'd130
; 
32'd11006: dataIn1 = 32'd175
; 
32'd11007: dataIn1 = 32'd225
; 
32'd11008: dataIn1 = 32'd232
; 
32'd11009: dataIn1 = 32'd277
; 
32'd11010: dataIn1 = 32'd319
; 
32'd11011: dataIn1 = 32'd131
; 
32'd11012: dataIn1 = 32'd132
; 
32'd11013: dataIn1 = 32'd222
; 
32'd11014: dataIn1 = 32'd233
; 
32'd11015: dataIn1 = 32'd282
; 
32'd11016: dataIn1 = 32'd287
; 
32'd11017: dataIn1 = 32'd292
; 
32'd11018: dataIn1 = 32'd316
; 
32'd11019: dataIn1 = 32'd320
; 
32'd11020: dataIn1 = 32'd132
; 
32'd11021: dataIn1 = 32'd183
; 
32'd11022: dataIn1 = 32'd199
; 
32'd11023: dataIn1 = 32'd234
; 
32'd11024: dataIn1 = 32'd287
; 
32'd11025: dataIn1 = 32'd293
; 
32'd11026: dataIn1 = 32'd303
; 
32'd11027: dataIn1 = 32'd134
; 
32'd11028: dataIn1 = 32'd200
; 
32'd11029: dataIn1 = 32'd201
; 
32'd11030: dataIn1 = 32'd235
; 
32'd11031: dataIn1 = 32'd251
; 
32'd11032: dataIn1 = 32'd316
; 
32'd11033: dataIn1 = 32'd321
; 
32'd11034: dataIn1 = 32'd337
; 
32'd11035: dataIn1 = 32'd135
; 
32'd11036: dataIn1 = 32'd136
; 
32'd11037: dataIn1 = 32'd226
; 
32'd11038: dataIn1 = 32'd236
; 
32'd11039: dataIn1 = 32'd254
; 
32'd11040: dataIn1 = 32'd261
; 
32'd11041: dataIn1 = 32'd273
; 
32'd11042: dataIn1 = 32'd294
; 
32'd11043: dataIn1 = 32'd322
; 
32'd11044: dataIn1 = 32'd145
; 
32'd11045: dataIn1 = 32'd148
; 
32'd11046: dataIn1 = 32'd176
; 
32'd11047: dataIn1 = 32'd237
; 
32'd11048: dataIn1 = 32'd283
; 
32'd11049: dataIn1 = 32'd313
; 
32'd11050: dataIn1 = 32'd148
; 
32'd11051: dataIn1 = 32'd167
; 
32'd11052: dataIn1 = 32'd225
; 
32'd11053: dataIn1 = 32'd238
; 
32'd11054: dataIn1 = 32'd245
; 
32'd11055: dataIn1 = 32'd266
; 
32'd11056: dataIn1 = 32'd289
; 
32'd11057: dataIn1 = 32'd149
; 
32'd11058: dataIn1 = 32'd206
; 
32'd11059: dataIn1 = 32'd215
; 
32'd11060: dataIn1 = 32'd239
; 
32'd11061: dataIn1 = 32'd246
; 
32'd11062: dataIn1 = 32'd282
; 
32'd11063: dataIn1 = 32'd295
; 
32'd11064: dataIn1 = 32'd308
; 
32'd11065: dataIn1 = 32'd156
; 
32'd11066: dataIn1 = 32'd166
; 
32'd11067: dataIn1 = 32'd205
; 
32'd11068: dataIn1 = 32'd240
; 
32'd11069: dataIn1 = 32'd264
; 
32'd11070: dataIn1 = 32'd304
; 
32'd11071: dataIn1 = 32'd166
; 
32'd11072: dataIn1 = 32'd219
; 
32'd11073: dataIn1 = 32'd231
; 
32'd11074: dataIn1 = 32'd241
; 
32'd11075: dataIn1 = 32'd252
; 
32'd11076: dataIn1 = 32'd301
; 
32'd11077: dataIn1 = 32'd315
; 
32'd11078: dataIn1 = 32'd359
; 
32'd11079: dataIn1 = 32'd162
; 
32'd11080: dataIn1 = 32'd174
; 
32'd11081: dataIn1 = 32'd181
; 
32'd11082: dataIn1 = 32'd242
; 
32'd11083: dataIn1 = 32'd247
; 
32'd11084: dataIn1 = 32'd300
; 
32'd11085: dataIn1 = 32'd312
; 
32'd11086: dataIn1 = 32'd317
; 
32'd11087: dataIn1 = 32'd161
; 
32'd11088: dataIn1 = 32'd194
; 
32'd11089: dataIn1 = 32'd227
; 
32'd11090: dataIn1 = 32'd243
; 
32'd11091: dataIn1 = 32'd323
; 
32'd11092: dataIn1 = 32'd193
; 
32'd11093: dataIn1 = 32'd220
; 
32'd11094: dataIn1 = 32'd229
; 
32'd11095: dataIn1 = 32'd244
; 
32'd11096: dataIn1 = 32'd285
; 
32'd11097: dataIn1 = 32'd291
; 
32'd11098: dataIn1 = 32'd310
; 
32'd11099: dataIn1 = 32'd318
; 
32'd11100: dataIn1 = 32'd360
; 
32'd11101: dataIn1 = 32'd148
; 
32'd11102: dataIn1 = 32'd213
; 
32'd11103: dataIn1 = 32'd238
; 
32'd11104: dataIn1 = 32'd245
; 
32'd11105: dataIn1 = 32'd254
; 
32'd11106: dataIn1 = 32'd266
; 
32'd11107: dataIn1 = 32'd313
; 
32'd11108: dataIn1 = 32'd324
; 
32'd11109: dataIn1 = 32'd162
; 
32'd11110: dataIn1 = 32'd223
; 
32'd11111: dataIn1 = 32'd239
; 
32'd11112: dataIn1 = 32'd246
; 
32'd11113: dataIn1 = 32'd270
; 
32'd11114: dataIn1 = 32'd317
; 
32'd11115: dataIn1 = 32'd325
; 
32'd11116: dataIn1 = 32'd218
; 
32'd11117: dataIn1 = 32'd230
; 
32'd11118: dataIn1 = 32'd242
; 
32'd11119: dataIn1 = 32'd247
; 
32'd11120: dataIn1 = 32'd256
; 
32'd11121: dataIn1 = 32'd300
; 
32'd11122: dataIn1 = 32'd312
; 
32'd11123: dataIn1 = 32'd314
; 
32'd11124: dataIn1 = 32'd326
; 
32'd11125: dataIn1 = 32'd343
; 
32'd11126: dataIn1 = 32'd355
; 
32'd11127: dataIn1 = 32'd361
; 
32'd11128: dataIn1 = 32'd389
; 
32'd11129: dataIn1 = 32'd404
; 
32'd11130: dataIn1 = 32'd112
; 
32'd11131: dataIn1 = 32'd169
; 
32'd11132: dataIn1 = 32'd203
; 
32'd11133: dataIn1 = 32'd248
; 
32'd11134: dataIn1 = 32'd300
; 
32'd11135: dataIn1 = 32'd198
; 
32'd11136: dataIn1 = 32'd200
; 
32'd11137: dataIn1 = 32'd223
; 
32'd11138: dataIn1 = 32'd249
; 
32'd11139: dataIn1 = 32'd292
; 
32'd11140: dataIn1 = 32'd327
; 
32'd11141: dataIn1 = 32'd358
; 
32'd11142: dataIn1 = 32'd183
; 
32'd11143: dataIn1 = 32'd190
; 
32'd11144: dataIn1 = 32'd202
; 
32'd11145: dataIn1 = 32'd250
; 
32'd11146: dataIn1 = 32'd259
; 
32'd11147: dataIn1 = 32'd157
; 
32'd11148: dataIn1 = 32'd160
; 
32'd11149: dataIn1 = 32'd235
; 
32'd11150: dataIn1 = 32'd251
; 
32'd11151: dataIn1 = 32'd311
; 
32'd11152: dataIn1 = 32'd328
; 
32'd11153: dataIn1 = 32'd348
; 
32'd11154: dataIn1 = 32'd154
; 
32'd11155: dataIn1 = 32'd164
; 
32'd11156: dataIn1 = 32'd241
; 
32'd11157: dataIn1 = 32'd252
; 
32'd11158: dataIn1 = 32'd301
; 
32'd11159: dataIn1 = 32'd159
; 
32'd11160: dataIn1 = 32'd176
; 
32'd11161: dataIn1 = 32'd197
; 
32'd11162: dataIn1 = 32'd253
; 
32'd11163: dataIn1 = 32'd280
; 
32'd11164: dataIn1 = 32'd329
; 
32'd11165: dataIn1 = 32'd336
; 
32'd11166: dataIn1 = 32'd346
; 
32'd11167: dataIn1 = 32'd357
; 
32'd11168: dataIn1 = 32'd225
; 
32'd11169: dataIn1 = 32'd236
; 
32'd11170: dataIn1 = 32'd245
; 
32'd11171: dataIn1 = 32'd254
; 
32'd11172: dataIn1 = 32'd273
; 
32'd11173: dataIn1 = 32'd324
; 
32'd11174: dataIn1 = 32'd330
; 
32'd11175: dataIn1 = 32'd339
; 
32'd11176: dataIn1 = 32'd191
; 
32'd11177: dataIn1 = 32'd214
; 
32'd11178: dataIn1 = 32'd228
; 
32'd11179: dataIn1 = 32'd255
; 
32'd11180: dataIn1 = 32'd278
; 
32'd11181: dataIn1 = 32'd290
; 
32'd11182: dataIn1 = 32'd302
; 
32'd11183: dataIn1 = 32'd319
; 
32'd11184: dataIn1 = 32'd331
; 
32'd11185: dataIn1 = 32'd197
; 
32'd11186: dataIn1 = 32'd227
; 
32'd11187: dataIn1 = 32'd247
; 
32'd11188: dataIn1 = 32'd256
; 
32'd11189: dataIn1 = 32'd297
; 
32'd11190: dataIn1 = 32'd329
; 
32'd11191: dataIn1 = 32'd355
; 
32'd11192: dataIn1 = 32'd423
; 
32'd11193: dataIn1 = 32'd156
; 
32'd11194: dataIn1 = 32'd157
; 
32'd11195: dataIn1 = 32'd212
; 
32'd11196: dataIn1 = 32'd257
; 
32'd11197: dataIn1 = 32'd328
; 
32'd11198: dataIn1 = 32'd349
; 
32'd11199: dataIn1 = 32'd351
; 
32'd11200: dataIn1 = 32'd157
; 
32'd11201: dataIn1 = 32'd208
; 
32'd11202: dataIn1 = 32'd217
; 
32'd11203: dataIn1 = 32'd258
; 
32'd11204: dataIn1 = 32'd296
; 
32'd11205: dataIn1 = 32'd333
; 
32'd11206: dataIn1 = 32'd348
; 
32'd11207: dataIn1 = 32'd362
; 
32'd11208: dataIn1 = 32'd167
; 
32'd11209: dataIn1 = 32'd202
; 
32'd11210: dataIn1 = 32'd250
; 
32'd11211: dataIn1 = 32'd259
; 
32'd11212: dataIn1 = 32'd277
; 
32'd11213: dataIn1 = 32'd307
; 
32'd11214: dataIn1 = 32'd332
; 
32'd11215: dataIn1 = 32'd363
; 
32'd11216: dataIn1 = 32'd171
; 
32'd11217: dataIn1 = 32'd204
; 
32'd11218: dataIn1 = 32'd220
; 
32'd11219: dataIn1 = 32'd260
; 
32'd11220: dataIn1 = 32'd263
; 
32'd11221: dataIn1 = 32'd296
; 
32'd11222: dataIn1 = 32'd318
; 
32'd11223: dataIn1 = 32'd354
; 
32'd11224: dataIn1 = 32'd364
; 
32'd11225: dataIn1 = 32'd189
; 
32'd11226: dataIn1 = 32'd226
; 
32'd11227: dataIn1 = 32'd236
; 
32'd11228: dataIn1 = 32'd261
; 
32'd11229: dataIn1 = 32'd275
; 
32'd11230: dataIn1 = 32'd286
; 
32'd11231: dataIn1 = 32'd294
; 
32'd11232: dataIn1 = 32'd322
; 
32'd11233: dataIn1 = 32'd182
; 
32'd11234: dataIn1 = 32'd203
; 
32'd11235: dataIn1 = 32'd226
; 
32'd11236: dataIn1 = 32'd262
; 
32'd11237: dataIn1 = 32'd267
; 
32'd11238: dataIn1 = 32'd276
; 
32'd11239: dataIn1 = 32'd334
; 
32'd11240: dataIn1 = 32'd342
; 
32'd11241: dataIn1 = 32'd365
; 
32'd11242: dataIn1 = 32'd171
; 
32'd11243: dataIn1 = 32'd222
; 
32'd11244: dataIn1 = 32'd260
; 
32'd11245: dataIn1 = 32'd263
; 
32'd11246: dataIn1 = 32'd279
; 
32'd11247: dataIn1 = 32'd288
; 
32'd11248: dataIn1 = 32'd321
; 
32'd11249: dataIn1 = 32'd362
; 
32'd11250: dataIn1 = 32'd364
; 
32'd11251: dataIn1 = 32'd366
; 
32'd11252: dataIn1 = 32'd376
; 
32'd11253: dataIn1 = 32'd156
; 
32'd11254: dataIn1 = 32'd177
; 
32'd11255: dataIn1 = 32'd240
; 
32'd11256: dataIn1 = 32'd264
; 
32'd11257: dataIn1 = 32'd274
; 
32'd11258: dataIn1 = 32'd328
; 
32'd11259: dataIn1 = 32'd345
; 
32'd11260: dataIn1 = 32'd351
; 
32'd11261: dataIn1 = 32'd367
; 
32'd11262: dataIn1 = 32'd102
; 
32'd11263: dataIn1 = 32'd179
; 
32'd11264: dataIn1 = 32'd182
; 
32'd11265: dataIn1 = 32'd265
; 
32'd11266: dataIn1 = 32'd275
; 
32'd11267: dataIn1 = 32'd306
; 
32'd11268: dataIn1 = 32'd335
; 
32'd11269: dataIn1 = 32'd148
; 
32'd11270: dataIn1 = 32'd238
; 
32'd11271: dataIn1 = 32'd245
; 
32'd11272: dataIn1 = 32'd266
; 
32'd11273: dataIn1 = 32'd324
; 
32'd11274: dataIn1 = 32'd333
; 
32'd11275: dataIn1 = 32'd349
; 
32'd11276: dataIn1 = 32'd368
; 
32'd11277: dataIn1 = 32'd152
; 
32'd11278: dataIn1 = 32'd214
; 
32'd11279: dataIn1 = 32'd262
; 
32'd11280: dataIn1 = 32'd267
; 
32'd11281: dataIn1 = 32'd302
; 
32'd11282: dataIn1 = 32'd322
; 
32'd11283: dataIn1 = 32'd334
; 
32'd11284: dataIn1 = 32'd154
; 
32'd11285: dataIn1 = 32'd206
; 
32'd11286: dataIn1 = 32'd210
; 
32'd11287: dataIn1 = 32'd268
; 
32'd11288: dataIn1 = 32'd306
; 
32'd11289: dataIn1 = 32'd359
; 
32'd11290: dataIn1 = 32'd369
; 
32'd11291: dataIn1 = 32'd371
; 
32'd11292: dataIn1 = 32'd159
; 
32'd11293: dataIn1 = 32'd179
; 
32'd11294: dataIn1 = 32'd221
; 
32'd11295: dataIn1 = 32'd269
; 
32'd11296: dataIn1 = 32'd299
; 
32'd11297: dataIn1 = 32'd329
; 
32'd11298: dataIn1 = 32'd370
; 
32'd11299: dataIn1 = 32'd375
; 
32'd11300: dataIn1 = 32'd388
; 
32'd11301: dataIn1 = 32'd406
; 
32'd11302: dataIn1 = 32'd162
; 
32'd11303: dataIn1 = 32'd169
; 
32'd11304: dataIn1 = 32'd246
; 
32'd11305: dataIn1 = 32'd270
; 
32'd11306: dataIn1 = 32'd272
; 
32'd11307: dataIn1 = 32'd308
; 
32'd11308: dataIn1 = 32'd350
; 
32'd11309: dataIn1 = 32'd167
; 
32'd11310: dataIn1 = 32'd202
; 
32'd11311: dataIn1 = 32'd212
; 
32'd11312: dataIn1 = 32'd271
; 
32'd11313: dataIn1 = 32'd304
; 
32'd11314: dataIn1 = 32'd332
; 
32'd11315: dataIn1 = 32'd349
; 
32'd11316: dataIn1 = 32'd356
; 
32'd11317: dataIn1 = 32'd169
; 
32'd11318: dataIn1 = 32'd206
; 
32'd11319: dataIn1 = 32'd270
; 
32'd11320: dataIn1 = 32'd272
; 
32'd11321: dataIn1 = 32'd305
; 
32'd11322: dataIn1 = 32'd371
; 
32'd11323: dataIn1 = 32'd175
; 
32'd11324: dataIn1 = 32'd236
; 
32'd11325: dataIn1 = 32'd254
; 
32'd11326: dataIn1 = 32'd273
; 
32'd11327: dataIn1 = 32'd319
; 
32'd11328: dataIn1 = 32'd339
; 
32'd11329: dataIn1 = 32'd156
; 
32'd11330: dataIn1 = 32'd177
; 
32'd11331: dataIn1 = 32'd264
; 
32'd11332: dataIn1 = 32'd274
; 
32'd11333: dataIn1 = 32'd179
; 
32'd11334: dataIn1 = 32'd261
; 
32'd11335: dataIn1 = 32'd265
; 
32'd11336: dataIn1 = 32'd275
; 
32'd11337: dataIn1 = 32'd335
; 
32'd11338: dataIn1 = 32'd342
; 
32'd11339: dataIn1 = 32'd370
; 
32'd11340: dataIn1 = 32'd372
; 
32'd11341: dataIn1 = 32'd182
; 
32'd11342: dataIn1 = 32'd196
; 
32'd11343: dataIn1 = 32'd262
; 
32'd11344: dataIn1 = 32'd276
; 
32'd11345: dataIn1 = 32'd306
; 
32'd11346: dataIn1 = 32'd183
; 
32'd11347: dataIn1 = 32'd232
; 
32'd11348: dataIn1 = 32'd259
; 
32'd11349: dataIn1 = 32'd277
; 
32'd11350: dataIn1 = 32'd307
; 
32'd11351: dataIn1 = 32'd363
; 
32'd11352: dataIn1 = 32'd373
; 
32'd11353: dataIn1 = 32'd191
; 
32'd11354: dataIn1 = 32'd228
; 
32'd11355: dataIn1 = 32'd255
; 
32'd11356: dataIn1 = 32'd278
; 
32'd11357: dataIn1 = 32'd279
; 
32'd11358: dataIn1 = 32'd293
; 
32'd11359: dataIn1 = 32'd331
; 
32'd11360: dataIn1 = 32'd192
; 
32'd11361: dataIn1 = 32'd263
; 
32'd11362: dataIn1 = 32'd278
; 
32'd11363: dataIn1 = 32'd279
; 
32'd11364: dataIn1 = 32'd288
; 
32'd11365: dataIn1 = 32'd338
; 
32'd11366: dataIn1 = 32'd344
; 
32'd11367: dataIn1 = 32'd353
; 
32'd11368: dataIn1 = 32'd197
; 
32'd11369: dataIn1 = 32'd204
; 
32'd11370: dataIn1 = 32'd253
; 
32'd11371: dataIn1 = 32'd280
; 
32'd11372: dataIn1 = 32'd297
; 
32'd11373: dataIn1 = 32'd336
; 
32'd11374: dataIn1 = 32'd354
; 
32'd11375: dataIn1 = 32'd198
; 
32'd11376: dataIn1 = 32'd207
; 
32'd11377: dataIn1 = 32'd218
; 
32'd11378: dataIn1 = 32'd281
; 
32'd11379: dataIn1 = 32'd314
; 
32'd11380: dataIn1 = 32'd199
; 
32'd11381: dataIn1 = 32'd233
; 
32'd11382: dataIn1 = 32'd239
; 
32'd11383: dataIn1 = 32'd282
; 
32'd11384: dataIn1 = 32'd320
; 
32'd11385: dataIn1 = 32'd325
; 
32'd11386: dataIn1 = 32'd340
; 
32'd11387: dataIn1 = 32'd204
; 
32'd11388: dataIn1 = 32'd208
; 
32'd11389: dataIn1 = 32'd237
; 
32'd11390: dataIn1 = 32'd283
; 
32'd11391: dataIn1 = 32'd296
; 
32'd11392: dataIn1 = 32'd336
; 
32'd11393: dataIn1 = 32'd354
; 
32'd11394: dataIn1 = 32'd143
; 
32'd11395: dataIn1 = 32'd205
; 
32'd11396: dataIn1 = 32'd231
; 
32'd11397: dataIn1 = 32'd284
; 
32'd11398: dataIn1 = 32'd298
; 
32'd11399: dataIn1 = 32'd211
; 
32'd11400: dataIn1 = 32'd228
; 
32'd11401: dataIn1 = 32'd244
; 
32'd11402: dataIn1 = 32'd285
; 
32'd11403: dataIn1 = 32'd309
; 
32'd11404: dataIn1 = 32'd344
; 
32'd11405: dataIn1 = 32'd360
; 
32'd11406: dataIn1 = 32'd378
; 
32'd11407: dataIn1 = 32'd179
; 
32'd11408: dataIn1 = 32'd213
; 
32'd11409: dataIn1 = 32'd261
; 
32'd11410: dataIn1 = 32'd286
; 
32'd11411: dataIn1 = 32'd299
; 
32'd11412: dataIn1 = 32'd216
; 
32'd11413: dataIn1 = 32'd233
; 
32'd11414: dataIn1 = 32'd234
; 
32'd11415: dataIn1 = 32'd287
; 
32'd11416: dataIn1 = 32'd293
; 
32'd11417: dataIn1 = 32'd303
; 
32'd11418: dataIn1 = 32'd338
; 
32'd11419: dataIn1 = 32'd347
; 
32'd11420: dataIn1 = 32'd352
; 
32'd11421: dataIn1 = 32'd220
; 
32'd11422: dataIn1 = 32'd263
; 
32'd11423: dataIn1 = 32'd279
; 
32'd11424: dataIn1 = 32'd288
; 
32'd11425: dataIn1 = 32'd344
; 
32'd11426: dataIn1 = 32'd167
; 
32'd11427: dataIn1 = 32'd225
; 
32'd11428: dataIn1 = 32'd238
; 
32'd11429: dataIn1 = 32'd289
; 
32'd11430: dataIn1 = 32'd339
; 
32'd11431: dataIn1 = 32'd356
; 
32'd11432: dataIn1 = 32'd211
; 
32'd11433: dataIn1 = 32'd228
; 
32'd11434: dataIn1 = 32'd255
; 
32'd11435: dataIn1 = 32'd290
; 
32'd11436: dataIn1 = 32'd302
; 
32'd11437: dataIn1 = 32'd309
; 
32'd11438: dataIn1 = 32'd331
; 
32'd11439: dataIn1 = 32'd229
; 
32'd11440: dataIn1 = 32'd230
; 
32'd11441: dataIn1 = 32'd244
; 
32'd11442: dataIn1 = 32'd291
; 
32'd11443: dataIn1 = 32'd310
; 
32'd11444: dataIn1 = 32'd223
; 
32'd11445: dataIn1 = 32'd233
; 
32'd11446: dataIn1 = 32'd249
; 
32'd11447: dataIn1 = 32'd292
; 
32'd11448: dataIn1 = 32'd320
; 
32'd11449: dataIn1 = 32'd337
; 
32'd11450: dataIn1 = 32'd234
; 
32'd11451: dataIn1 = 32'd278
; 
32'd11452: dataIn1 = 32'd287
; 
32'd11453: dataIn1 = 32'd293
; 
32'd11454: dataIn1 = 32'd338
; 
32'd11455: dataIn1 = 32'd347
; 
32'd11456: dataIn1 = 32'd213
; 
32'd11457: dataIn1 = 32'd236
; 
32'd11458: dataIn1 = 32'd261
; 
32'd11459: dataIn1 = 32'd294
; 
32'd11460: dataIn1 = 32'd330
; 
32'd11461: dataIn1 = 32'd199
; 
32'd11462: dataIn1 = 32'd206
; 
32'd11463: dataIn1 = 32'd239
; 
32'd11464: dataIn1 = 32'd295
; 
32'd11465: dataIn1 = 32'd371
; 
32'd11466: dataIn1 = 32'd374
; 
32'd11467: dataIn1 = 32'd377
; 
32'd11468: dataIn1 = 32'd391
; 
32'd11469: dataIn1 = 32'd258
; 
32'd11470: dataIn1 = 32'd260
; 
32'd11471: dataIn1 = 32'd283
; 
32'd11472: dataIn1 = 32'd296
; 
32'd11473: dataIn1 = 32'd229
; 
32'd11474: dataIn1 = 32'd256
; 
32'd11475: dataIn1 = 32'd280
; 
32'd11476: dataIn1 = 32'd297
; 
32'd11477: dataIn1 = 32'd326
; 
32'd11478: dataIn1 = 32'd346
; 
32'd11479: dataIn1 = 32'd355
; 
32'd11480: dataIn1 = 32'd407
; 
32'd11481: dataIn1 = 32'd428
; 
32'd11482: dataIn1 = 32'd429
; 
32'd11483: dataIn1 = 32'd177
; 
32'd11484: dataIn1 = 32'd207
; 
32'd11485: dataIn1 = 32'd284
; 
32'd11486: dataIn1 = 32'd298
; 
32'd11487: dataIn1 = 32'd323
; 
32'd11488: dataIn1 = 32'd345
; 
32'd11489: dataIn1 = 32'd408
; 
32'd11490: dataIn1 = 32'd213
; 
32'd11491: dataIn1 = 32'd269
; 
32'd11492: dataIn1 = 32'd286
; 
32'd11493: dataIn1 = 32'd299
; 
32'd11494: dataIn1 = 32'd370
; 
32'd11495: dataIn1 = 32'd375
; 
32'd11496: dataIn1 = 32'd396
; 
32'd11497: dataIn1 = 32'd242
; 
32'd11498: dataIn1 = 32'd247
; 
32'd11499: dataIn1 = 32'd248
; 
32'd11500: dataIn1 = 32'd300
; 
32'd11501: dataIn1 = 32'd305
; 
32'd11502: dataIn1 = 32'd310
; 
32'd11503: dataIn1 = 32'd389
; 
32'd11504: dataIn1 = 32'd409
; 
32'd11505: dataIn1 = 32'd202
; 
32'd11506: dataIn1 = 32'd241
; 
32'd11507: dataIn1 = 32'd252
; 
32'd11508: dataIn1 = 32'd301
; 
32'd11509: dataIn1 = 32'd307
; 
32'd11510: dataIn1 = 32'd359
; 
32'd11511: dataIn1 = 32'd385
; 
32'd11512: dataIn1 = 32'd387
; 
32'd11513: dataIn1 = 32'd394
; 
32'd11514: dataIn1 = 32'd401
; 
32'd11515: dataIn1 = 32'd255
; 
32'd11516: dataIn1 = 32'd267
; 
32'd11517: dataIn1 = 32'd290
; 
32'd11518: dataIn1 = 32'd302
; 
32'd11519: dataIn1 = 32'd410
; 
32'd11520: dataIn1 = 32'd431
; 
32'd11521: dataIn1 = 32'd199
; 
32'd11522: dataIn1 = 32'd234
; 
32'd11523: dataIn1 = 32'd287
; 
32'd11524: dataIn1 = 32'd303
; 
32'd11525: dataIn1 = 32'd374
; 
32'd11526: dataIn1 = 32'd202
; 
32'd11527: dataIn1 = 32'd240
; 
32'd11528: dataIn1 = 32'd271
; 
32'd11529: dataIn1 = 32'd304
; 
32'd11530: dataIn1 = 32'd351
; 
32'd11531: dataIn1 = 32'd203
; 
32'd11532: dataIn1 = 32'd272
; 
32'd11533: dataIn1 = 32'd300
; 
32'd11534: dataIn1 = 32'd305
; 
32'd11535: dataIn1 = 32'd341
; 
32'd11536: dataIn1 = 32'd265
; 
32'd11537: dataIn1 = 32'd268
; 
32'd11538: dataIn1 = 32'd276
; 
32'd11539: dataIn1 = 32'd306
; 
32'd11540: dataIn1 = 32'd342
; 
32'd11541: dataIn1 = 32'd369
; 
32'd11542: dataIn1 = 32'd259
; 
32'd11543: dataIn1 = 32'd277
; 
32'd11544: dataIn1 = 32'd301
; 
32'd11545: dataIn1 = 32'd307
; 
32'd11546: dataIn1 = 32'd363
; 
32'd11547: dataIn1 = 32'd385
; 
32'd11548: dataIn1 = 32'd402
; 
32'd11549: dataIn1 = 32'd206
; 
32'd11550: dataIn1 = 32'd239
; 
32'd11551: dataIn1 = 32'd270
; 
32'd11552: dataIn1 = 32'd308
; 
32'd11553: dataIn1 = 32'd350
; 
32'd11554: dataIn1 = 32'd211
; 
32'd11555: dataIn1 = 32'd285
; 
32'd11556: dataIn1 = 32'd290
; 
32'd11557: dataIn1 = 32'd309
; 
32'd11558: dataIn1 = 32'd341
; 
32'd11559: dataIn1 = 32'd411
; 
32'd11560: dataIn1 = 32'd448
; 
32'd11561: dataIn1 = 32'd244
; 
32'd11562: dataIn1 = 32'd291
; 
32'd11563: dataIn1 = 32'd300
; 
32'd11564: dataIn1 = 32'd310
; 
32'd11565: dataIn1 = 32'd389
; 
32'd11566: dataIn1 = 32'd403
; 
32'd11567: dataIn1 = 32'd177
; 
32'd11568: dataIn1 = 32'd200
; 
32'd11569: dataIn1 = 32'd251
; 
32'd11570: dataIn1 = 32'd311
; 
32'd11571: dataIn1 = 32'd327
; 
32'd11572: dataIn1 = 32'd337
; 
32'd11573: dataIn1 = 32'd345
; 
32'd11574: dataIn1 = 32'd405
; 
32'd11575: dataIn1 = 32'd412
; 
32'd11576: dataIn1 = 32'd198
; 
32'd11577: dataIn1 = 32'd242
; 
32'd11578: dataIn1 = 32'd247
; 
32'd11579: dataIn1 = 32'd312
; 
32'd11580: dataIn1 = 32'd343
; 
32'd11581: dataIn1 = 32'd213
; 
32'd11582: dataIn1 = 32'd237
; 
32'd11583: dataIn1 = 32'd245
; 
32'd11584: dataIn1 = 32'd313
; 
32'd11585: dataIn1 = 32'd330
; 
32'd11586: dataIn1 = 32'd333
; 
32'd11587: dataIn1 = 32'd357
; 
32'd11588: dataIn1 = 32'd368
; 
32'd11589: dataIn1 = 32'd395
; 
32'd11590: dataIn1 = 32'd218
; 
32'd11591: dataIn1 = 32'd247
; 
32'd11592: dataIn1 = 32'd281
; 
32'd11593: dataIn1 = 32'd314
; 
32'd11594: dataIn1 = 32'd361
; 
32'd11595: dataIn1 = 32'd221
; 
32'd11596: dataIn1 = 32'd231
; 
32'd11597: dataIn1 = 32'd241
; 
32'd11598: dataIn1 = 32'd315
; 
32'd11599: dataIn1 = 32'd383
; 
32'd11600: dataIn1 = 32'd392
; 
32'd11601: dataIn1 = 32'd413
; 
32'd11602: dataIn1 = 32'd414
; 
32'd11603: dataIn1 = 32'd458
; 
32'd11604: dataIn1 = 32'd222
; 
32'd11605: dataIn1 = 32'd233
; 
32'd11606: dataIn1 = 32'd235
; 
32'd11607: dataIn1 = 32'd316
; 
32'd11608: dataIn1 = 32'd321
; 
32'd11609: dataIn1 = 32'd352
; 
32'd11610: dataIn1 = 32'd223
; 
32'd11611: dataIn1 = 32'd242
; 
32'd11612: dataIn1 = 32'd246
; 
32'd11613: dataIn1 = 32'd317
; 
32'd11614: dataIn1 = 32'd325
; 
32'd11615: dataIn1 = 32'd343
; 
32'd11616: dataIn1 = 32'd350
; 
32'd11617: dataIn1 = 32'd229
; 
32'd11618: dataIn1 = 32'd244
; 
32'd11619: dataIn1 = 32'd260
; 
32'd11620: dataIn1 = 32'd318
; 
32'd11621: dataIn1 = 32'd360
; 
32'd11622: dataIn1 = 32'd399
; 
32'd11623: dataIn1 = 32'd407
; 
32'd11624: dataIn1 = 32'd232
; 
32'd11625: dataIn1 = 32'd255
; 
32'd11626: dataIn1 = 32'd273
; 
32'd11627: dataIn1 = 32'd319
; 
32'd11628: dataIn1 = 32'd373
; 
32'd11629: dataIn1 = 32'd233
; 
32'd11630: dataIn1 = 32'd282
; 
32'd11631: dataIn1 = 32'd292
; 
32'd11632: dataIn1 = 32'd320
; 
32'd11633: dataIn1 = 32'd340
; 
32'd11634: dataIn1 = 32'd352
; 
32'd11635: dataIn1 = 32'd384
; 
32'd11636: dataIn1 = 32'd393
; 
32'd11637: dataIn1 = 32'd400
; 
32'd11638: dataIn1 = 32'd235
; 
32'd11639: dataIn1 = 32'd263
; 
32'd11640: dataIn1 = 32'd316
; 
32'd11641: dataIn1 = 32'd321
; 
32'd11642: dataIn1 = 32'd366
; 
32'd11643: dataIn1 = 32'd236
; 
32'd11644: dataIn1 = 32'd261
; 
32'd11645: dataIn1 = 32'd267
; 
32'd11646: dataIn1 = 32'd322
; 
32'd11647: dataIn1 = 32'd365
; 
32'd11648: dataIn1 = 32'd372
; 
32'd11649: dataIn1 = 32'd379
; 
32'd11650: dataIn1 = 32'd221
; 
32'd11651: dataIn1 = 32'd243
; 
32'd11652: dataIn1 = 32'd298
; 
32'd11653: dataIn1 = 32'd323
; 
32'd11654: dataIn1 = 32'd388
; 
32'd11655: dataIn1 = 32'd414
; 
32'd11656: dataIn1 = 32'd459
; 
32'd11657: dataIn1 = 32'd245
; 
32'd11658: dataIn1 = 32'd254
; 
32'd11659: dataIn1 = 32'd266
; 
32'd11660: dataIn1 = 32'd324
; 
32'd11661: dataIn1 = 32'd368
; 
32'd11662: dataIn1 = 32'd380
; 
32'd11663: dataIn1 = 32'd246
; 
32'd11664: dataIn1 = 32'd282
; 
32'd11665: dataIn1 = 32'd317
; 
32'd11666: dataIn1 = 32'd325
; 
32'd11667: dataIn1 = 32'd340
; 
32'd11668: dataIn1 = 32'd230
; 
32'd11669: dataIn1 = 32'd247
; 
32'd11670: dataIn1 = 32'd297
; 
32'd11671: dataIn1 = 32'd326
; 
32'd11672: dataIn1 = 32'd198
; 
32'd11673: dataIn1 = 32'd249
; 
32'd11674: dataIn1 = 32'd311
; 
32'd11675: dataIn1 = 32'd327
; 
32'd11676: dataIn1 = 32'd358
; 
32'd11677: dataIn1 = 32'd408
; 
32'd11678: dataIn1 = 32'd412
; 
32'd11679: dataIn1 = 32'd415
; 
32'd11680: dataIn1 = 32'd251
; 
32'd11681: dataIn1 = 32'd257
; 
32'd11682: dataIn1 = 32'd264
; 
32'd11683: dataIn1 = 32'd328
; 
32'd11684: dataIn1 = 32'd348
; 
32'd11685: dataIn1 = 32'd367
; 
32'd11686: dataIn1 = 32'd253
; 
32'd11687: dataIn1 = 32'd256
; 
32'd11688: dataIn1 = 32'd269
; 
32'd11689: dataIn1 = 32'd329
; 
32'd11690: dataIn1 = 32'd346
; 
32'd11691: dataIn1 = 32'd388
; 
32'd11692: dataIn1 = 32'd254
; 
32'd11693: dataIn1 = 32'd294
; 
32'd11694: dataIn1 = 32'd313
; 
32'd11695: dataIn1 = 32'd330
; 
32'd11696: dataIn1 = 32'd379
; 
32'd11697: dataIn1 = 32'd380
; 
32'd11698: dataIn1 = 32'd396
; 
32'd11699: dataIn1 = 32'd416
; 
32'd11700: dataIn1 = 32'd452
; 
32'd11701: dataIn1 = 32'd255
; 
32'd11702: dataIn1 = 32'd278
; 
32'd11703: dataIn1 = 32'd290
; 
32'd11704: dataIn1 = 32'd331
; 
32'd11705: dataIn1 = 32'd353
; 
32'd11706: dataIn1 = 32'd410
; 
32'd11707: dataIn1 = 32'd427
; 
32'd11708: dataIn1 = 32'd202
; 
32'd11709: dataIn1 = 32'd259
; 
32'd11710: dataIn1 = 32'd271
; 
32'd11711: dataIn1 = 32'd332
; 
32'd11712: dataIn1 = 32'd385
; 
32'd11713: dataIn1 = 32'd387
; 
32'd11714: dataIn1 = 32'd390
; 
32'd11715: dataIn1 = 32'd258
; 
32'd11716: dataIn1 = 32'd266
; 
32'd11717: dataIn1 = 32'd313
; 
32'd11718: dataIn1 = 32'd333
; 
32'd11719: dataIn1 = 32'd381
; 
32'd11720: dataIn1 = 32'd397
; 
32'd11721: dataIn1 = 32'd417
; 
32'd11722: dataIn1 = 32'd440
; 
32'd11723: dataIn1 = 32'd203
; 
32'd11724: dataIn1 = 32'd262
; 
32'd11725: dataIn1 = 32'd267
; 
32'd11726: dataIn1 = 32'd334
; 
32'd11727: dataIn1 = 32'd341
; 
32'd11728: dataIn1 = 32'd221
; 
32'd11729: dataIn1 = 32'd265
; 
32'd11730: dataIn1 = 32'd275
; 
32'd11731: dataIn1 = 32'd335
; 
32'd11732: dataIn1 = 32'd369
; 
32'd11733: dataIn1 = 32'd406
; 
32'd11734: dataIn1 = 32'd418
; 
32'd11735: dataIn1 = 32'd460
; 
32'd11736: dataIn1 = 32'd253
; 
32'd11737: dataIn1 = 32'd280
; 
32'd11738: dataIn1 = 32'd283
; 
32'd11739: dataIn1 = 32'd336
; 
32'd11740: dataIn1 = 32'd357
; 
32'd11741: dataIn1 = 32'd381
; 
32'd11742: dataIn1 = 32'd235
; 
32'd11743: dataIn1 = 32'd292
; 
32'd11744: dataIn1 = 32'd311
; 
32'd11745: dataIn1 = 32'd337
; 
32'd11746: dataIn1 = 32'd384
; 
32'd11747: dataIn1 = 32'd419
; 
32'd11748: dataIn1 = 32'd464
; 
32'd11749: dataIn1 = 32'd279
; 
32'd11750: dataIn1 = 32'd287
; 
32'd11751: dataIn1 = 32'd293
; 
32'd11752: dataIn1 = 32'd338
; 
32'd11753: dataIn1 = 32'd347
; 
32'd11754: dataIn1 = 32'd376
; 
32'd11755: dataIn1 = 32'd386
; 
32'd11756: dataIn1 = 32'd254
; 
32'd11757: dataIn1 = 32'd273
; 
32'd11758: dataIn1 = 32'd289
; 
32'd11759: dataIn1 = 32'd339
; 
32'd11760: dataIn1 = 32'd380
; 
32'd11761: dataIn1 = 32'd382
; 
32'd11762: dataIn1 = 32'd398
; 
32'd11763: dataIn1 = 32'd282
; 
32'd11764: dataIn1 = 32'd320
; 
32'd11765: dataIn1 = 32'd325
; 
32'd11766: dataIn1 = 32'd340
; 
32'd11767: dataIn1 = 32'd374
; 
32'd11768: dataIn1 = 32'd377
; 
32'd11769: dataIn1 = 32'd393
; 
32'd11770: dataIn1 = 32'd305
; 
32'd11771: dataIn1 = 32'd309
; 
32'd11772: dataIn1 = 32'd334
; 
32'd11773: dataIn1 = 32'd341
; 
32'd11774: dataIn1 = 32'd403
; 
32'd11775: dataIn1 = 32'd420
; 
32'd11776: dataIn1 = 32'd262
; 
32'd11777: dataIn1 = 32'd275
; 
32'd11778: dataIn1 = 32'd306
; 
32'd11779: dataIn1 = 32'd342
; 
32'd11780: dataIn1 = 32'd365
; 
32'd11781: dataIn1 = 32'd418
; 
32'd11782: dataIn1 = 32'd420
; 
32'd11783: dataIn1 = 32'd421
; 
32'd11784: dataIn1 = 32'd439
; 
32'd11785: dataIn1 = 32'd247
; 
32'd11786: dataIn1 = 32'd312
; 
32'd11787: dataIn1 = 32'd317
; 
32'd11788: dataIn1 = 32'd343
; 
32'd11789: dataIn1 = 32'd358
; 
32'd11790: dataIn1 = 32'd361
; 
32'd11791: dataIn1 = 32'd422
; 
32'd11792: dataIn1 = 32'd457
; 
32'd11793: dataIn1 = 32'd279
; 
32'd11794: dataIn1 = 32'd285
; 
32'd11795: dataIn1 = 32'd288
; 
32'd11796: dataIn1 = 32'd344
; 
32'd11797: dataIn1 = 32'd353
; 
32'd11798: dataIn1 = 32'd364
; 
32'd11799: dataIn1 = 32'd378
; 
32'd11800: dataIn1 = 32'd264
; 
32'd11801: dataIn1 = 32'd298
; 
32'd11802: dataIn1 = 32'd311
; 
32'd11803: dataIn1 = 32'd345
; 
32'd11804: dataIn1 = 32'd413
; 
32'd11805: dataIn1 = 32'd444
; 
32'd11806: dataIn1 = 32'd253
; 
32'd11807: dataIn1 = 32'd297
; 
32'd11808: dataIn1 = 32'd329
; 
32'd11809: dataIn1 = 32'd346
; 
32'd11810: dataIn1 = 32'd423
; 
32'd11811: dataIn1 = 32'd428
; 
32'd11812: dataIn1 = 32'd432
; 
32'd11813: dataIn1 = 32'd436
; 
32'd11814: dataIn1 = 32'd287
; 
32'd11815: dataIn1 = 32'd293
; 
32'd11816: dataIn1 = 32'd338
; 
32'd11817: dataIn1 = 32'd347
; 
32'd11818: dataIn1 = 32'd402
; 
32'd11819: dataIn1 = 32'd424
; 
32'd11820: dataIn1 = 32'd455
; 
32'd11821: dataIn1 = 32'd251
; 
32'd11822: dataIn1 = 32'd258
; 
32'd11823: dataIn1 = 32'd328
; 
32'd11824: dataIn1 = 32'd348
; 
32'd11825: dataIn1 = 32'd362
; 
32'd11826: dataIn1 = 32'd397
; 
32'd11827: dataIn1 = 32'd405
; 
32'd11828: dataIn1 = 32'd461
; 
32'd11829: dataIn1 = 32'd257
; 
32'd11830: dataIn1 = 32'd266
; 
32'd11831: dataIn1 = 32'd271
; 
32'd11832: dataIn1 = 32'd349
; 
32'd11833: dataIn1 = 32'd356
; 
32'd11834: dataIn1 = 32'd397
; 
32'd11835: dataIn1 = 32'd426
; 
32'd11836: dataIn1 = 32'd270
; 
32'd11837: dataIn1 = 32'd308
; 
32'd11838: dataIn1 = 32'd317
; 
32'd11839: dataIn1 = 32'd350
; 
32'd11840: dataIn1 = 32'd422
; 
32'd11841: dataIn1 = 32'd425
; 
32'd11842: dataIn1 = 32'd257
; 
32'd11843: dataIn1 = 32'd264
; 
32'd11844: dataIn1 = 32'd304
; 
32'd11845: dataIn1 = 32'd351
; 
32'd11846: dataIn1 = 32'd367
; 
32'd11847: dataIn1 = 32'd392
; 
32'd11848: dataIn1 = 32'd426
; 
32'd11849: dataIn1 = 32'd462
; 
32'd11850: dataIn1 = 32'd287
; 
32'd11851: dataIn1 = 32'd316
; 
32'd11852: dataIn1 = 32'd320
; 
32'd11853: dataIn1 = 32'd352
; 
32'd11854: dataIn1 = 32'd384
; 
32'd11855: dataIn1 = 32'd279
; 
32'd11856: dataIn1 = 32'd331
; 
32'd11857: dataIn1 = 32'd344
; 
32'd11858: dataIn1 = 32'd353
; 
32'd11859: dataIn1 = 32'd376
; 
32'd11860: dataIn1 = 32'd386
; 
32'd11861: dataIn1 = 32'd427
; 
32'd11862: dataIn1 = 32'd260
; 
32'd11863: dataIn1 = 32'd280
; 
32'd11864: dataIn1 = 32'd283
; 
32'd11865: dataIn1 = 32'd354
; 
32'd11866: dataIn1 = 32'd399
; 
32'd11867: dataIn1 = 32'd417
; 
32'd11868: dataIn1 = 32'd428
; 
32'd11869: dataIn1 = 32'd247
; 
32'd11870: dataIn1 = 32'd256
; 
32'd11871: dataIn1 = 32'd297
; 
32'd11872: dataIn1 = 32'd355
; 
32'd11873: dataIn1 = 32'd404
; 
32'd11874: dataIn1 = 32'd429
; 
32'd11875: dataIn1 = 32'd443
; 
32'd11876: dataIn1 = 32'd271
; 
32'd11877: dataIn1 = 32'd289
; 
32'd11878: dataIn1 = 32'd349
; 
32'd11879: dataIn1 = 32'd356
; 
32'd11880: dataIn1 = 32'd382
; 
32'd11881: dataIn1 = 32'd390
; 
32'd11882: dataIn1 = 32'd430
; 
32'd11883: dataIn1 = 32'd442
; 
32'd11884: dataIn1 = 32'd453
; 
32'd11885: dataIn1 = 32'd463
; 
32'd11886: dataIn1 = 32'd253
; 
32'd11887: dataIn1 = 32'd313
; 
32'd11888: dataIn1 = 32'd336
; 
32'd11889: dataIn1 = 32'd357
; 
32'd11890: dataIn1 = 32'd375
; 
32'd11891: dataIn1 = 32'd381
; 
32'd11892: dataIn1 = 32'd249
; 
32'd11893: dataIn1 = 32'd327
; 
32'd11894: dataIn1 = 32'd343
; 
32'd11895: dataIn1 = 32'd358
; 
32'd11896: dataIn1 = 32'd393
; 
32'd11897: dataIn1 = 32'd412
; 
32'd11898: dataIn1 = 32'd415
; 
32'd11899: dataIn1 = 32'd422
; 
32'd11900: dataIn1 = 32'd464
; 
32'd11901: dataIn1 = 32'd479
; 
32'd11902: dataIn1 = 32'd241
; 
32'd11903: dataIn1 = 32'd268
; 
32'd11904: dataIn1 = 32'd301
; 
32'd11905: dataIn1 = 32'd359
; 
32'd11906: dataIn1 = 32'd383
; 
32'd11907: dataIn1 = 32'd401
; 
32'd11908: dataIn1 = 32'd435
; 
32'd11909: dataIn1 = 32'd465
; 
32'd11910: dataIn1 = 32'd244
; 
32'd11911: dataIn1 = 32'd285
; 
32'd11912: dataIn1 = 32'd318
; 
32'd11913: dataIn1 = 32'd360
; 
32'd11914: dataIn1 = 32'd378
; 
32'd11915: dataIn1 = 32'd411
; 
32'd11916: dataIn1 = 32'd247
; 
32'd11917: dataIn1 = 32'd314
; 
32'd11918: dataIn1 = 32'd343
; 
32'd11919: dataIn1 = 32'd361
; 
32'd11920: dataIn1 = 32'd404
; 
32'd11921: dataIn1 = 32'd415
; 
32'd11922: dataIn1 = 32'd457
; 
32'd11923: dataIn1 = 32'd258
; 
32'd11924: dataIn1 = 32'd263
; 
32'd11925: dataIn1 = 32'd348
; 
32'd11926: dataIn1 = 32'd362
; 
32'd11927: dataIn1 = 32'd366
; 
32'd11928: dataIn1 = 32'd417
; 
32'd11929: dataIn1 = 32'd447
; 
32'd11930: dataIn1 = 32'd466
; 
32'd11931: dataIn1 = 32'd259
; 
32'd11932: dataIn1 = 32'd277
; 
32'd11933: dataIn1 = 32'd307
; 
32'd11934: dataIn1 = 32'd363
; 
32'd11935: dataIn1 = 32'd373
; 
32'd11936: dataIn1 = 32'd398
; 
32'd11937: dataIn1 = 32'd438
; 
32'd11938: dataIn1 = 32'd260
; 
32'd11939: dataIn1 = 32'd263
; 
32'd11940: dataIn1 = 32'd344
; 
32'd11941: dataIn1 = 32'd364
; 
32'd11942: dataIn1 = 32'd399
; 
32'd11943: dataIn1 = 32'd262
; 
32'd11944: dataIn1 = 32'd322
; 
32'd11945: dataIn1 = 32'd342
; 
32'd11946: dataIn1 = 32'd365
; 
32'd11947: dataIn1 = 32'd431
; 
32'd11948: dataIn1 = 32'd439
; 
32'd11949: dataIn1 = 32'd263
; 
32'd11950: dataIn1 = 32'd321
; 
32'd11951: dataIn1 = 32'd362
; 
32'd11952: dataIn1 = 32'd366
; 
32'd11953: dataIn1 = 32'd419
; 
32'd11954: dataIn1 = 32'd264
; 
32'd11955: dataIn1 = 32'd328
; 
32'd11956: dataIn1 = 32'd351
; 
32'd11957: dataIn1 = 32'd367
; 
32'd11958: dataIn1 = 32'd392
; 
32'd11959: dataIn1 = 32'd405
; 
32'd11960: dataIn1 = 32'd462
; 
32'd11961: dataIn1 = 32'd475
; 
32'd11962: dataIn1 = 32'd266
; 
32'd11963: dataIn1 = 32'd313
; 
32'd11964: dataIn1 = 32'd324
; 
32'd11965: dataIn1 = 32'd368
; 
32'd11966: dataIn1 = 32'd395
; 
32'd11967: dataIn1 = 32'd430
; 
32'd11968: dataIn1 = 32'd268
; 
32'd11969: dataIn1 = 32'd306
; 
32'd11970: dataIn1 = 32'd335
; 
32'd11971: dataIn1 = 32'd369
; 
32'd11972: dataIn1 = 32'd383
; 
32'd11973: dataIn1 = 32'd421
; 
32'd11974: dataIn1 = 32'd269
; 
32'd11975: dataIn1 = 32'd275
; 
32'd11976: dataIn1 = 32'd299
; 
32'd11977: dataIn1 = 32'd370
; 
32'd11978: dataIn1 = 32'd372
; 
32'd11979: dataIn1 = 32'd416
; 
32'd11980: dataIn1 = 32'd446
; 
32'd11981: dataIn1 = 32'd268
; 
32'd11982: dataIn1 = 32'd272
; 
32'd11983: dataIn1 = 32'd295
; 
32'd11984: dataIn1 = 32'd371
; 
32'd11985: dataIn1 = 32'd421
; 
32'd11986: dataIn1 = 32'd425
; 
32'd11987: dataIn1 = 32'd435
; 
32'd11988: dataIn1 = 32'd437
; 
32'd11989: dataIn1 = 32'd275
; 
32'd11990: dataIn1 = 32'd322
; 
32'd11991: dataIn1 = 32'd370
; 
32'd11992: dataIn1 = 32'd372
; 
32'd11993: dataIn1 = 32'd379
; 
32'd11994: dataIn1 = 32'd416
; 
32'd11995: dataIn1 = 32'd418
; 
32'd11996: dataIn1 = 32'd439
; 
32'd11997: dataIn1 = 32'd446
; 
32'd11998: dataIn1 = 32'd277
; 
32'd11999: dataIn1 = 32'd319
; 
32'd12000: dataIn1 = 32'd363
; 
32'd12001: dataIn1 = 32'd373
; 
32'd12002: dataIn1 = 32'd424
; 
32'd12003: dataIn1 = 32'd295
; 
32'd12004: dataIn1 = 32'd303
; 
32'd12005: dataIn1 = 32'd340
; 
32'd12006: dataIn1 = 32'd374
; 
32'd12007: dataIn1 = 32'd377
; 
32'd12008: dataIn1 = 32'd391
; 
32'd12009: dataIn1 = 32'd400
; 
32'd12010: dataIn1 = 32'd269
; 
32'd12011: dataIn1 = 32'd299
; 
32'd12012: dataIn1 = 32'd357
; 
32'd12013: dataIn1 = 32'd375
; 
32'd12014: dataIn1 = 32'd396
; 
32'd12015: dataIn1 = 32'd432
; 
32'd12016: dataIn1 = 32'd445
; 
32'd12017: dataIn1 = 32'd489
; 
32'd12018: dataIn1 = 32'd263
; 
32'd12019: dataIn1 = 32'd338
; 
32'd12020: dataIn1 = 32'd353
; 
32'd12021: dataIn1 = 32'd376
; 
32'd12022: dataIn1 = 32'd386
; 
32'd12023: dataIn1 = 32'd447
; 
32'd12024: dataIn1 = 32'd468
; 
32'd12025: dataIn1 = 32'd488
; 
32'd12026: dataIn1 = 32'd295
; 
32'd12027: dataIn1 = 32'd340
; 
32'd12028: dataIn1 = 32'd374
; 
32'd12029: dataIn1 = 32'd377
; 
32'd12030: dataIn1 = 32'd391
; 
32'd12031: dataIn1 = 32'd437
; 
32'd12032: dataIn1 = 32'd467
; 
32'd12033: dataIn1 = 32'd472
; 
32'd12034: dataIn1 = 32'd285
; 
32'd12035: dataIn1 = 32'd344
; 
32'd12036: dataIn1 = 32'd360
; 
32'd12037: dataIn1 = 32'd378
; 
32'd12038: dataIn1 = 32'd427
; 
32'd12039: dataIn1 = 32'd468
; 
32'd12040: dataIn1 = 32'd322
; 
32'd12041: dataIn1 = 32'd330
; 
32'd12042: dataIn1 = 32'd372
; 
32'd12043: dataIn1 = 32'd379
; 
32'd12044: dataIn1 = 32'd452
; 
32'd12045: dataIn1 = 32'd456
; 
32'd12046: dataIn1 = 32'd486
; 
32'd12047: dataIn1 = 32'd324
; 
32'd12048: dataIn1 = 32'd330
; 
32'd12049: dataIn1 = 32'd339
; 
32'd12050: dataIn1 = 32'd380
; 
32'd12051: dataIn1 = 32'd382
; 
32'd12052: dataIn1 = 32'd395
; 
32'd12053: dataIn1 = 32'd450
; 
32'd12054: dataIn1 = 32'd453
; 
32'd12055: dataIn1 = 32'd333
; 
32'd12056: dataIn1 = 32'd336
; 
32'd12057: dataIn1 = 32'd357
; 
32'd12058: dataIn1 = 32'd381
; 
32'd12059: dataIn1 = 32'd432
; 
32'd12060: dataIn1 = 32'd440
; 
32'd12061: dataIn1 = 32'd339
; 
32'd12062: dataIn1 = 32'd356
; 
32'd12063: dataIn1 = 32'd380
; 
32'd12064: dataIn1 = 32'd382
; 
32'd12065: dataIn1 = 32'd398
; 
32'd12066: dataIn1 = 32'd450
; 
32'd12067: dataIn1 = 32'd453
; 
32'd12068: dataIn1 = 32'd315
; 
32'd12069: dataIn1 = 32'd359
; 
32'd12070: dataIn1 = 32'd369
; 
32'd12071: dataIn1 = 32'd383
; 
32'd12072: dataIn1 = 32'd435
; 
32'd12073: dataIn1 = 32'd458
; 
32'd12074: dataIn1 = 32'd504
; 
32'd12075: dataIn1 = 32'd518
; 
32'd12076: dataIn1 = 32'd320
; 
32'd12077: dataIn1 = 32'd337
; 
32'd12078: dataIn1 = 32'd352
; 
32'd12079: dataIn1 = 32'd384
; 
32'd12080: dataIn1 = 32'd419
; 
32'd12081: dataIn1 = 32'd469
; 
32'd12082: dataIn1 = 32'd301
; 
32'd12083: dataIn1 = 32'd307
; 
32'd12084: dataIn1 = 32'd332
; 
32'd12085: dataIn1 = 32'd385
; 
32'd12086: dataIn1 = 32'd387
; 
32'd12087: dataIn1 = 32'd394
; 
32'd12088: dataIn1 = 32'd434
; 
32'd12089: dataIn1 = 32'd438
; 
32'd12090: dataIn1 = 32'd442
; 
32'd12091: dataIn1 = 32'd338
; 
32'd12092: dataIn1 = 32'd353
; 
32'd12093: dataIn1 = 32'd376
; 
32'd12094: dataIn1 = 32'd386
; 
32'd12095: dataIn1 = 32'd433
; 
32'd12096: dataIn1 = 32'd469
; 
32'd12097: dataIn1 = 32'd488
; 
32'd12098: dataIn1 = 32'd499
; 
32'd12099: dataIn1 = 32'd301
; 
32'd12100: dataIn1 = 32'd332
; 
32'd12101: dataIn1 = 32'd385
; 
32'd12102: dataIn1 = 32'd387
; 
32'd12103: dataIn1 = 32'd390
; 
32'd12104: dataIn1 = 32'd401
; 
32'd12105: dataIn1 = 32'd269
; 
32'd12106: dataIn1 = 32'd323
; 
32'd12107: dataIn1 = 32'd329
; 
32'd12108: dataIn1 = 32'd388
; 
32'd12109: dataIn1 = 32'd406
; 
32'd12110: dataIn1 = 32'd436
; 
32'd12111: dataIn1 = 32'd247
; 
32'd12112: dataIn1 = 32'd300
; 
32'd12113: dataIn1 = 32'd310
; 
32'd12114: dataIn1 = 32'd389
; 
32'd12115: dataIn1 = 32'd403
; 
32'd12116: dataIn1 = 32'd409
; 
32'd12117: dataIn1 = 32'd443
; 
32'd12118: dataIn1 = 32'd470
; 
32'd12119: dataIn1 = 32'd332
; 
32'd12120: dataIn1 = 32'd356
; 
32'd12121: dataIn1 = 32'd387
; 
32'd12122: dataIn1 = 32'd390
; 
32'd12123: dataIn1 = 32'd426
; 
32'd12124: dataIn1 = 32'd434
; 
32'd12125: dataIn1 = 32'd463
; 
32'd12126: dataIn1 = 32'd471
; 
32'd12127: dataIn1 = 32'd295
; 
32'd12128: dataIn1 = 32'd374
; 
32'd12129: dataIn1 = 32'd377
; 
32'd12130: dataIn1 = 32'd391
; 
32'd12131: dataIn1 = 32'd394
; 
32'd12132: dataIn1 = 32'd315
; 
32'd12133: dataIn1 = 32'd351
; 
32'd12134: dataIn1 = 32'd367
; 
32'd12135: dataIn1 = 32'd392
; 
32'd12136: dataIn1 = 32'd471
; 
32'd12137: dataIn1 = 32'd497
; 
32'd12138: dataIn1 = 32'd498
; 
32'd12139: dataIn1 = 32'd527
; 
32'd12140: dataIn1 = 32'd320
; 
32'd12141: dataIn1 = 32'd340
; 
32'd12142: dataIn1 = 32'd358
; 
32'd12143: dataIn1 = 32'd393
; 
32'd12144: dataIn1 = 32'd400
; 
32'd12145: dataIn1 = 32'd467
; 
32'd12146: dataIn1 = 32'd301
; 
32'd12147: dataIn1 = 32'd385
; 
32'd12148: dataIn1 = 32'd391
; 
32'd12149: dataIn1 = 32'd394
; 
32'd12150: dataIn1 = 32'd402
; 
32'd12151: dataIn1 = 32'd438
; 
32'd12152: dataIn1 = 32'd455
; 
32'd12153: dataIn1 = 32'd465
; 
32'd12154: dataIn1 = 32'd472
; 
32'd12155: dataIn1 = 32'd485
; 
32'd12156: dataIn1 = 32'd487
; 
32'd12157: dataIn1 = 32'd313
; 
32'd12158: dataIn1 = 32'd368
; 
32'd12159: dataIn1 = 32'd380
; 
32'd12160: dataIn1 = 32'd395
; 
32'd12161: dataIn1 = 32'd445
; 
32'd12162: dataIn1 = 32'd482
; 
32'd12163: dataIn1 = 32'd299
; 
32'd12164: dataIn1 = 32'd330
; 
32'd12165: dataIn1 = 32'd375
; 
32'd12166: dataIn1 = 32'd396
; 
32'd12167: dataIn1 = 32'd333
; 
32'd12168: dataIn1 = 32'd348
; 
32'd12169: dataIn1 = 32'd349
; 
32'd12170: dataIn1 = 32'd397
; 
32'd12171: dataIn1 = 32'd430
; 
32'd12172: dataIn1 = 32'd462
; 
32'd12173: dataIn1 = 32'd466
; 
32'd12174: dataIn1 = 32'd483
; 
32'd12175: dataIn1 = 32'd490
; 
32'd12176: dataIn1 = 32'd546
; 
32'd12177: dataIn1 = 32'd339
; 
32'd12178: dataIn1 = 32'd363
; 
32'd12179: dataIn1 = 32'd382
; 
32'd12180: dataIn1 = 32'd398
; 
32'd12181: dataIn1 = 32'd410
; 
32'd12182: dataIn1 = 32'd318
; 
32'd12183: dataIn1 = 32'd354
; 
32'd12184: dataIn1 = 32'd364
; 
32'd12185: dataIn1 = 32'd399
; 
32'd12186: dataIn1 = 32'd407
; 
32'd12187: dataIn1 = 32'd441
; 
32'd12188: dataIn1 = 32'd451
; 
32'd12189: dataIn1 = 32'd495
; 
32'd12190: dataIn1 = 32'd320
; 
32'd12191: dataIn1 = 32'd374
; 
32'd12192: dataIn1 = 32'd393
; 
32'd12193: dataIn1 = 32'd400
; 
32'd12194: dataIn1 = 32'd469
; 
32'd12195: dataIn1 = 32'd301
; 
32'd12196: dataIn1 = 32'd359
; 
32'd12197: dataIn1 = 32'd387
; 
32'd12198: dataIn1 = 32'd401
; 
32'd12199: dataIn1 = 32'd434
; 
32'd12200: dataIn1 = 32'd458
; 
32'd12201: dataIn1 = 32'd494
; 
32'd12202: dataIn1 = 32'd307
; 
32'd12203: dataIn1 = 32'd347
; 
32'd12204: dataIn1 = 32'd394
; 
32'd12205: dataIn1 = 32'd402
; 
32'd12206: dataIn1 = 32'd424
; 
32'd12207: dataIn1 = 32'd455
; 
32'd12208: dataIn1 = 32'd310
; 
32'd12209: dataIn1 = 32'd341
; 
32'd12210: dataIn1 = 32'd389
; 
32'd12211: dataIn1 = 32'd403
; 
32'd12212: dataIn1 = 32'd409
; 
32'd12213: dataIn1 = 32'd411
; 
32'd12214: dataIn1 = 32'd420
; 
32'd12215: dataIn1 = 32'd448
; 
32'd12216: dataIn1 = 32'd449
; 
32'd12217: dataIn1 = 32'd470
; 
32'd12218: dataIn1 = 32'd473
; 
32'd12219: dataIn1 = 32'd493
; 
32'd12220: dataIn1 = 32'd505
; 
32'd12221: dataIn1 = 32'd547
; 
32'd12222: dataIn1 = 32'd569
; 
32'd12223: dataIn1 = 32'd571
; 
32'd12224: dataIn1 = 32'd247
; 
32'd12225: dataIn1 = 32'd355
; 
32'd12226: dataIn1 = 32'd361
; 
32'd12227: dataIn1 = 32'd404
; 
32'd12228: dataIn1 = 32'd408
; 
32'd12229: dataIn1 = 32'd423
; 
32'd12230: dataIn1 = 32'd454
; 
32'd12231: dataIn1 = 32'd459
; 
32'd12232: dataIn1 = 32'd474
; 
32'd12233: dataIn1 = 32'd506
; 
32'd12234: dataIn1 = 32'd311
; 
32'd12235: dataIn1 = 32'd348
; 
32'd12236: dataIn1 = 32'd367
; 
32'd12237: dataIn1 = 32'd405
; 
32'd12238: dataIn1 = 32'd461
; 
32'd12239: dataIn1 = 32'd475
; 
32'd12240: dataIn1 = 32'd269
; 
32'd12241: dataIn1 = 32'd335
; 
32'd12242: dataIn1 = 32'd388
; 
32'd12243: dataIn1 = 32'd406
; 
32'd12244: dataIn1 = 32'd414
; 
32'd12245: dataIn1 = 32'd459
; 
32'd12246: dataIn1 = 32'd489
; 
32'd12247: dataIn1 = 32'd507
; 
32'd12248: dataIn1 = 32'd297
; 
32'd12249: dataIn1 = 32'd318
; 
32'd12250: dataIn1 = 32'd399
; 
32'd12251: dataIn1 = 32'd407
; 
32'd12252: dataIn1 = 32'd441
; 
32'd12253: dataIn1 = 32'd443
; 
32'd12254: dataIn1 = 32'd449
; 
32'd12255: dataIn1 = 32'd451
; 
32'd12256: dataIn1 = 32'd508
; 
32'd12257: dataIn1 = 32'd298
; 
32'd12258: dataIn1 = 32'd327
; 
32'd12259: dataIn1 = 32'd404
; 
32'd12260: dataIn1 = 32'd408
; 
32'd12261: dataIn1 = 32'd413
; 
32'd12262: dataIn1 = 32'd444
; 
32'd12263: dataIn1 = 32'd474
; 
32'd12264: dataIn1 = 32'd476
; 
32'd12265: dataIn1 = 32'd300
; 
32'd12266: dataIn1 = 32'd389
; 
32'd12267: dataIn1 = 32'd403
; 
32'd12268: dataIn1 = 32'd409
; 
32'd12269: dataIn1 = 32'd302
; 
32'd12270: dataIn1 = 32'd331
; 
32'd12271: dataIn1 = 32'd398
; 
32'd12272: dataIn1 = 32'd410
; 
32'd12273: dataIn1 = 32'd431
; 
32'd12274: dataIn1 = 32'd433
; 
32'd12275: dataIn1 = 32'd450
; 
32'd12276: dataIn1 = 32'd480
; 
32'd12277: dataIn1 = 32'd509
; 
32'd12278: dataIn1 = 32'd309
; 
32'd12279: dataIn1 = 32'd360
; 
32'd12280: dataIn1 = 32'd403
; 
32'd12281: dataIn1 = 32'd411
; 
32'd12282: dataIn1 = 32'd441
; 
32'd12283: dataIn1 = 32'd448
; 
32'd12284: dataIn1 = 32'd449
; 
32'd12285: dataIn1 = 32'd501
; 
32'd12286: dataIn1 = 32'd311
; 
32'd12287: dataIn1 = 32'd327
; 
32'd12288: dataIn1 = 32'd358
; 
32'd12289: dataIn1 = 32'd412
; 
32'd12290: dataIn1 = 32'd444
; 
32'd12291: dataIn1 = 32'd464
; 
32'd12292: dataIn1 = 32'd492
; 
32'd12293: dataIn1 = 32'd315
; 
32'd12294: dataIn1 = 32'd345
; 
32'd12295: dataIn1 = 32'd408
; 
32'd12296: dataIn1 = 32'd413
; 
32'd12297: dataIn1 = 32'd476
; 
32'd12298: dataIn1 = 32'd315
; 
32'd12299: dataIn1 = 32'd323
; 
32'd12300: dataIn1 = 32'd406
; 
32'd12301: dataIn1 = 32'd414
; 
32'd12302: dataIn1 = 32'd510
; 
32'd12303: dataIn1 = 32'd517
; 
32'd12304: dataIn1 = 32'd327
; 
32'd12305: dataIn1 = 32'd358
; 
32'd12306: dataIn1 = 32'd361
; 
32'd12307: dataIn1 = 32'd415
; 
32'd12308: dataIn1 = 32'd457
; 
32'd12309: dataIn1 = 32'd474
; 
32'd12310: dataIn1 = 32'd330
; 
32'd12311: dataIn1 = 32'd370
; 
32'd12312: dataIn1 = 32'd372
; 
32'd12313: dataIn1 = 32'd416
; 
32'd12314: dataIn1 = 32'd452
; 
32'd12315: dataIn1 = 32'd477
; 
32'd12316: dataIn1 = 32'd333
; 
32'd12317: dataIn1 = 32'd354
; 
32'd12318: dataIn1 = 32'd362
; 
32'd12319: dataIn1 = 32'd417
; 
32'd12320: dataIn1 = 32'd440
; 
32'd12321: dataIn1 = 32'd466
; 
32'd12322: dataIn1 = 32'd521
; 
32'd12323: dataIn1 = 32'd548
; 
32'd12324: dataIn1 = 32'd335
; 
32'd12325: dataIn1 = 32'd342
; 
32'd12326: dataIn1 = 32'd372
; 
32'd12327: dataIn1 = 32'd418
; 
32'd12328: dataIn1 = 32'd446
; 
32'd12329: dataIn1 = 32'd460
; 
32'd12330: dataIn1 = 32'd337
; 
32'd12331: dataIn1 = 32'd366
; 
32'd12332: dataIn1 = 32'd384
; 
32'd12333: dataIn1 = 32'd419
; 
32'd12334: dataIn1 = 32'd447
; 
32'd12335: dataIn1 = 32'd461
; 
32'd12336: dataIn1 = 32'd478
; 
32'd12337: dataIn1 = 32'd500
; 
32'd12338: dataIn1 = 32'd341
; 
32'd12339: dataIn1 = 32'd342
; 
32'd12340: dataIn1 = 32'd403
; 
32'd12341: dataIn1 = 32'd420
; 
32'd12342: dataIn1 = 32'd425
; 
32'd12343: dataIn1 = 32'd484
; 
32'd12344: dataIn1 = 32'd493
; 
32'd12345: dataIn1 = 32'd511
; 
32'd12346: dataIn1 = 32'd532
; 
32'd12347: dataIn1 = 32'd342
; 
32'd12348: dataIn1 = 32'd369
; 
32'd12349: dataIn1 = 32'd371
; 
32'd12350: dataIn1 = 32'd421
; 
32'd12351: dataIn1 = 32'd460
; 
32'd12352: dataIn1 = 32'd484
; 
32'd12353: dataIn1 = 32'd512
; 
32'd12354: dataIn1 = 32'd518
; 
32'd12355: dataIn1 = 32'd343
; 
32'd12356: dataIn1 = 32'd350
; 
32'd12357: dataIn1 = 32'd358
; 
32'd12358: dataIn1 = 32'd422
; 
32'd12359: dataIn1 = 32'd467
; 
32'd12360: dataIn1 = 32'd470
; 
32'd12361: dataIn1 = 32'd479
; 
32'd12362: dataIn1 = 32'd256
; 
32'd12363: dataIn1 = 32'd346
; 
32'd12364: dataIn1 = 32'd404
; 
32'd12365: dataIn1 = 32'd423
; 
32'd12366: dataIn1 = 32'd429
; 
32'd12367: dataIn1 = 32'd436
; 
32'd12368: dataIn1 = 32'd347
; 
32'd12369: dataIn1 = 32'd373
; 
32'd12370: dataIn1 = 32'd402
; 
32'd12371: dataIn1 = 32'd424
; 
32'd12372: dataIn1 = 32'd433
; 
32'd12373: dataIn1 = 32'd350
; 
32'd12374: dataIn1 = 32'd371
; 
32'd12375: dataIn1 = 32'd420
; 
32'd12376: dataIn1 = 32'd425
; 
32'd12377: dataIn1 = 32'd484
; 
32'd12378: dataIn1 = 32'd493
; 
32'd12379: dataIn1 = 32'd535
; 
32'd12380: dataIn1 = 32'd349
; 
32'd12381: dataIn1 = 32'd351
; 
32'd12382: dataIn1 = 32'd390
; 
32'd12383: dataIn1 = 32'd426
; 
32'd12384: dataIn1 = 32'd463
; 
32'd12385: dataIn1 = 32'd471
; 
32'd12386: dataIn1 = 32'd331
; 
32'd12387: dataIn1 = 32'd353
; 
32'd12388: dataIn1 = 32'd378
; 
32'd12389: dataIn1 = 32'd427
; 
32'd12390: dataIn1 = 32'd480
; 
32'd12391: dataIn1 = 32'd297
; 
32'd12392: dataIn1 = 32'd346
; 
32'd12393: dataIn1 = 32'd354
; 
32'd12394: dataIn1 = 32'd428
; 
32'd12395: dataIn1 = 32'd451
; 
32'd12396: dataIn1 = 32'd481
; 
32'd12397: dataIn1 = 32'd297
; 
32'd12398: dataIn1 = 32'd355
; 
32'd12399: dataIn1 = 32'd423
; 
32'd12400: dataIn1 = 32'd429
; 
32'd12401: dataIn1 = 32'd454
; 
32'd12402: dataIn1 = 32'd356
; 
32'd12403: dataIn1 = 32'd368
; 
32'd12404: dataIn1 = 32'd397
; 
32'd12405: dataIn1 = 32'd430
; 
32'd12406: dataIn1 = 32'd483
; 
32'd12407: dataIn1 = 32'd549
; 
32'd12408: dataIn1 = 32'd563
; 
32'd12409: dataIn1 = 32'd302
; 
32'd12410: dataIn1 = 32'd365
; 
32'd12411: dataIn1 = 32'd410
; 
32'd12412: dataIn1 = 32'd431
; 
32'd12413: dataIn1 = 32'd473
; 
32'd12414: dataIn1 = 32'd486
; 
32'd12415: dataIn1 = 32'd346
; 
32'd12416: dataIn1 = 32'd375
; 
32'd12417: dataIn1 = 32'd381
; 
32'd12418: dataIn1 = 32'd432
; 
32'd12419: dataIn1 = 32'd445
; 
32'd12420: dataIn1 = 32'd481
; 
32'd12421: dataIn1 = 32'd491
; 
32'd12422: dataIn1 = 32'd502
; 
32'd12423: dataIn1 = 32'd386
; 
32'd12424: dataIn1 = 32'd410
; 
32'd12425: dataIn1 = 32'd424
; 
32'd12426: dataIn1 = 32'd433
; 
32'd12427: dataIn1 = 32'd385
; 
32'd12428: dataIn1 = 32'd390
; 
32'd12429: dataIn1 = 32'd401
; 
32'd12430: dataIn1 = 32'd434
; 
32'd12431: dataIn1 = 32'd465
; 
32'd12432: dataIn1 = 32'd485
; 
32'd12433: dataIn1 = 32'd494
; 
32'd12434: dataIn1 = 32'd359
; 
32'd12435: dataIn1 = 32'd371
; 
32'd12436: dataIn1 = 32'd383
; 
32'd12437: dataIn1 = 32'd435
; 
32'd12438: dataIn1 = 32'd437
; 
32'd12439: dataIn1 = 32'd504
; 
32'd12440: dataIn1 = 32'd346
; 
32'd12441: dataIn1 = 32'd388
; 
32'd12442: dataIn1 = 32'd423
; 
32'd12443: dataIn1 = 32'd436
; 
32'd12444: dataIn1 = 32'd481
; 
32'd12445: dataIn1 = 32'd491
; 
32'd12446: dataIn1 = 32'd371
; 
32'd12447: dataIn1 = 32'd377
; 
32'd12448: dataIn1 = 32'd435
; 
32'd12449: dataIn1 = 32'd437
; 
32'd12450: dataIn1 = 32'd472
; 
32'd12451: dataIn1 = 32'd520
; 
32'd12452: dataIn1 = 32'd531
; 
32'd12453: dataIn1 = 32'd363
; 
32'd12454: dataIn1 = 32'd385
; 
32'd12455: dataIn1 = 32'd394
; 
32'd12456: dataIn1 = 32'd438
; 
32'd12457: dataIn1 = 32'd442
; 
32'd12458: dataIn1 = 32'd485
; 
32'd12459: dataIn1 = 32'd487
; 
32'd12460: dataIn1 = 32'd509
; 
32'd12461: dataIn1 = 32'd342
; 
32'd12462: dataIn1 = 32'd365
; 
32'd12463: dataIn1 = 32'd372
; 
32'd12464: dataIn1 = 32'd439
; 
32'd12465: dataIn1 = 32'd456
; 
32'd12466: dataIn1 = 32'd511
; 
32'd12467: dataIn1 = 32'd512
; 
32'd12468: dataIn1 = 32'd333
; 
32'd12469: dataIn1 = 32'd381
; 
32'd12470: dataIn1 = 32'd417
; 
32'd12471: dataIn1 = 32'd440
; 
32'd12472: dataIn1 = 32'd483
; 
32'd12473: dataIn1 = 32'd399
; 
32'd12474: dataIn1 = 32'd407
; 
32'd12475: dataIn1 = 32'd411
; 
32'd12476: dataIn1 = 32'd441
; 
32'd12477: dataIn1 = 32'd513
; 
32'd12478: dataIn1 = 32'd536
; 
32'd12479: dataIn1 = 32'd356
; 
32'd12480: dataIn1 = 32'd385
; 
32'd12481: dataIn1 = 32'd438
; 
32'd12482: dataIn1 = 32'd442
; 
32'd12483: dataIn1 = 32'd514
; 
32'd12484: dataIn1 = 32'd355
; 
32'd12485: dataIn1 = 32'd389
; 
32'd12486: dataIn1 = 32'd407
; 
32'd12487: dataIn1 = 32'd443
; 
32'd12488: dataIn1 = 32'd454
; 
32'd12489: dataIn1 = 32'd503
; 
32'd12490: dataIn1 = 32'd505
; 
32'd12491: dataIn1 = 32'd345
; 
32'd12492: dataIn1 = 32'd408
; 
32'd12493: dataIn1 = 32'd412
; 
32'd12494: dataIn1 = 32'd444
; 
32'd12495: dataIn1 = 32'd497
; 
32'd12496: dataIn1 = 32'd519
; 
32'd12497: dataIn1 = 32'd375
; 
32'd12498: dataIn1 = 32'd395
; 
32'd12499: dataIn1 = 32'd432
; 
32'd12500: dataIn1 = 32'd445
; 
32'd12501: dataIn1 = 32'd477
; 
32'd12502: dataIn1 = 32'd482
; 
32'd12503: dataIn1 = 32'd550
; 
32'd12504: dataIn1 = 32'd559
; 
32'd12505: dataIn1 = 32'd370
; 
32'd12506: dataIn1 = 32'd372
; 
32'd12507: dataIn1 = 32'd418
; 
32'd12508: dataIn1 = 32'd446
; 
32'd12509: dataIn1 = 32'd456
; 
32'd12510: dataIn1 = 32'd477
; 
32'd12511: dataIn1 = 32'd496
; 
32'd12512: dataIn1 = 32'd362
; 
32'd12513: dataIn1 = 32'd376
; 
32'd12514: dataIn1 = 32'd419
; 
32'd12515: dataIn1 = 32'd447
; 
32'd12516: dataIn1 = 32'd468
; 
32'd12517: dataIn1 = 32'd495
; 
32'd12518: dataIn1 = 32'd541
; 
32'd12519: dataIn1 = 32'd544
; 
32'd12520: dataIn1 = 32'd551
; 
32'd12521: dataIn1 = 32'd309
; 
32'd12522: dataIn1 = 32'd403
; 
32'd12523: dataIn1 = 32'd411
; 
32'd12524: dataIn1 = 32'd448
; 
32'd12525: dataIn1 = 32'd473
; 
32'd12526: dataIn1 = 32'd480
; 
32'd12527: dataIn1 = 32'd501
; 
32'd12528: dataIn1 = 32'd403
; 
32'd12529: dataIn1 = 32'd407
; 
32'd12530: dataIn1 = 32'd411
; 
32'd12531: dataIn1 = 32'd449
; 
32'd12532: dataIn1 = 32'd501
; 
32'd12533: dataIn1 = 32'd515
; 
32'd12534: dataIn1 = 32'd380
; 
32'd12535: dataIn1 = 32'd382
; 
32'd12536: dataIn1 = 32'd410
; 
32'd12537: dataIn1 = 32'd450
; 
32'd12538: dataIn1 = 32'd486
; 
32'd12539: dataIn1 = 32'd509
; 
32'd12540: dataIn1 = 32'd538
; 
32'd12541: dataIn1 = 32'd399
; 
32'd12542: dataIn1 = 32'd407
; 
32'd12543: dataIn1 = 32'd428
; 
32'd12544: dataIn1 = 32'd451
; 
32'd12545: dataIn1 = 32'd502
; 
32'd12546: dataIn1 = 32'd515
; 
32'd12547: dataIn1 = 32'd330
; 
32'd12548: dataIn1 = 32'd379
; 
32'd12549: dataIn1 = 32'd416
; 
32'd12550: dataIn1 = 32'd452
; 
32'd12551: dataIn1 = 32'd482
; 
32'd12552: dataIn1 = 32'd356
; 
32'd12553: dataIn1 = 32'd380
; 
32'd12554: dataIn1 = 32'd382
; 
32'd12555: dataIn1 = 32'd453
; 
32'd12556: dataIn1 = 32'd514
; 
32'd12557: dataIn1 = 32'd549
; 
32'd12558: dataIn1 = 32'd404
; 
32'd12559: dataIn1 = 32'd429
; 
32'd12560: dataIn1 = 32'd443
; 
32'd12561: dataIn1 = 32'd454
; 
32'd12562: dataIn1 = 32'd508
; 
32'd12563: dataIn1 = 32'd540
; 
32'd12564: dataIn1 = 32'd566
; 
32'd12565: dataIn1 = 32'd347
; 
32'd12566: dataIn1 = 32'd394
; 
32'd12567: dataIn1 = 32'd402
; 
32'd12568: dataIn1 = 32'd455
; 
32'd12569: dataIn1 = 32'd379
; 
32'd12570: dataIn1 = 32'd439
; 
32'd12571: dataIn1 = 32'd446
; 
32'd12572: dataIn1 = 32'd456
; 
32'd12573: dataIn1 = 32'd516
; 
32'd12574: dataIn1 = 32'd525
; 
32'd12575: dataIn1 = 32'd530
; 
32'd12576: dataIn1 = 32'd343
; 
32'd12577: dataIn1 = 32'd361
; 
32'd12578: dataIn1 = 32'd415
; 
32'd12579: dataIn1 = 32'd457
; 
32'd12580: dataIn1 = 32'd479
; 
32'd12581: dataIn1 = 32'd503
; 
32'd12582: dataIn1 = 32'd315
; 
32'd12583: dataIn1 = 32'd383
; 
32'd12584: dataIn1 = 32'd401
; 
32'd12585: dataIn1 = 32'd458
; 
32'd12586: dataIn1 = 32'd510
; 
32'd12587: dataIn1 = 32'd517
; 
32'd12588: dataIn1 = 32'd526
; 
32'd12589: dataIn1 = 32'd542
; 
32'd12590: dataIn1 = 32'd576
; 
32'd12591: dataIn1 = 32'd580
; 
32'd12592: dataIn1 = 32'd588
; 
32'd12593: dataIn1 = 32'd323
; 
32'd12594: dataIn1 = 32'd404
; 
32'd12595: dataIn1 = 32'd406
; 
32'd12596: dataIn1 = 32'd459
; 
32'd12597: dataIn1 = 32'd476
; 
32'd12598: dataIn1 = 32'd506
; 
32'd12599: dataIn1 = 32'd507
; 
32'd12600: dataIn1 = 32'd537
; 
32'd12601: dataIn1 = 32'd558
; 
32'd12602: dataIn1 = 32'd598
; 
32'd12603: dataIn1 = 32'd335
; 
32'd12604: dataIn1 = 32'd418
; 
32'd12605: dataIn1 = 32'd421
; 
32'd12606: dataIn1 = 32'd460
; 
32'd12607: dataIn1 = 32'd507
; 
32'd12608: dataIn1 = 32'd510
; 
32'd12609: dataIn1 = 32'd512
; 
32'd12610: dataIn1 = 32'd518
; 
32'd12611: dataIn1 = 32'd552
; 
32'd12612: dataIn1 = 32'd348
; 
32'd12613: dataIn1 = 32'd405
; 
32'd12614: dataIn1 = 32'd419
; 
32'd12615: dataIn1 = 32'd461
; 
32'd12616: dataIn1 = 32'd475
; 
32'd12617: dataIn1 = 32'd519
; 
32'd12618: dataIn1 = 32'd534
; 
32'd12619: dataIn1 = 32'd544
; 
32'd12620: dataIn1 = 32'd546
; 
32'd12621: dataIn1 = 32'd351
; 
32'd12622: dataIn1 = 32'd367
; 
32'd12623: dataIn1 = 32'd397
; 
32'd12624: dataIn1 = 32'd462
; 
32'd12625: dataIn1 = 32'd490
; 
32'd12626: dataIn1 = 32'd356
; 
32'd12627: dataIn1 = 32'd390
; 
32'd12628: dataIn1 = 32'd426
; 
32'd12629: dataIn1 = 32'd463
; 
32'd12630: dataIn1 = 32'd490
; 
32'd12631: dataIn1 = 32'd514
; 
32'd12632: dataIn1 = 32'd337
; 
32'd12633: dataIn1 = 32'd358
; 
32'd12634: dataIn1 = 32'd412
; 
32'd12635: dataIn1 = 32'd464
; 
32'd12636: dataIn1 = 32'd478
; 
32'd12637: dataIn1 = 32'd492
; 
32'd12638: dataIn1 = 32'd534
; 
32'd12639: dataIn1 = 32'd359
; 
32'd12640: dataIn1 = 32'd394
; 
32'd12641: dataIn1 = 32'd434
; 
32'd12642: dataIn1 = 32'd465
; 
32'd12643: dataIn1 = 32'd504
; 
32'd12644: dataIn1 = 32'd520
; 
32'd12645: dataIn1 = 32'd533
; 
32'd12646: dataIn1 = 32'd362
; 
32'd12647: dataIn1 = 32'd397
; 
32'd12648: dataIn1 = 32'd417
; 
32'd12649: dataIn1 = 32'd466
; 
32'd12650: dataIn1 = 32'd521
; 
32'd12651: dataIn1 = 32'd544
; 
32'd12652: dataIn1 = 32'd553
; 
32'd12653: dataIn1 = 32'd377
; 
32'd12654: dataIn1 = 32'd393
; 
32'd12655: dataIn1 = 32'd422
; 
32'd12656: dataIn1 = 32'd467
; 
32'd12657: dataIn1 = 32'd531
; 
32'd12658: dataIn1 = 32'd535
; 
32'd12659: dataIn1 = 32'd543
; 
32'd12660: dataIn1 = 32'd554
; 
32'd12661: dataIn1 = 32'd560
; 
32'd12662: dataIn1 = 32'd592
; 
32'd12663: dataIn1 = 32'd376
; 
32'd12664: dataIn1 = 32'd378
; 
32'd12665: dataIn1 = 32'd447
; 
32'd12666: dataIn1 = 32'd468
; 
32'd12667: dataIn1 = 32'd495
; 
32'd12668: dataIn1 = 32'd499
; 
32'd12669: dataIn1 = 32'd513
; 
32'd12670: dataIn1 = 32'd529
; 
32'd12671: dataIn1 = 32'd551
; 
32'd12672: dataIn1 = 32'd384
; 
32'd12673: dataIn1 = 32'd386
; 
32'd12674: dataIn1 = 32'd400
; 
32'd12675: dataIn1 = 32'd469
; 
32'd12676: dataIn1 = 32'd478
; 
32'd12677: dataIn1 = 32'd488
; 
32'd12678: dataIn1 = 32'd555
; 
32'd12679: dataIn1 = 32'd389
; 
32'd12680: dataIn1 = 32'd403
; 
32'd12681: dataIn1 = 32'd422
; 
32'd12682: dataIn1 = 32'd470
; 
32'd12683: dataIn1 = 32'd503
; 
32'd12684: dataIn1 = 32'd539
; 
32'd12685: dataIn1 = 32'd569
; 
32'd12686: dataIn1 = 32'd390
; 
32'd12687: dataIn1 = 32'd392
; 
32'd12688: dataIn1 = 32'd426
; 
32'd12689: dataIn1 = 32'd471
; 
32'd12690: dataIn1 = 32'd494
; 
32'd12691: dataIn1 = 32'd377
; 
32'd12692: dataIn1 = 32'd394
; 
32'd12693: dataIn1 = 32'd437
; 
32'd12694: dataIn1 = 32'd472
; 
32'd12695: dataIn1 = 32'd554
; 
32'd12696: dataIn1 = 32'd556
; 
32'd12697: dataIn1 = 32'd583
; 
32'd12698: dataIn1 = 32'd403
; 
32'd12699: dataIn1 = 32'd431
; 
32'd12700: dataIn1 = 32'd448
; 
32'd12701: dataIn1 = 32'd473
; 
32'd12702: dataIn1 = 32'd511
; 
32'd12703: dataIn1 = 32'd523
; 
32'd12704: dataIn1 = 32'd524
; 
32'd12705: dataIn1 = 32'd547
; 
32'd12706: dataIn1 = 32'd404
; 
32'd12707: dataIn1 = 32'd408
; 
32'd12708: dataIn1 = 32'd415
; 
32'd12709: dataIn1 = 32'd474
; 
32'd12710: dataIn1 = 32'd506
; 
32'd12711: dataIn1 = 32'd528
; 
32'd12712: dataIn1 = 32'd557
; 
32'd12713: dataIn1 = 32'd603
; 
32'd12714: dataIn1 = 32'd367
; 
32'd12715: dataIn1 = 32'd405
; 
32'd12716: dataIn1 = 32'd461
; 
32'd12717: dataIn1 = 32'd475
; 
32'd12718: dataIn1 = 32'd497
; 
32'd12719: dataIn1 = 32'd498
; 
32'd12720: dataIn1 = 32'd545
; 
32'd12721: dataIn1 = 32'd408
; 
32'd12722: dataIn1 = 32'd413
; 
32'd12723: dataIn1 = 32'd459
; 
32'd12724: dataIn1 = 32'd476
; 
32'd12725: dataIn1 = 32'd517
; 
32'd12726: dataIn1 = 32'd527
; 
32'd12727: dataIn1 = 32'd557
; 
32'd12728: dataIn1 = 32'd558
; 
32'd12729: dataIn1 = 32'd593
; 
32'd12730: dataIn1 = 32'd618
; 
32'd12731: dataIn1 = 32'd416
; 
32'd12732: dataIn1 = 32'd445
; 
32'd12733: dataIn1 = 32'd446
; 
32'd12734: dataIn1 = 32'd477
; 
32'd12735: dataIn1 = 32'd489
; 
32'd12736: dataIn1 = 32'd496
; 
32'd12737: dataIn1 = 32'd559
; 
32'd12738: dataIn1 = 32'd419
; 
32'd12739: dataIn1 = 32'd464
; 
32'd12740: dataIn1 = 32'd469
; 
32'd12741: dataIn1 = 32'd478
; 
32'd12742: dataIn1 = 32'd500
; 
32'd12743: dataIn1 = 32'd534
; 
32'd12744: dataIn1 = 32'd554
; 
32'd12745: dataIn1 = 32'd560
; 
32'd12746: dataIn1 = 32'd358
; 
32'd12747: dataIn1 = 32'd422
; 
32'd12748: dataIn1 = 32'd457
; 
32'd12749: dataIn1 = 32'd479
; 
32'd12750: dataIn1 = 32'd492
; 
32'd12751: dataIn1 = 32'd528
; 
32'd12752: dataIn1 = 32'd561
; 
32'd12753: dataIn1 = 32'd410
; 
32'd12754: dataIn1 = 32'd427
; 
32'd12755: dataIn1 = 32'd448
; 
32'd12756: dataIn1 = 32'd480
; 
32'd12757: dataIn1 = 32'd522
; 
32'd12758: dataIn1 = 32'd428
; 
32'd12759: dataIn1 = 32'd432
; 
32'd12760: dataIn1 = 32'd436
; 
32'd12761: dataIn1 = 32'd481
; 
32'd12762: dataIn1 = 32'd502
; 
32'd12763: dataIn1 = 32'd508
; 
32'd12764: dataIn1 = 32'd395
; 
32'd12765: dataIn1 = 32'd445
; 
32'd12766: dataIn1 = 32'd452
; 
32'd12767: dataIn1 = 32'd482
; 
32'd12768: dataIn1 = 32'd516
; 
32'd12769: dataIn1 = 32'd538
; 
32'd12770: dataIn1 = 32'd549
; 
32'd12771: dataIn1 = 32'd562
; 
32'd12772: dataIn1 = 32'd397
; 
32'd12773: dataIn1 = 32'd430
; 
32'd12774: dataIn1 = 32'd440
; 
32'd12775: dataIn1 = 32'd483
; 
32'd12776: dataIn1 = 32'd548
; 
32'd12777: dataIn1 = 32'd550
; 
32'd12778: dataIn1 = 32'd553
; 
32'd12779: dataIn1 = 32'd563
; 
32'd12780: dataIn1 = 32'd420
; 
32'd12781: dataIn1 = 32'd421
; 
32'd12782: dataIn1 = 32'd425
; 
32'd12783: dataIn1 = 32'd484
; 
32'd12784: dataIn1 = 32'd531
; 
32'd12785: dataIn1 = 32'd532
; 
32'd12786: dataIn1 = 32'd567
; 
32'd12787: dataIn1 = 32'd594
; 
32'd12788: dataIn1 = 32'd596
; 
32'd12789: dataIn1 = 32'd605
; 
32'd12790: dataIn1 = 32'd394
; 
32'd12791: dataIn1 = 32'd434
; 
32'd12792: dataIn1 = 32'd438
; 
32'd12793: dataIn1 = 32'd485
; 
32'd12794: dataIn1 = 32'd487
; 
32'd12795: dataIn1 = 32'd533
; 
32'd12796: dataIn1 = 32'd584
; 
32'd12797: dataIn1 = 32'd379
; 
32'd12798: dataIn1 = 32'd431
; 
32'd12799: dataIn1 = 32'd450
; 
32'd12800: dataIn1 = 32'd486
; 
32'd12801: dataIn1 = 32'd516
; 
32'd12802: dataIn1 = 32'd564
; 
32'd12803: dataIn1 = 32'd394
; 
32'd12804: dataIn1 = 32'd438
; 
32'd12805: dataIn1 = 32'd485
; 
32'd12806: dataIn1 = 32'd487
; 
32'd12807: dataIn1 = 32'd555
; 
32'd12808: dataIn1 = 32'd556
; 
32'd12809: dataIn1 = 32'd595
; 
32'd12810: dataIn1 = 32'd617
; 
32'd12811: dataIn1 = 32'd376
; 
32'd12812: dataIn1 = 32'd386
; 
32'd12813: dataIn1 = 32'd469
; 
32'd12814: dataIn1 = 32'd488
; 
32'd12815: dataIn1 = 32'd499
; 
32'd12816: dataIn1 = 32'd500
; 
32'd12817: dataIn1 = 32'd541
; 
32'd12818: dataIn1 = 32'd375
; 
32'd12819: dataIn1 = 32'd406
; 
32'd12820: dataIn1 = 32'd477
; 
32'd12821: dataIn1 = 32'd489
; 
32'd12822: dataIn1 = 32'd491
; 
32'd12823: dataIn1 = 32'd496
; 
32'd12824: dataIn1 = 32'd537
; 
32'd12825: dataIn1 = 32'd559
; 
32'd12826: dataIn1 = 32'd397
; 
32'd12827: dataIn1 = 32'd462
; 
32'd12828: dataIn1 = 32'd463
; 
32'd12829: dataIn1 = 32'd490
; 
32'd12830: dataIn1 = 32'd498
; 
32'd12831: dataIn1 = 32'd585
; 
32'd12832: dataIn1 = 32'd587
; 
32'd12833: dataIn1 = 32'd432
; 
32'd12834: dataIn1 = 32'd436
; 
32'd12835: dataIn1 = 32'd489
; 
32'd12836: dataIn1 = 32'd491
; 
32'd12837: dataIn1 = 32'd540
; 
32'd12838: dataIn1 = 32'd570
; 
32'd12839: dataIn1 = 32'd412
; 
32'd12840: dataIn1 = 32'd464
; 
32'd12841: dataIn1 = 32'd479
; 
32'd12842: dataIn1 = 32'd492
; 
32'd12843: dataIn1 = 32'd519
; 
32'd12844: dataIn1 = 32'd561
; 
32'd12845: dataIn1 = 32'd403
; 
32'd12846: dataIn1 = 32'd420
; 
32'd12847: dataIn1 = 32'd425
; 
32'd12848: dataIn1 = 32'd493
; 
32'd12849: dataIn1 = 32'd547
; 
32'd12850: dataIn1 = 32'd569
; 
32'd12851: dataIn1 = 32'd596
; 
32'd12852: dataIn1 = 32'd401
; 
32'd12853: dataIn1 = 32'd434
; 
32'd12854: dataIn1 = 32'd471
; 
32'd12855: dataIn1 = 32'd494
; 
32'd12856: dataIn1 = 32'd533
; 
32'd12857: dataIn1 = 32'd576
; 
32'd12858: dataIn1 = 32'd585
; 
32'd12859: dataIn1 = 32'd606
; 
32'd12860: dataIn1 = 32'd399
; 
32'd12861: dataIn1 = 32'd447
; 
32'd12862: dataIn1 = 32'd468
; 
32'd12863: dataIn1 = 32'd495
; 
32'd12864: dataIn1 = 32'd521
; 
32'd12865: dataIn1 = 32'd536
; 
32'd12866: dataIn1 = 32'd551
; 
32'd12867: dataIn1 = 32'd446
; 
32'd12868: dataIn1 = 32'd477
; 
32'd12869: dataIn1 = 32'd489
; 
32'd12870: dataIn1 = 32'd496
; 
32'd12871: dataIn1 = 32'd525
; 
32'd12872: dataIn1 = 32'd575
; 
32'd12873: dataIn1 = 32'd392
; 
32'd12874: dataIn1 = 32'd444
; 
32'd12875: dataIn1 = 32'd475
; 
32'd12876: dataIn1 = 32'd497
; 
32'd12877: dataIn1 = 32'd527
; 
32'd12878: dataIn1 = 32'd545
; 
32'd12879: dataIn1 = 32'd392
; 
32'd12880: dataIn1 = 32'd475
; 
32'd12881: dataIn1 = 32'd490
; 
32'd12882: dataIn1 = 32'd498
; 
32'd12883: dataIn1 = 32'd386
; 
32'd12884: dataIn1 = 32'd468
; 
32'd12885: dataIn1 = 32'd488
; 
32'd12886: dataIn1 = 32'd499
; 
32'd12887: dataIn1 = 32'd529
; 
32'd12888: dataIn1 = 32'd577
; 
32'd12889: dataIn1 = 32'd621
; 
32'd12890: dataIn1 = 32'd419
; 
32'd12891: dataIn1 = 32'd478
; 
32'd12892: dataIn1 = 32'd488
; 
32'd12893: dataIn1 = 32'd500
; 
32'd12894: dataIn1 = 32'd541
; 
32'd12895: dataIn1 = 32'd590
; 
32'd12896: dataIn1 = 32'd411
; 
32'd12897: dataIn1 = 32'd448
; 
32'd12898: dataIn1 = 32'd449
; 
32'd12899: dataIn1 = 32'd501
; 
32'd12900: dataIn1 = 32'd513
; 
32'd12901: dataIn1 = 32'd432
; 
32'd12902: dataIn1 = 32'd451
; 
32'd12903: dataIn1 = 32'd481
; 
32'd12904: dataIn1 = 32'd502
; 
32'd12905: dataIn1 = 32'd548
; 
32'd12906: dataIn1 = 32'd565
; 
32'd12907: dataIn1 = 32'd570
; 
32'd12908: dataIn1 = 32'd573
; 
32'd12909: dataIn1 = 32'd443
; 
32'd12910: dataIn1 = 32'd457
; 
32'd12911: dataIn1 = 32'd470
; 
32'd12912: dataIn1 = 32'd503
; 
32'd12913: dataIn1 = 32'd505
; 
32'd12914: dataIn1 = 32'd528
; 
32'd12915: dataIn1 = 32'd539
; 
32'd12916: dataIn1 = 32'd566
; 
32'd12917: dataIn1 = 32'd383
; 
32'd12918: dataIn1 = 32'd435
; 
32'd12919: dataIn1 = 32'd465
; 
32'd12920: dataIn1 = 32'd504
; 
32'd12921: dataIn1 = 32'd520
; 
32'd12922: dataIn1 = 32'd542
; 
32'd12923: dataIn1 = 32'd567
; 
32'd12924: dataIn1 = 32'd572
; 
32'd12925: dataIn1 = 32'd403
; 
32'd12926: dataIn1 = 32'd443
; 
32'd12927: dataIn1 = 32'd503
; 
32'd12928: dataIn1 = 32'd505
; 
32'd12929: dataIn1 = 32'd597
; 
32'd12930: dataIn1 = 32'd607
; 
32'd12931: dataIn1 = 32'd619
; 
32'd12932: dataIn1 = 32'd644
; 
32'd12933: dataIn1 = 32'd404
; 
32'd12934: dataIn1 = 32'd459
; 
32'd12935: dataIn1 = 32'd474
; 
32'd12936: dataIn1 = 32'd506
; 
32'd12937: dataIn1 = 32'd598
; 
32'd12938: dataIn1 = 32'd406
; 
32'd12939: dataIn1 = 32'd459
; 
32'd12940: dataIn1 = 32'd460
; 
32'd12941: dataIn1 = 32'd507
; 
32'd12942: dataIn1 = 32'd537
; 
32'd12943: dataIn1 = 32'd552
; 
32'd12944: dataIn1 = 32'd582
; 
32'd12945: dataIn1 = 32'd599
; 
32'd12946: dataIn1 = 32'd407
; 
32'd12947: dataIn1 = 32'd454
; 
32'd12948: dataIn1 = 32'd481
; 
32'd12949: dataIn1 = 32'd508
; 
32'd12950: dataIn1 = 32'd515
; 
32'd12951: dataIn1 = 32'd410
; 
32'd12952: dataIn1 = 32'd438
; 
32'd12953: dataIn1 = 32'd450
; 
32'd12954: dataIn1 = 32'd509
; 
32'd12955: dataIn1 = 32'd522
; 
32'd12956: dataIn1 = 32'd564
; 
32'd12957: dataIn1 = 32'd595
; 
32'd12958: dataIn1 = 32'd414
; 
32'd12959: dataIn1 = 32'd458
; 
32'd12960: dataIn1 = 32'd460
; 
32'd12961: dataIn1 = 32'd510
; 
32'd12962: dataIn1 = 32'd526
; 
32'd12963: dataIn1 = 32'd420
; 
32'd12964: dataIn1 = 32'd439
; 
32'd12965: dataIn1 = 32'd473
; 
32'd12966: dataIn1 = 32'd511
; 
32'd12967: dataIn1 = 32'd530
; 
32'd12968: dataIn1 = 32'd532
; 
32'd12969: dataIn1 = 32'd594
; 
32'd12970: dataIn1 = 32'd421
; 
32'd12971: dataIn1 = 32'd439
; 
32'd12972: dataIn1 = 32'd460
; 
32'd12973: dataIn1 = 32'd512
; 
32'd12974: dataIn1 = 32'd525
; 
32'd12975: dataIn1 = 32'd594
; 
32'd12976: dataIn1 = 32'd441
; 
32'd12977: dataIn1 = 32'd468
; 
32'd12978: dataIn1 = 32'd501
; 
32'd12979: dataIn1 = 32'd513
; 
32'd12980: dataIn1 = 32'd522
; 
32'd12981: dataIn1 = 32'd523
; 
32'd12982: dataIn1 = 32'd529
; 
32'd12983: dataIn1 = 32'd597
; 
32'd12984: dataIn1 = 32'd604
; 
32'd12985: dataIn1 = 32'd442
; 
32'd12986: dataIn1 = 32'd453
; 
32'd12987: dataIn1 = 32'd463
; 
32'd12988: dataIn1 = 32'd514
; 
32'd12989: dataIn1 = 32'd584
; 
32'd12990: dataIn1 = 32'd585
; 
32'd12991: dataIn1 = 32'd600
; 
32'd12992: dataIn1 = 32'd620
; 
32'd12993: dataIn1 = 32'd634
; 
32'd12994: dataIn1 = 32'd449
; 
32'd12995: dataIn1 = 32'd451
; 
32'd12996: dataIn1 = 32'd508
; 
32'd12997: dataIn1 = 32'd515
; 
32'd12998: dataIn1 = 32'd536
; 
32'd12999: dataIn1 = 32'd565
; 
32'd13000: dataIn1 = 32'd597
; 
32'd13001: dataIn1 = 32'd456
; 
32'd13002: dataIn1 = 32'd482
; 
32'd13003: dataIn1 = 32'd486
; 
32'd13004: dataIn1 = 32'd516
; 
32'd13005: dataIn1 = 32'd538
; 
32'd13006: dataIn1 = 32'd562
; 
32'd13007: dataIn1 = 32'd564
; 
32'd13008: dataIn1 = 32'd591
; 
32'd13009: dataIn1 = 32'd601
; 
32'd13010: dataIn1 = 32'd414
; 
32'd13011: dataIn1 = 32'd458
; 
32'd13012: dataIn1 = 32'd476
; 
32'd13013: dataIn1 = 32'd517
; 
32'd13014: dataIn1 = 32'd558
; 
32'd13015: dataIn1 = 32'd582
; 
32'd13016: dataIn1 = 32'd588
; 
32'd13017: dataIn1 = 32'd383
; 
32'd13018: dataIn1 = 32'd421
; 
32'd13019: dataIn1 = 32'd460
; 
32'd13020: dataIn1 = 32'd518
; 
32'd13021: dataIn1 = 32'd526
; 
32'd13022: dataIn1 = 32'd552
; 
32'd13023: dataIn1 = 32'd444
; 
32'd13024: dataIn1 = 32'd461
; 
32'd13025: dataIn1 = 32'd492
; 
32'd13026: dataIn1 = 32'd519
; 
32'd13027: dataIn1 = 32'd545
; 
32'd13028: dataIn1 = 32'd557
; 
32'd13029: dataIn1 = 32'd589
; 
32'd13030: dataIn1 = 32'd437
; 
32'd13031: dataIn1 = 32'd465
; 
32'd13032: dataIn1 = 32'd504
; 
32'd13033: dataIn1 = 32'd520
; 
32'd13034: dataIn1 = 32'd581
; 
32'd13035: dataIn1 = 32'd417
; 
32'd13036: dataIn1 = 32'd466
; 
32'd13037: dataIn1 = 32'd495
; 
32'd13038: dataIn1 = 32'd521
; 
32'd13039: dataIn1 = 32'd568
; 
32'd13040: dataIn1 = 32'd579
; 
32'd13041: dataIn1 = 32'd480
; 
32'd13042: dataIn1 = 32'd509
; 
32'd13043: dataIn1 = 32'd513
; 
32'd13044: dataIn1 = 32'd522
; 
32'd13045: dataIn1 = 32'd523
; 
32'd13046: dataIn1 = 32'd524
; 
32'd13047: dataIn1 = 32'd604
; 
32'd13048: dataIn1 = 32'd621
; 
32'd13049: dataIn1 = 32'd628
; 
32'd13050: dataIn1 = 32'd645
; 
32'd13051: dataIn1 = 32'd652
; 
32'd13052: dataIn1 = 32'd473
; 
32'd13053: dataIn1 = 32'd513
; 
32'd13054: dataIn1 = 32'd522
; 
32'd13055: dataIn1 = 32'd523
; 
32'd13056: dataIn1 = 32'd524
; 
32'd13057: dataIn1 = 32'd571
; 
32'd13058: dataIn1 = 32'd578
; 
32'd13059: dataIn1 = 32'd473
; 
32'd13060: dataIn1 = 32'd522
; 
32'd13061: dataIn1 = 32'd523
; 
32'd13062: dataIn1 = 32'd524
; 
32'd13063: dataIn1 = 32'd578
; 
32'd13064: dataIn1 = 32'd628
; 
32'd13065: dataIn1 = 32'd629
; 
32'd13066: dataIn1 = 32'd645
; 
32'd13067: dataIn1 = 32'd456
; 
32'd13068: dataIn1 = 32'd496
; 
32'd13069: dataIn1 = 32'd512
; 
32'd13070: dataIn1 = 32'd525
; 
32'd13071: dataIn1 = 32'd530
; 
32'd13072: dataIn1 = 32'd591
; 
32'd13073: dataIn1 = 32'd625
; 
32'd13074: dataIn1 = 32'd646
; 
32'd13075: dataIn1 = 32'd458
; 
32'd13076: dataIn1 = 32'd510
; 
32'd13077: dataIn1 = 32'd518
; 
32'd13078: dataIn1 = 32'd526
; 
32'd13079: dataIn1 = 32'd580
; 
32'd13080: dataIn1 = 32'd392
; 
32'd13081: dataIn1 = 32'd476
; 
32'd13082: dataIn1 = 32'd497
; 
32'd13083: dataIn1 = 32'd527
; 
32'd13084: dataIn1 = 32'd588
; 
32'd13085: dataIn1 = 32'd602
; 
32'd13086: dataIn1 = 32'd474
; 
32'd13087: dataIn1 = 32'd479
; 
32'd13088: dataIn1 = 32'd503
; 
32'd13089: dataIn1 = 32'd528
; 
32'd13090: dataIn1 = 32'd539
; 
32'd13091: dataIn1 = 32'd566
; 
32'd13092: dataIn1 = 32'd574
; 
32'd13093: dataIn1 = 32'd603
; 
32'd13094: dataIn1 = 32'd468
; 
32'd13095: dataIn1 = 32'd499
; 
32'd13096: dataIn1 = 32'd513
; 
32'd13097: dataIn1 = 32'd529
; 
32'd13098: dataIn1 = 32'd586
; 
32'd13099: dataIn1 = 32'd604
; 
32'd13100: dataIn1 = 32'd621
; 
32'd13101: dataIn1 = 32'd640
; 
32'd13102: dataIn1 = 32'd456
; 
32'd13103: dataIn1 = 32'd511
; 
32'd13104: dataIn1 = 32'd525
; 
32'd13105: dataIn1 = 32'd530
; 
32'd13106: dataIn1 = 32'd591
; 
32'd13107: dataIn1 = 32'd625
; 
32'd13108: dataIn1 = 32'd629
; 
32'd13109: dataIn1 = 32'd437
; 
32'd13110: dataIn1 = 32'd467
; 
32'd13111: dataIn1 = 32'd484
; 
32'd13112: dataIn1 = 32'd531
; 
32'd13113: dataIn1 = 32'd535
; 
32'd13114: dataIn1 = 32'd583
; 
32'd13115: dataIn1 = 32'd605
; 
32'd13116: dataIn1 = 32'd420
; 
32'd13117: dataIn1 = 32'd484
; 
32'd13118: dataIn1 = 32'd511
; 
32'd13119: dataIn1 = 32'd532
; 
32'd13120: dataIn1 = 32'd596
; 
32'd13121: dataIn1 = 32'd465
; 
32'd13122: dataIn1 = 32'd485
; 
32'd13123: dataIn1 = 32'd494
; 
32'd13124: dataIn1 = 32'd533
; 
32'd13125: dataIn1 = 32'd542
; 
32'd13126: dataIn1 = 32'd572
; 
32'd13127: dataIn1 = 32'd584
; 
32'd13128: dataIn1 = 32'd606
; 
32'd13129: dataIn1 = 32'd631
; 
32'd13130: dataIn1 = 32'd633
; 
32'd13131: dataIn1 = 32'd461
; 
32'd13132: dataIn1 = 32'd464
; 
32'd13133: dataIn1 = 32'd478
; 
32'd13134: dataIn1 = 32'd534
; 
32'd13135: dataIn1 = 32'd560
; 
32'd13136: dataIn1 = 32'd589
; 
32'd13137: dataIn1 = 32'd590
; 
32'd13138: dataIn1 = 32'd630
; 
32'd13139: dataIn1 = 32'd425
; 
32'd13140: dataIn1 = 32'd467
; 
32'd13141: dataIn1 = 32'd531
; 
32'd13142: dataIn1 = 32'd535
; 
32'd13143: dataIn1 = 32'd543
; 
32'd13144: dataIn1 = 32'd441
; 
32'd13145: dataIn1 = 32'd495
; 
32'd13146: dataIn1 = 32'd515
; 
32'd13147: dataIn1 = 32'd536
; 
32'd13148: dataIn1 = 32'd568
; 
32'd13149: dataIn1 = 32'd459
; 
32'd13150: dataIn1 = 32'd489
; 
32'd13151: dataIn1 = 32'd507
; 
32'd13152: dataIn1 = 32'd537
; 
32'd13153: dataIn1 = 32'd540
; 
32'd13154: dataIn1 = 32'd575
; 
32'd13155: dataIn1 = 32'd599
; 
32'd13156: dataIn1 = 32'd623
; 
32'd13157: dataIn1 = 32'd660
; 
32'd13158: dataIn1 = 32'd450
; 
32'd13159: dataIn1 = 32'd482
; 
32'd13160: dataIn1 = 32'd516
; 
32'd13161: dataIn1 = 32'd538
; 
32'd13162: dataIn1 = 32'd470
; 
32'd13163: dataIn1 = 32'd503
; 
32'd13164: dataIn1 = 32'd528
; 
32'd13165: dataIn1 = 32'd539
; 
32'd13166: dataIn1 = 32'd543
; 
32'd13167: dataIn1 = 32'd607
; 
32'd13168: dataIn1 = 32'd454
; 
32'd13169: dataIn1 = 32'd491
; 
32'd13170: dataIn1 = 32'd537
; 
32'd13171: dataIn1 = 32'd540
; 
32'd13172: dataIn1 = 32'd565
; 
32'd13173: dataIn1 = 32'd608
; 
32'd13174: dataIn1 = 32'd660
; 
32'd13175: dataIn1 = 32'd447
; 
32'd13176: dataIn1 = 32'd488
; 
32'd13177: dataIn1 = 32'd500
; 
32'd13178: dataIn1 = 32'd541
; 
32'd13179: dataIn1 = 32'd577
; 
32'd13180: dataIn1 = 32'd586
; 
32'd13181: dataIn1 = 32'd609
; 
32'd13182: dataIn1 = 32'd458
; 
32'd13183: dataIn1 = 32'd504
; 
32'd13184: dataIn1 = 32'd533
; 
32'd13185: dataIn1 = 32'd542
; 
32'd13186: dataIn1 = 32'd576
; 
32'd13187: dataIn1 = 32'd610
; 
32'd13188: dataIn1 = 32'd467
; 
32'd13189: dataIn1 = 32'd535
; 
32'd13190: dataIn1 = 32'd539
; 
32'd13191: dataIn1 = 32'd543
; 
32'd13192: dataIn1 = 32'd592
; 
32'd13193: dataIn1 = 32'd622
; 
32'd13194: dataIn1 = 32'd627
; 
32'd13195: dataIn1 = 32'd447
; 
32'd13196: dataIn1 = 32'd461
; 
32'd13197: dataIn1 = 32'd466
; 
32'd13198: dataIn1 = 32'd544
; 
32'd13199: dataIn1 = 32'd590
; 
32'd13200: dataIn1 = 32'd611
; 
32'd13201: dataIn1 = 32'd614
; 
32'd13202: dataIn1 = 32'd666
; 
32'd13203: dataIn1 = 32'd475
; 
32'd13204: dataIn1 = 32'd497
; 
32'd13205: dataIn1 = 32'd519
; 
32'd13206: dataIn1 = 32'd545
; 
32'd13207: dataIn1 = 32'd546
; 
32'd13208: dataIn1 = 32'd589
; 
32'd13209: dataIn1 = 32'd593
; 
32'd13210: dataIn1 = 32'd611
; 
32'd13211: dataIn1 = 32'd636
; 
32'd13212: dataIn1 = 32'd638
; 
32'd13213: dataIn1 = 32'd397
; 
32'd13214: dataIn1 = 32'd461
; 
32'd13215: dataIn1 = 32'd545
; 
32'd13216: dataIn1 = 32'd546
; 
32'd13217: dataIn1 = 32'd587
; 
32'd13218: dataIn1 = 32'd611
; 
32'd13219: dataIn1 = 32'd403
; 
32'd13220: dataIn1 = 32'd473
; 
32'd13221: dataIn1 = 32'd493
; 
32'd13222: dataIn1 = 32'd547
; 
32'd13223: dataIn1 = 32'd571
; 
32'd13224: dataIn1 = 32'd578
; 
32'd13225: dataIn1 = 32'd619
; 
32'd13226: dataIn1 = 32'd417
; 
32'd13227: dataIn1 = 32'd483
; 
32'd13228: dataIn1 = 32'd502
; 
32'd13229: dataIn1 = 32'd548
; 
32'd13230: dataIn1 = 32'd550
; 
32'd13231: dataIn1 = 32'd553
; 
32'd13232: dataIn1 = 32'd612
; 
32'd13233: dataIn1 = 32'd430
; 
32'd13234: dataIn1 = 32'd453
; 
32'd13235: dataIn1 = 32'd482
; 
32'd13236: dataIn1 = 32'd549
; 
32'd13237: dataIn1 = 32'd563
; 
32'd13238: dataIn1 = 32'd600
; 
32'd13239: dataIn1 = 32'd613
; 
32'd13240: dataIn1 = 32'd445
; 
32'd13241: dataIn1 = 32'd483
; 
32'd13242: dataIn1 = 32'd548
; 
32'd13243: dataIn1 = 32'd550
; 
32'd13244: dataIn1 = 32'd573
; 
32'd13245: dataIn1 = 32'd612
; 
32'd13246: dataIn1 = 32'd447
; 
32'd13247: dataIn1 = 32'd468
; 
32'd13248: dataIn1 = 32'd495
; 
32'd13249: dataIn1 = 32'd551
; 
32'd13250: dataIn1 = 32'd579
; 
32'd13251: dataIn1 = 32'd586
; 
32'd13252: dataIn1 = 32'd460
; 
32'd13253: dataIn1 = 32'd507
; 
32'd13254: dataIn1 = 32'd518
; 
32'd13255: dataIn1 = 32'd552
; 
32'd13256: dataIn1 = 32'd567
; 
32'd13257: dataIn1 = 32'd580
; 
32'd13258: dataIn1 = 32'd582
; 
32'd13259: dataIn1 = 32'd632
; 
32'd13260: dataIn1 = 32'd646
; 
32'd13261: dataIn1 = 32'd647
; 
32'd13262: dataIn1 = 32'd692
; 
32'd13263: dataIn1 = 32'd717
; 
32'd13264: dataIn1 = 32'd466
; 
32'd13265: dataIn1 = 32'd483
; 
32'd13266: dataIn1 = 32'd548
; 
32'd13267: dataIn1 = 32'd553
; 
32'd13268: dataIn1 = 32'd612
; 
32'd13269: dataIn1 = 32'd614
; 
32'd13270: dataIn1 = 32'd639
; 
32'd13271: dataIn1 = 32'd648
; 
32'd13272: dataIn1 = 32'd467
; 
32'd13273: dataIn1 = 32'd472
; 
32'd13274: dataIn1 = 32'd478
; 
32'd13275: dataIn1 = 32'd554
; 
32'd13276: dataIn1 = 32'd555
; 
32'd13277: dataIn1 = 32'd583
; 
32'd13278: dataIn1 = 32'd615
; 
32'd13279: dataIn1 = 32'd469
; 
32'd13280: dataIn1 = 32'd487
; 
32'd13281: dataIn1 = 32'd554
; 
32'd13282: dataIn1 = 32'd555
; 
32'd13283: dataIn1 = 32'd556
; 
32'd13284: dataIn1 = 32'd577
; 
32'd13285: dataIn1 = 32'd616
; 
32'd13286: dataIn1 = 32'd617
; 
32'd13287: dataIn1 = 32'd472
; 
32'd13288: dataIn1 = 32'd487
; 
32'd13289: dataIn1 = 32'd555
; 
32'd13290: dataIn1 = 32'd556
; 
32'd13291: dataIn1 = 32'd581
; 
32'd13292: dataIn1 = 32'd616
; 
32'd13293: dataIn1 = 32'd617
; 
32'd13294: dataIn1 = 32'd474
; 
32'd13295: dataIn1 = 32'd476
; 
32'd13296: dataIn1 = 32'd519
; 
32'd13297: dataIn1 = 32'd557
; 
32'd13298: dataIn1 = 32'd574
; 
32'd13299: dataIn1 = 32'd593
; 
32'd13300: dataIn1 = 32'd603
; 
32'd13301: dataIn1 = 32'd618
; 
32'd13302: dataIn1 = 32'd626
; 
32'd13303: dataIn1 = 32'd649
; 
32'd13304: dataIn1 = 32'd693
; 
32'd13305: dataIn1 = 32'd459
; 
32'd13306: dataIn1 = 32'd476
; 
32'd13307: dataIn1 = 32'd517
; 
32'd13308: dataIn1 = 32'd558
; 
32'd13309: dataIn1 = 32'd598
; 
32'd13310: dataIn1 = 32'd599
; 
32'd13311: dataIn1 = 32'd618
; 
32'd13312: dataIn1 = 32'd661
; 
32'd13313: dataIn1 = 32'd445
; 
32'd13314: dataIn1 = 32'd477
; 
32'd13315: dataIn1 = 32'd489
; 
32'd13316: dataIn1 = 32'd559
; 
32'd13317: dataIn1 = 32'd562
; 
32'd13318: dataIn1 = 32'd570
; 
32'd13319: dataIn1 = 32'd575
; 
32'd13320: dataIn1 = 32'd467
; 
32'd13321: dataIn1 = 32'd478
; 
32'd13322: dataIn1 = 32'd534
; 
32'd13323: dataIn1 = 32'd560
; 
32'd13324: dataIn1 = 32'd561
; 
32'd13325: dataIn1 = 32'd630
; 
32'd13326: dataIn1 = 32'd650
; 
32'd13327: dataIn1 = 32'd479
; 
32'd13328: dataIn1 = 32'd492
; 
32'd13329: dataIn1 = 32'd560
; 
32'd13330: dataIn1 = 32'd561
; 
32'd13331: dataIn1 = 32'd574
; 
32'd13332: dataIn1 = 32'd627
; 
32'd13333: dataIn1 = 32'd482
; 
32'd13334: dataIn1 = 32'd516
; 
32'd13335: dataIn1 = 32'd559
; 
32'd13336: dataIn1 = 32'd562
; 
32'd13337: dataIn1 = 32'd613
; 
32'd13338: dataIn1 = 32'd624
; 
32'd13339: dataIn1 = 32'd651
; 
32'd13340: dataIn1 = 32'd430
; 
32'd13341: dataIn1 = 32'd483
; 
32'd13342: dataIn1 = 32'd549
; 
32'd13343: dataIn1 = 32'd563
; 
32'd13344: dataIn1 = 32'd641
; 
32'd13345: dataIn1 = 32'd486
; 
32'd13346: dataIn1 = 32'd509
; 
32'd13347: dataIn1 = 32'd516
; 
32'd13348: dataIn1 = 32'd564
; 
32'd13349: dataIn1 = 32'd601
; 
32'd13350: dataIn1 = 32'd620
; 
32'd13351: dataIn1 = 32'd652
; 
32'd13352: dataIn1 = 32'd502
; 
32'd13353: dataIn1 = 32'd515
; 
32'd13354: dataIn1 = 32'd540
; 
32'd13355: dataIn1 = 32'd565
; 
32'd13356: dataIn1 = 32'd568
; 
32'd13357: dataIn1 = 32'd608
; 
32'd13358: dataIn1 = 32'd653
; 
32'd13359: dataIn1 = 32'd654
; 
32'd13360: dataIn1 = 32'd659
; 
32'd13361: dataIn1 = 32'd665
; 
32'd13362: dataIn1 = 32'd687
; 
32'd13363: dataIn1 = 32'd694
; 
32'd13364: dataIn1 = 32'd454
; 
32'd13365: dataIn1 = 32'd503
; 
32'd13366: dataIn1 = 32'd528
; 
32'd13367: dataIn1 = 32'd566
; 
32'd13368: dataIn1 = 32'd607
; 
32'd13369: dataIn1 = 32'd608
; 
32'd13370: dataIn1 = 32'd626
; 
32'd13371: dataIn1 = 32'd484
; 
32'd13372: dataIn1 = 32'd504
; 
32'd13373: dataIn1 = 32'd552
; 
32'd13374: dataIn1 = 32'd567
; 
32'd13375: dataIn1 = 32'd572
; 
32'd13376: dataIn1 = 32'd610
; 
32'd13377: dataIn1 = 32'd643
; 
32'd13378: dataIn1 = 32'd521
; 
32'd13379: dataIn1 = 32'd536
; 
32'd13380: dataIn1 = 32'd565
; 
32'd13381: dataIn1 = 32'd568
; 
32'd13382: dataIn1 = 32'd579
; 
32'd13383: dataIn1 = 32'd642
; 
32'd13384: dataIn1 = 32'd653
; 
32'd13385: dataIn1 = 32'd654
; 
32'd13386: dataIn1 = 32'd687
; 
32'd13387: dataIn1 = 32'd691
; 
32'd13388: dataIn1 = 32'd695
; 
32'd13389: dataIn1 = 32'd403
; 
32'd13390: dataIn1 = 32'd470
; 
32'd13391: dataIn1 = 32'd493
; 
32'd13392: dataIn1 = 32'd569
; 
32'd13393: dataIn1 = 32'd619
; 
32'd13394: dataIn1 = 32'd491
; 
32'd13395: dataIn1 = 32'd502
; 
32'd13396: dataIn1 = 32'd559
; 
32'd13397: dataIn1 = 32'd570
; 
32'd13398: dataIn1 = 32'd573
; 
32'd13399: dataIn1 = 32'd623
; 
32'd13400: dataIn1 = 32'd403
; 
32'd13401: dataIn1 = 32'd523
; 
32'd13402: dataIn1 = 32'd547
; 
32'd13403: dataIn1 = 32'd571
; 
32'd13404: dataIn1 = 32'd504
; 
32'd13405: dataIn1 = 32'd533
; 
32'd13406: dataIn1 = 32'd567
; 
32'd13407: dataIn1 = 32'd572
; 
32'd13408: dataIn1 = 32'd581
; 
32'd13409: dataIn1 = 32'd631
; 
32'd13410: dataIn1 = 32'd643
; 
32'd13411: dataIn1 = 32'd502
; 
32'd13412: dataIn1 = 32'd550
; 
32'd13413: dataIn1 = 32'd570
; 
32'd13414: dataIn1 = 32'd573
; 
32'd13415: dataIn1 = 32'd653
; 
32'd13416: dataIn1 = 32'd655
; 
32'd13417: dataIn1 = 32'd528
; 
32'd13418: dataIn1 = 32'd557
; 
32'd13419: dataIn1 = 32'd561
; 
32'd13420: dataIn1 = 32'd574
; 
32'd13421: dataIn1 = 32'd649
; 
32'd13422: dataIn1 = 32'd496
; 
32'd13423: dataIn1 = 32'd537
; 
32'd13424: dataIn1 = 32'd559
; 
32'd13425: dataIn1 = 32'd575
; 
32'd13426: dataIn1 = 32'd623
; 
32'd13427: dataIn1 = 32'd646
; 
32'd13428: dataIn1 = 32'd651
; 
32'd13429: dataIn1 = 32'd458
; 
32'd13430: dataIn1 = 32'd494
; 
32'd13431: dataIn1 = 32'd542
; 
32'd13432: dataIn1 = 32'd576
; 
32'd13433: dataIn1 = 32'd633
; 
32'd13434: dataIn1 = 32'd499
; 
32'd13435: dataIn1 = 32'd541
; 
32'd13436: dataIn1 = 32'd555
; 
32'd13437: dataIn1 = 32'd577
; 
32'd13438: dataIn1 = 32'd615
; 
32'd13439: dataIn1 = 32'd635
; 
32'd13440: dataIn1 = 32'd656
; 
32'd13441: dataIn1 = 32'd696
; 
32'd13442: dataIn1 = 32'd523
; 
32'd13443: dataIn1 = 32'd524
; 
32'd13444: dataIn1 = 32'd547
; 
32'd13445: dataIn1 = 32'd578
; 
32'd13446: dataIn1 = 32'd628
; 
32'd13447: dataIn1 = 32'd644
; 
32'd13448: dataIn1 = 32'd657
; 
32'd13449: dataIn1 = 32'd670
; 
32'd13450: dataIn1 = 32'd671
; 
32'd13451: dataIn1 = 32'd697
; 
32'd13452: dataIn1 = 32'd521
; 
32'd13453: dataIn1 = 32'd551
; 
32'd13454: dataIn1 = 32'd568
; 
32'd13455: dataIn1 = 32'd579
; 
32'd13456: dataIn1 = 32'd609
; 
32'd13457: dataIn1 = 32'd614
; 
32'd13458: dataIn1 = 32'd642
; 
32'd13459: dataIn1 = 32'd458
; 
32'd13460: dataIn1 = 32'd526
; 
32'd13461: dataIn1 = 32'd552
; 
32'd13462: dataIn1 = 32'd580
; 
32'd13463: dataIn1 = 32'd610
; 
32'd13464: dataIn1 = 32'd520
; 
32'd13465: dataIn1 = 32'd556
; 
32'd13466: dataIn1 = 32'd572
; 
32'd13467: dataIn1 = 32'd581
; 
32'd13468: dataIn1 = 32'd637
; 
32'd13469: dataIn1 = 32'd507
; 
32'd13470: dataIn1 = 32'd517
; 
32'd13471: dataIn1 = 32'd552
; 
32'd13472: dataIn1 = 32'd582
; 
32'd13473: dataIn1 = 32'd632
; 
32'd13474: dataIn1 = 32'd472
; 
32'd13475: dataIn1 = 32'd531
; 
32'd13476: dataIn1 = 32'd554
; 
32'd13477: dataIn1 = 32'd583
; 
32'd13478: dataIn1 = 32'd592
; 
32'd13479: dataIn1 = 32'd616
; 
32'd13480: dataIn1 = 32'd637
; 
32'd13481: dataIn1 = 32'd658
; 
32'd13482: dataIn1 = 32'd485
; 
32'd13483: dataIn1 = 32'd514
; 
32'd13484: dataIn1 = 32'd533
; 
32'd13485: dataIn1 = 32'd584
; 
32'd13486: dataIn1 = 32'd595
; 
32'd13487: dataIn1 = 32'd631
; 
32'd13488: dataIn1 = 32'd634
; 
32'd13489: dataIn1 = 32'd672
; 
32'd13490: dataIn1 = 32'd490
; 
32'd13491: dataIn1 = 32'd494
; 
32'd13492: dataIn1 = 32'd514
; 
32'd13493: dataIn1 = 32'd585
; 
32'd13494: dataIn1 = 32'd587
; 
32'd13495: dataIn1 = 32'd600
; 
32'd13496: dataIn1 = 32'd602
; 
32'd13497: dataIn1 = 32'd606
; 
32'd13498: dataIn1 = 32'd634
; 
32'd13499: dataIn1 = 32'd641
; 
32'd13500: dataIn1 = 32'd681
; 
32'd13501: dataIn1 = 32'd698
; 
32'd13502: dataIn1 = 32'd529
; 
32'd13503: dataIn1 = 32'd541
; 
32'd13504: dataIn1 = 32'd551
; 
32'd13505: dataIn1 = 32'd586
; 
32'd13506: dataIn1 = 32'd640
; 
32'd13507: dataIn1 = 32'd642
; 
32'd13508: dataIn1 = 32'd490
; 
32'd13509: dataIn1 = 32'd546
; 
32'd13510: dataIn1 = 32'd585
; 
32'd13511: dataIn1 = 32'd587
; 
32'd13512: dataIn1 = 32'd638
; 
32'd13513: dataIn1 = 32'd639
; 
32'd13514: dataIn1 = 32'd641
; 
32'd13515: dataIn1 = 32'd684
; 
32'd13516: dataIn1 = 32'd458
; 
32'd13517: dataIn1 = 32'd517
; 
32'd13518: dataIn1 = 32'd527
; 
32'd13519: dataIn1 = 32'd588
; 
32'd13520: dataIn1 = 32'd602
; 
32'd13521: dataIn1 = 32'd632
; 
32'd13522: dataIn1 = 32'd668
; 
32'd13523: dataIn1 = 32'd519
; 
32'd13524: dataIn1 = 32'd534
; 
32'd13525: dataIn1 = 32'd545
; 
32'd13526: dataIn1 = 32'd589
; 
32'd13527: dataIn1 = 32'd649
; 
32'd13528: dataIn1 = 32'd677
; 
32'd13529: dataIn1 = 32'd699
; 
32'd13530: dataIn1 = 32'd740
; 
32'd13531: dataIn1 = 32'd500
; 
32'd13532: dataIn1 = 32'd534
; 
32'd13533: dataIn1 = 32'd544
; 
32'd13534: dataIn1 = 32'd590
; 
32'd13535: dataIn1 = 32'd609
; 
32'd13536: dataIn1 = 32'd615
; 
32'd13537: dataIn1 = 32'd630
; 
32'd13538: dataIn1 = 32'd669
; 
32'd13539: dataIn1 = 32'd699
; 
32'd13540: dataIn1 = 32'd700
; 
32'd13541: dataIn1 = 32'd716
; 
32'd13542: dataIn1 = 32'd516
; 
32'd13543: dataIn1 = 32'd525
; 
32'd13544: dataIn1 = 32'd530
; 
32'd13545: dataIn1 = 32'd591
; 
32'd13546: dataIn1 = 32'd629
; 
32'd13547: dataIn1 = 32'd678
; 
32'd13548: dataIn1 = 32'd686
; 
32'd13549: dataIn1 = 32'd734
; 
32'd13550: dataIn1 = 32'd467
; 
32'd13551: dataIn1 = 32'd543
; 
32'd13552: dataIn1 = 32'd583
; 
32'd13553: dataIn1 = 32'd592
; 
32'd13554: dataIn1 = 32'd627
; 
32'd13555: dataIn1 = 32'd658
; 
32'd13556: dataIn1 = 32'd663
; 
32'd13557: dataIn1 = 32'd664
; 
32'd13558: dataIn1 = 32'd683
; 
32'd13559: dataIn1 = 32'd741
; 
32'd13560: dataIn1 = 32'd476
; 
32'd13561: dataIn1 = 32'd545
; 
32'd13562: dataIn1 = 32'd557
; 
32'd13563: dataIn1 = 32'd593
; 
32'd13564: dataIn1 = 32'd484
; 
32'd13565: dataIn1 = 32'd511
; 
32'd13566: dataIn1 = 32'd512
; 
32'd13567: dataIn1 = 32'd594
; 
32'd13568: dataIn1 = 32'd625
; 
32'd13569: dataIn1 = 32'd657
; 
32'd13570: dataIn1 = 32'd487
; 
32'd13571: dataIn1 = 32'd509
; 
32'd13572: dataIn1 = 32'd584
; 
32'd13573: dataIn1 = 32'd595
; 
32'd13574: dataIn1 = 32'd620
; 
32'd13575: dataIn1 = 32'd656
; 
32'd13576: dataIn1 = 32'd484
; 
32'd13577: dataIn1 = 32'd493
; 
32'd13578: dataIn1 = 32'd532
; 
32'd13579: dataIn1 = 32'd596
; 
32'd13580: dataIn1 = 32'd605
; 
32'd13581: dataIn1 = 32'd622
; 
32'd13582: dataIn1 = 32'd657
; 
32'd13583: dataIn1 = 32'd663
; 
32'd13584: dataIn1 = 32'd505
; 
32'd13585: dataIn1 = 32'd513
; 
32'd13586: dataIn1 = 32'd515
; 
32'd13587: dataIn1 = 32'd597
; 
32'd13588: dataIn1 = 32'd654
; 
32'd13589: dataIn1 = 32'd659
; 
32'd13590: dataIn1 = 32'd662
; 
32'd13591: dataIn1 = 32'd671
; 
32'd13592: dataIn1 = 32'd673
; 
32'd13593: dataIn1 = 32'd459
; 
32'd13594: dataIn1 = 32'd506
; 
32'd13595: dataIn1 = 32'd558
; 
32'd13596: dataIn1 = 32'd598
; 
32'd13597: dataIn1 = 32'd660
; 
32'd13598: dataIn1 = 32'd661
; 
32'd13599: dataIn1 = 32'd507
; 
32'd13600: dataIn1 = 32'd537
; 
32'd13601: dataIn1 = 32'd558
; 
32'd13602: dataIn1 = 32'd599
; 
32'd13603: dataIn1 = 32'd661
; 
32'd13604: dataIn1 = 32'd682
; 
32'd13605: dataIn1 = 32'd685
; 
32'd13606: dataIn1 = 32'd701
; 
32'd13607: dataIn1 = 32'd514
; 
32'd13608: dataIn1 = 32'd549
; 
32'd13609: dataIn1 = 32'd585
; 
32'd13610: dataIn1 = 32'd600
; 
32'd13611: dataIn1 = 32'd601
; 
32'd13612: dataIn1 = 32'd613
; 
32'd13613: dataIn1 = 32'd698
; 
32'd13614: dataIn1 = 32'd702
; 
32'd13615: dataIn1 = 32'd713
; 
32'd13616: dataIn1 = 32'd723
; 
32'd13617: dataIn1 = 32'd516
; 
32'd13618: dataIn1 = 32'd564
; 
32'd13619: dataIn1 = 32'd600
; 
32'd13620: dataIn1 = 32'd601
; 
32'd13621: dataIn1 = 32'd678
; 
32'd13622: dataIn1 = 32'd688
; 
32'd13623: dataIn1 = 32'd703
; 
32'd13624: dataIn1 = 32'd527
; 
32'd13625: dataIn1 = 32'd585
; 
32'd13626: dataIn1 = 32'd588
; 
32'd13627: dataIn1 = 32'd602
; 
32'd13628: dataIn1 = 32'd636
; 
32'd13629: dataIn1 = 32'd638
; 
32'd13630: dataIn1 = 32'd667
; 
32'd13631: dataIn1 = 32'd675
; 
32'd13632: dataIn1 = 32'd729
; 
32'd13633: dataIn1 = 32'd744
; 
32'd13634: dataIn1 = 32'd474
; 
32'd13635: dataIn1 = 32'd528
; 
32'd13636: dataIn1 = 32'd557
; 
32'd13637: dataIn1 = 32'd603
; 
32'd13638: dataIn1 = 32'd513
; 
32'd13639: dataIn1 = 32'd522
; 
32'd13640: dataIn1 = 32'd529
; 
32'd13641: dataIn1 = 32'd604
; 
32'd13642: dataIn1 = 32'd662
; 
32'd13643: dataIn1 = 32'd671
; 
32'd13644: dataIn1 = 32'd676
; 
32'd13645: dataIn1 = 32'd704
; 
32'd13646: dataIn1 = 32'd484
; 
32'd13647: dataIn1 = 32'd531
; 
32'd13648: dataIn1 = 32'd596
; 
32'd13649: dataIn1 = 32'd605
; 
32'd13650: dataIn1 = 32'd647
; 
32'd13651: dataIn1 = 32'd663
; 
32'd13652: dataIn1 = 32'd683
; 
32'd13653: dataIn1 = 32'd705
; 
32'd13654: dataIn1 = 32'd714
; 
32'd13655: dataIn1 = 32'd494
; 
32'd13656: dataIn1 = 32'd533
; 
32'd13657: dataIn1 = 32'd585
; 
32'd13658: dataIn1 = 32'd606
; 
32'd13659: dataIn1 = 32'd633
; 
32'd13660: dataIn1 = 32'd675
; 
32'd13661: dataIn1 = 32'd505
; 
32'd13662: dataIn1 = 32'd539
; 
32'd13663: dataIn1 = 32'd566
; 
32'd13664: dataIn1 = 32'd607
; 
32'd13665: dataIn1 = 32'd659
; 
32'd13666: dataIn1 = 32'd664
; 
32'd13667: dataIn1 = 32'd689
; 
32'd13668: dataIn1 = 32'd706
; 
32'd13669: dataIn1 = 32'd736
; 
32'd13670: dataIn1 = 32'd765
; 
32'd13671: dataIn1 = 32'd540
; 
32'd13672: dataIn1 = 32'd565
; 
32'd13673: dataIn1 = 32'd566
; 
32'd13674: dataIn1 = 32'd608
; 
32'd13675: dataIn1 = 32'd626
; 
32'd13676: dataIn1 = 32'd665
; 
32'd13677: dataIn1 = 32'd707
; 
32'd13678: dataIn1 = 32'd541
; 
32'd13679: dataIn1 = 32'd579
; 
32'd13680: dataIn1 = 32'd590
; 
32'd13681: dataIn1 = 32'd609
; 
32'd13682: dataIn1 = 32'd666
; 
32'd13683: dataIn1 = 32'd679
; 
32'd13684: dataIn1 = 32'd542
; 
32'd13685: dataIn1 = 32'd567
; 
32'd13686: dataIn1 = 32'd580
; 
32'd13687: dataIn1 = 32'd610
; 
32'd13688: dataIn1 = 32'd643
; 
32'd13689: dataIn1 = 32'd667
; 
32'd13690: dataIn1 = 32'd680
; 
32'd13691: dataIn1 = 32'd690
; 
32'd13692: dataIn1 = 32'd544
; 
32'd13693: dataIn1 = 32'd545
; 
32'd13694: dataIn1 = 32'd546
; 
32'd13695: dataIn1 = 32'd611
; 
32'd13696: dataIn1 = 32'd639
; 
32'd13697: dataIn1 = 32'd699
; 
32'd13698: dataIn1 = 32'd708
; 
32'd13699: dataIn1 = 32'd548
; 
32'd13700: dataIn1 = 32'd550
; 
32'd13701: dataIn1 = 32'd553
; 
32'd13702: dataIn1 = 32'd612
; 
32'd13703: dataIn1 = 32'd624
; 
32'd13704: dataIn1 = 32'd648
; 
32'd13705: dataIn1 = 32'd702
; 
32'd13706: dataIn1 = 32'd709
; 
32'd13707: dataIn1 = 32'd549
; 
32'd13708: dataIn1 = 32'd562
; 
32'd13709: dataIn1 = 32'd600
; 
32'd13710: dataIn1 = 32'd613
; 
32'd13711: dataIn1 = 32'd624
; 
32'd13712: dataIn1 = 32'd544
; 
32'd13713: dataIn1 = 32'd553
; 
32'd13714: dataIn1 = 32'd579
; 
32'd13715: dataIn1 = 32'd614
; 
32'd13716: dataIn1 = 32'd648
; 
32'd13717: dataIn1 = 32'd666
; 
32'd13718: dataIn1 = 32'd554
; 
32'd13719: dataIn1 = 32'd577
; 
32'd13720: dataIn1 = 32'd590
; 
32'd13721: dataIn1 = 32'd615
; 
32'd13722: dataIn1 = 32'd635
; 
32'd13723: dataIn1 = 32'd658
; 
32'd13724: dataIn1 = 32'd669
; 
32'd13725: dataIn1 = 32'd555
; 
32'd13726: dataIn1 = 32'd556
; 
32'd13727: dataIn1 = 32'd583
; 
32'd13728: dataIn1 = 32'd616
; 
32'd13729: dataIn1 = 32'd635
; 
32'd13730: dataIn1 = 32'd637
; 
32'd13731: dataIn1 = 32'd487
; 
32'd13732: dataIn1 = 32'd555
; 
32'd13733: dataIn1 = 32'd556
; 
32'd13734: dataIn1 = 32'd617
; 
32'd13735: dataIn1 = 32'd712
; 
32'd13736: dataIn1 = 32'd476
; 
32'd13737: dataIn1 = 32'd557
; 
32'd13738: dataIn1 = 32'd558
; 
32'd13739: dataIn1 = 32'd618
; 
32'd13740: dataIn1 = 32'd636
; 
32'd13741: dataIn1 = 32'd668
; 
32'd13742: dataIn1 = 32'd674
; 
32'd13743: dataIn1 = 32'd505
; 
32'd13744: dataIn1 = 32'd547
; 
32'd13745: dataIn1 = 32'd569
; 
32'd13746: dataIn1 = 32'd619
; 
32'd13747: dataIn1 = 32'd622
; 
32'd13748: dataIn1 = 32'd644
; 
32'd13749: dataIn1 = 32'd514
; 
32'd13750: dataIn1 = 32'd564
; 
32'd13751: dataIn1 = 32'd595
; 
32'd13752: dataIn1 = 32'd620
; 
32'd13753: dataIn1 = 32'd652
; 
32'd13754: dataIn1 = 32'd672
; 
32'd13755: dataIn1 = 32'd703
; 
32'd13756: dataIn1 = 32'd499
; 
32'd13757: dataIn1 = 32'd522
; 
32'd13758: dataIn1 = 32'd529
; 
32'd13759: dataIn1 = 32'd621
; 
32'd13760: dataIn1 = 32'd640
; 
32'd13761: dataIn1 = 32'd696
; 
32'd13762: dataIn1 = 32'd704
; 
32'd13763: dataIn1 = 32'd543
; 
32'd13764: dataIn1 = 32'd596
; 
32'd13765: dataIn1 = 32'd619
; 
32'd13766: dataIn1 = 32'd622
; 
32'd13767: dataIn1 = 32'd664
; 
32'd13768: dataIn1 = 32'd706
; 
32'd13769: dataIn1 = 32'd537
; 
32'd13770: dataIn1 = 32'd570
; 
32'd13771: dataIn1 = 32'd575
; 
32'd13772: dataIn1 = 32'd623
; 
32'd13773: dataIn1 = 32'd651
; 
32'd13774: dataIn1 = 32'd655
; 
32'd13775: dataIn1 = 32'd665
; 
32'd13776: dataIn1 = 32'd710
; 
32'd13777: dataIn1 = 32'd719
; 
32'd13778: dataIn1 = 32'd562
; 
32'd13779: dataIn1 = 32'd612
; 
32'd13780: dataIn1 = 32'd613
; 
32'd13781: dataIn1 = 32'd624
; 
32'd13782: dataIn1 = 32'd655
; 
32'd13783: dataIn1 = 32'd688
; 
32'd13784: dataIn1 = 32'd709
; 
32'd13785: dataIn1 = 32'd525
; 
32'd13786: dataIn1 = 32'd530
; 
32'd13787: dataIn1 = 32'd594
; 
32'd13788: dataIn1 = 32'd625
; 
32'd13789: dataIn1 = 32'd686
; 
32'd13790: dataIn1 = 32'd692
; 
32'd13791: dataIn1 = 32'd557
; 
32'd13792: dataIn1 = 32'd566
; 
32'd13793: dataIn1 = 32'd608
; 
32'd13794: dataIn1 = 32'd626
; 
32'd13795: dataIn1 = 32'd674
; 
32'd13796: dataIn1 = 32'd689
; 
32'd13797: dataIn1 = 32'd707
; 
32'd13798: dataIn1 = 32'd711
; 
32'd13799: dataIn1 = 32'd543
; 
32'd13800: dataIn1 = 32'd561
; 
32'd13801: dataIn1 = 32'd592
; 
32'd13802: dataIn1 = 32'd627
; 
32'd13803: dataIn1 = 32'd522
; 
32'd13804: dataIn1 = 32'd524
; 
32'd13805: dataIn1 = 32'd578
; 
32'd13806: dataIn1 = 32'd628
; 
32'd13807: dataIn1 = 32'd645
; 
32'd13808: dataIn1 = 32'd676
; 
32'd13809: dataIn1 = 32'd524
; 
32'd13810: dataIn1 = 32'd530
; 
32'd13811: dataIn1 = 32'd591
; 
32'd13812: dataIn1 = 32'd629
; 
32'd13813: dataIn1 = 32'd670
; 
32'd13814: dataIn1 = 32'd686
; 
32'd13815: dataIn1 = 32'd534
; 
32'd13816: dataIn1 = 32'd560
; 
32'd13817: dataIn1 = 32'd590
; 
32'd13818: dataIn1 = 32'd630
; 
32'd13819: dataIn1 = 32'd650
; 
32'd13820: dataIn1 = 32'd533
; 
32'd13821: dataIn1 = 32'd572
; 
32'd13822: dataIn1 = 32'd584
; 
32'd13823: dataIn1 = 32'd631
; 
32'd13824: dataIn1 = 32'd680
; 
32'd13825: dataIn1 = 32'd712
; 
32'd13826: dataIn1 = 32'd552
; 
32'd13827: dataIn1 = 32'd582
; 
32'd13828: dataIn1 = 32'd588
; 
32'd13829: dataIn1 = 32'd632
; 
32'd13830: dataIn1 = 32'd682
; 
32'd13831: dataIn1 = 32'd685
; 
32'd13832: dataIn1 = 32'd717
; 
32'd13833: dataIn1 = 32'd742
; 
32'd13834: dataIn1 = 32'd754
; 
32'd13835: dataIn1 = 32'd533
; 
32'd13836: dataIn1 = 32'd576
; 
32'd13837: dataIn1 = 32'd606
; 
32'd13838: dataIn1 = 32'd633
; 
32'd13839: dataIn1 = 32'd667
; 
32'd13840: dataIn1 = 32'd680
; 
32'd13841: dataIn1 = 32'd514
; 
32'd13842: dataIn1 = 32'd584
; 
32'd13843: dataIn1 = 32'd585
; 
32'd13844: dataIn1 = 32'd634
; 
32'd13845: dataIn1 = 32'd672
; 
32'd13846: dataIn1 = 32'd698
; 
32'd13847: dataIn1 = 32'd577
; 
32'd13848: dataIn1 = 32'd615
; 
32'd13849: dataIn1 = 32'd616
; 
32'd13850: dataIn1 = 32'd635
; 
32'd13851: dataIn1 = 32'd656
; 
32'd13852: dataIn1 = 32'd669
; 
32'd13853: dataIn1 = 32'd724
; 
32'd13854: dataIn1 = 32'd725
; 
32'd13855: dataIn1 = 32'd731
; 
32'd13856: dataIn1 = 32'd739
; 
32'd13857: dataIn1 = 32'd743
; 
32'd13858: dataIn1 = 32'd788
; 
32'd13859: dataIn1 = 32'd832
; 
32'd13860: dataIn1 = 32'd545
; 
32'd13861: dataIn1 = 32'd602
; 
32'd13862: dataIn1 = 32'd618
; 
32'd13863: dataIn1 = 32'd636
; 
32'd13864: dataIn1 = 32'd668
; 
32'd13865: dataIn1 = 32'd677
; 
32'd13866: dataIn1 = 32'd729
; 
32'd13867: dataIn1 = 32'd581
; 
32'd13868: dataIn1 = 32'd583
; 
32'd13869: dataIn1 = 32'd616
; 
32'd13870: dataIn1 = 32'd637
; 
32'd13871: dataIn1 = 32'd724
; 
32'd13872: dataIn1 = 32'd545
; 
32'd13873: dataIn1 = 32'd587
; 
32'd13874: dataIn1 = 32'd602
; 
32'd13875: dataIn1 = 32'd638
; 
32'd13876: dataIn1 = 32'd677
; 
32'd13877: dataIn1 = 32'd681
; 
32'd13878: dataIn1 = 32'd708
; 
32'd13879: dataIn1 = 32'd744
; 
32'd13880: dataIn1 = 32'd553
; 
32'd13881: dataIn1 = 32'd587
; 
32'd13882: dataIn1 = 32'd611
; 
32'd13883: dataIn1 = 32'd639
; 
32'd13884: dataIn1 = 32'd684
; 
32'd13885: dataIn1 = 32'd708
; 
32'd13886: dataIn1 = 32'd529
; 
32'd13887: dataIn1 = 32'd586
; 
32'd13888: dataIn1 = 32'd621
; 
32'd13889: dataIn1 = 32'd640
; 
32'd13890: dataIn1 = 32'd679
; 
32'd13891: dataIn1 = 32'd563
; 
32'd13892: dataIn1 = 32'd585
; 
32'd13893: dataIn1 = 32'd587
; 
32'd13894: dataIn1 = 32'd641
; 
32'd13895: dataIn1 = 32'd681
; 
32'd13896: dataIn1 = 32'd684
; 
32'd13897: dataIn1 = 32'd568
; 
32'd13898: dataIn1 = 32'd579
; 
32'd13899: dataIn1 = 32'd586
; 
32'd13900: dataIn1 = 32'd642
; 
32'd13901: dataIn1 = 32'd662
; 
32'd13902: dataIn1 = 32'd695
; 
32'd13903: dataIn1 = 32'd567
; 
32'd13904: dataIn1 = 32'd572
; 
32'd13905: dataIn1 = 32'd610
; 
32'd13906: dataIn1 = 32'd643
; 
32'd13907: dataIn1 = 32'd647
; 
32'd13908: dataIn1 = 32'd690
; 
32'd13909: dataIn1 = 32'd714
; 
32'd13910: dataIn1 = 32'd505
; 
32'd13911: dataIn1 = 32'd578
; 
32'd13912: dataIn1 = 32'd619
; 
32'd13913: dataIn1 = 32'd644
; 
32'd13914: dataIn1 = 32'd673
; 
32'd13915: dataIn1 = 32'd522
; 
32'd13916: dataIn1 = 32'd524
; 
32'd13917: dataIn1 = 32'd628
; 
32'd13918: dataIn1 = 32'd645
; 
32'd13919: dataIn1 = 32'd670
; 
32'd13920: dataIn1 = 32'd678
; 
32'd13921: dataIn1 = 32'd745
; 
32'd13922: dataIn1 = 32'd525
; 
32'd13923: dataIn1 = 32'd552
; 
32'd13924: dataIn1 = 32'd575
; 
32'd13925: dataIn1 = 32'd646
; 
32'd13926: dataIn1 = 32'd682
; 
32'd13927: dataIn1 = 32'd552
; 
32'd13928: dataIn1 = 32'd605
; 
32'd13929: dataIn1 = 32'd643
; 
32'd13930: dataIn1 = 32'd647
; 
32'd13931: dataIn1 = 32'd690
; 
32'd13932: dataIn1 = 32'd692
; 
32'd13933: dataIn1 = 32'd705
; 
32'd13934: dataIn1 = 32'd715
; 
32'd13935: dataIn1 = 32'd746
; 
32'd13936: dataIn1 = 32'd553
; 
32'd13937: dataIn1 = 32'd612
; 
32'd13938: dataIn1 = 32'd614
; 
32'd13939: dataIn1 = 32'd648
; 
32'd13940: dataIn1 = 32'd691
; 
32'd13941: dataIn1 = 32'd720
; 
32'd13942: dataIn1 = 32'd728
; 
32'd13943: dataIn1 = 32'd747
; 
32'd13944: dataIn1 = 32'd768
; 
32'd13945: dataIn1 = 32'd557
; 
32'd13946: dataIn1 = 32'd574
; 
32'd13947: dataIn1 = 32'd589
; 
32'd13948: dataIn1 = 32'd649
; 
32'd13949: dataIn1 = 32'd650
; 
32'd13950: dataIn1 = 32'd689
; 
32'd13951: dataIn1 = 32'd560
; 
32'd13952: dataIn1 = 32'd630
; 
32'd13953: dataIn1 = 32'd649
; 
32'd13954: dataIn1 = 32'd650
; 
32'd13955: dataIn1 = 32'd725
; 
32'd13956: dataIn1 = 32'd740
; 
32'd13957: dataIn1 = 32'd741
; 
32'd13958: dataIn1 = 32'd748
; 
32'd13959: dataIn1 = 32'd755
; 
32'd13960: dataIn1 = 32'd786
; 
32'd13961: dataIn1 = 32'd562
; 
32'd13962: dataIn1 = 32'd575
; 
32'd13963: dataIn1 = 32'd623
; 
32'd13964: dataIn1 = 32'd651
; 
32'd13965: dataIn1 = 32'd688
; 
32'd13966: dataIn1 = 32'd719
; 
32'd13967: dataIn1 = 32'd733
; 
32'd13968: dataIn1 = 32'd522
; 
32'd13969: dataIn1 = 32'd564
; 
32'd13970: dataIn1 = 32'd620
; 
32'd13971: dataIn1 = 32'd652
; 
32'd13972: dataIn1 = 32'd745
; 
32'd13973: dataIn1 = 32'd749
; 
32'd13974: dataIn1 = 32'd759
; 
32'd13975: dataIn1 = 32'd565
; 
32'd13976: dataIn1 = 32'd568
; 
32'd13977: dataIn1 = 32'd573
; 
32'd13978: dataIn1 = 32'd653
; 
32'd13979: dataIn1 = 32'd691
; 
32'd13980: dataIn1 = 32'd565
; 
32'd13981: dataIn1 = 32'd568
; 
32'd13982: dataIn1 = 32'd597
; 
32'd13983: dataIn1 = 32'd654
; 
32'd13984: dataIn1 = 32'd687
; 
32'd13985: dataIn1 = 32'd573
; 
32'd13986: dataIn1 = 32'd623
; 
32'd13987: dataIn1 = 32'd624
; 
32'd13988: dataIn1 = 32'd655
; 
32'd13989: dataIn1 = 32'd709
; 
32'd13990: dataIn1 = 32'd710
; 
32'd13991: dataIn1 = 32'd721
; 
32'd13992: dataIn1 = 32'd750
; 
32'd13993: dataIn1 = 32'd577
; 
32'd13994: dataIn1 = 32'd595
; 
32'd13995: dataIn1 = 32'd635
; 
32'd13996: dataIn1 = 32'd656
; 
32'd13997: dataIn1 = 32'd696
; 
32'd13998: dataIn1 = 32'd578
; 
32'd13999: dataIn1 = 32'd594
; 
32'd14000: dataIn1 = 32'd596
; 
32'd14001: dataIn1 = 32'd657
; 
32'd14002: dataIn1 = 32'd697
; 
32'd14003: dataIn1 = 32'd705
; 
32'd14004: dataIn1 = 32'd726
; 
32'd14005: dataIn1 = 32'd583
; 
32'd14006: dataIn1 = 32'd592
; 
32'd14007: dataIn1 = 32'd615
; 
32'd14008: dataIn1 = 32'd658
; 
32'd14009: dataIn1 = 32'd565
; 
32'd14010: dataIn1 = 32'd597
; 
32'd14011: dataIn1 = 32'd607
; 
32'd14012: dataIn1 = 32'd659
; 
32'd14013: dataIn1 = 32'd673
; 
32'd14014: dataIn1 = 32'd694
; 
32'd14015: dataIn1 = 32'd707
; 
32'd14016: dataIn1 = 32'd736
; 
32'd14017: dataIn1 = 32'd751
; 
32'd14018: dataIn1 = 32'd763
; 
32'd14019: dataIn1 = 32'd793
; 
32'd14020: dataIn1 = 32'd537
; 
32'd14021: dataIn1 = 32'd540
; 
32'd14022: dataIn1 = 32'd598
; 
32'd14023: dataIn1 = 32'd660
; 
32'd14024: dataIn1 = 32'd701
; 
32'd14025: dataIn1 = 32'd558
; 
32'd14026: dataIn1 = 32'd598
; 
32'd14027: dataIn1 = 32'd599
; 
32'd14028: dataIn1 = 32'd661
; 
32'd14029: dataIn1 = 32'd674
; 
32'd14030: dataIn1 = 32'd685
; 
32'd14031: dataIn1 = 32'd597
; 
32'd14032: dataIn1 = 32'd604
; 
32'd14033: dataIn1 = 32'd642
; 
32'd14034: dataIn1 = 32'd662
; 
32'd14035: dataIn1 = 32'd679
; 
32'd14036: dataIn1 = 32'd751
; 
32'd14037: dataIn1 = 32'd752
; 
32'd14038: dataIn1 = 32'd771
; 
32'd14039: dataIn1 = 32'd796
; 
32'd14040: dataIn1 = 32'd592
; 
32'd14041: dataIn1 = 32'd596
; 
32'd14042: dataIn1 = 32'd605
; 
32'd14043: dataIn1 = 32'd663
; 
32'd14044: dataIn1 = 32'd683
; 
32'd14045: dataIn1 = 32'd753
; 
32'd14046: dataIn1 = 32'd592
; 
32'd14047: dataIn1 = 32'd607
; 
32'd14048: dataIn1 = 32'd622
; 
32'd14049: dataIn1 = 32'd664
; 
32'd14050: dataIn1 = 32'd741
; 
32'd14051: dataIn1 = 32'd753
; 
32'd14052: dataIn1 = 32'd765
; 
32'd14053: dataIn1 = 32'd766
; 
32'd14054: dataIn1 = 32'd565
; 
32'd14055: dataIn1 = 32'd608
; 
32'd14056: dataIn1 = 32'd623
; 
32'd14057: dataIn1 = 32'd665
; 
32'd14058: dataIn1 = 32'd694
; 
32'd14059: dataIn1 = 32'd710
; 
32'd14060: dataIn1 = 32'd544
; 
32'd14061: dataIn1 = 32'd609
; 
32'd14062: dataIn1 = 32'd614
; 
32'd14063: dataIn1 = 32'd666
; 
32'd14064: dataIn1 = 32'd700
; 
32'd14065: dataIn1 = 32'd602
; 
32'd14066: dataIn1 = 32'd610
; 
32'd14067: dataIn1 = 32'd633
; 
32'd14068: dataIn1 = 32'd667
; 
32'd14069: dataIn1 = 32'd675
; 
32'd14070: dataIn1 = 32'd742
; 
32'd14071: dataIn1 = 32'd588
; 
32'd14072: dataIn1 = 32'd618
; 
32'd14073: dataIn1 = 32'd636
; 
32'd14074: dataIn1 = 32'd668
; 
32'd14075: dataIn1 = 32'd729
; 
32'd14076: dataIn1 = 32'd754
; 
32'd14077: dataIn1 = 32'd590
; 
32'd14078: dataIn1 = 32'd615
; 
32'd14079: dataIn1 = 32'd635
; 
32'd14080: dataIn1 = 32'd669
; 
32'd14081: dataIn1 = 32'd716
; 
32'd14082: dataIn1 = 32'd730
; 
32'd14083: dataIn1 = 32'd755
; 
32'd14084: dataIn1 = 32'd578
; 
32'd14085: dataIn1 = 32'd629
; 
32'd14086: dataIn1 = 32'd645
; 
32'd14087: dataIn1 = 32'd670
; 
32'd14088: dataIn1 = 32'd718
; 
32'd14089: dataIn1 = 32'd727
; 
32'd14090: dataIn1 = 32'd770
; 
32'd14091: dataIn1 = 32'd578
; 
32'd14092: dataIn1 = 32'd597
; 
32'd14093: dataIn1 = 32'd604
; 
32'd14094: dataIn1 = 32'd671
; 
32'd14095: dataIn1 = 32'd676
; 
32'd14096: dataIn1 = 32'd727
; 
32'd14097: dataIn1 = 32'd752
; 
32'd14098: dataIn1 = 32'd777
; 
32'd14099: dataIn1 = 32'd584
; 
32'd14100: dataIn1 = 32'd620
; 
32'd14101: dataIn1 = 32'd634
; 
32'd14102: dataIn1 = 32'd672
; 
32'd14103: dataIn1 = 32'd712
; 
32'd14104: dataIn1 = 32'd735
; 
32'd14105: dataIn1 = 32'd739
; 
32'd14106: dataIn1 = 32'd756
; 
32'd14107: dataIn1 = 32'd826
; 
32'd14108: dataIn1 = 32'd597
; 
32'd14109: dataIn1 = 32'd644
; 
32'd14110: dataIn1 = 32'd659
; 
32'd14111: dataIn1 = 32'd673
; 
32'd14112: dataIn1 = 32'd697
; 
32'd14113: dataIn1 = 32'd706
; 
32'd14114: dataIn1 = 32'd751
; 
32'd14115: dataIn1 = 32'd777
; 
32'd14116: dataIn1 = 32'd618
; 
32'd14117: dataIn1 = 32'd626
; 
32'd14118: dataIn1 = 32'd661
; 
32'd14119: dataIn1 = 32'd674
; 
32'd14120: dataIn1 = 32'd701
; 
32'd14121: dataIn1 = 32'd754
; 
32'd14122: dataIn1 = 32'd757
; 
32'd14123: dataIn1 = 32'd769
; 
32'd14124: dataIn1 = 32'd772
; 
32'd14125: dataIn1 = 32'd785
; 
32'd14126: dataIn1 = 32'd602
; 
32'd14127: dataIn1 = 32'd606
; 
32'd14128: dataIn1 = 32'd667
; 
32'd14129: dataIn1 = 32'd675
; 
32'd14130: dataIn1 = 32'd756
; 
32'd14131: dataIn1 = 32'd604
; 
32'd14132: dataIn1 = 32'd628
; 
32'd14133: dataIn1 = 32'd671
; 
32'd14134: dataIn1 = 32'd676
; 
32'd14135: dataIn1 = 32'd589
; 
32'd14136: dataIn1 = 32'd636
; 
32'd14137: dataIn1 = 32'd638
; 
32'd14138: dataIn1 = 32'd677
; 
32'd14139: dataIn1 = 32'd693
; 
32'd14140: dataIn1 = 32'd758
; 
32'd14141: dataIn1 = 32'd773
; 
32'd14142: dataIn1 = 32'd799
; 
32'd14143: dataIn1 = 32'd804
; 
32'd14144: dataIn1 = 32'd591
; 
32'd14145: dataIn1 = 32'd601
; 
32'd14146: dataIn1 = 32'd645
; 
32'd14147: dataIn1 = 32'd678
; 
32'd14148: dataIn1 = 32'd703
; 
32'd14149: dataIn1 = 32'd745
; 
32'd14150: dataIn1 = 32'd759
; 
32'd14151: dataIn1 = 32'd764
; 
32'd14152: dataIn1 = 32'd770
; 
32'd14153: dataIn1 = 32'd815
; 
32'd14154: dataIn1 = 32'd609
; 
32'd14155: dataIn1 = 32'd640
; 
32'd14156: dataIn1 = 32'd662
; 
32'd14157: dataIn1 = 32'd679
; 
32'd14158: dataIn1 = 32'd743
; 
32'd14159: dataIn1 = 32'd760
; 
32'd14160: dataIn1 = 32'd771
; 
32'd14161: dataIn1 = 32'd778
; 
32'd14162: dataIn1 = 32'd610
; 
32'd14163: dataIn1 = 32'd631
; 
32'd14164: dataIn1 = 32'd633
; 
32'd14165: dataIn1 = 32'd680
; 
32'd14166: dataIn1 = 32'd732
; 
32'd14167: dataIn1 = 32'd585
; 
32'd14168: dataIn1 = 32'd638
; 
32'd14169: dataIn1 = 32'd641
; 
32'd14170: dataIn1 = 32'd681
; 
32'd14171: dataIn1 = 32'd735
; 
32'd14172: dataIn1 = 32'd744
; 
32'd14173: dataIn1 = 32'd758
; 
32'd14174: dataIn1 = 32'd779
; 
32'd14175: dataIn1 = 32'd800
; 
32'd14176: dataIn1 = 32'd599
; 
32'd14177: dataIn1 = 32'd632
; 
32'd14178: dataIn1 = 32'd646
; 
32'd14179: dataIn1 = 32'd682
; 
32'd14180: dataIn1 = 32'd719
; 
32'd14181: dataIn1 = 32'd733
; 
32'd14182: dataIn1 = 32'd761
; 
32'd14183: dataIn1 = 32'd787
; 
32'd14184: dataIn1 = 32'd801
; 
32'd14185: dataIn1 = 32'd848
; 
32'd14186: dataIn1 = 32'd592
; 
32'd14187: dataIn1 = 32'd605
; 
32'd14188: dataIn1 = 32'd663
; 
32'd14189: dataIn1 = 32'd683
; 
32'd14190: dataIn1 = 32'd714
; 
32'd14191: dataIn1 = 32'd724
; 
32'd14192: dataIn1 = 32'd738
; 
32'd14193: dataIn1 = 32'd762
; 
32'd14194: dataIn1 = 32'd784
; 
32'd14195: dataIn1 = 32'd587
; 
32'd14196: dataIn1 = 32'd639
; 
32'd14197: dataIn1 = 32'd641
; 
32'd14198: dataIn1 = 32'd684
; 
32'd14199: dataIn1 = 32'd702
; 
32'd14200: dataIn1 = 32'd722
; 
32'd14201: dataIn1 = 32'd768
; 
32'd14202: dataIn1 = 32'd599
; 
32'd14203: dataIn1 = 32'd632
; 
32'd14204: dataIn1 = 32'd661
; 
32'd14205: dataIn1 = 32'd685
; 
32'd14206: dataIn1 = 32'd761
; 
32'd14207: dataIn1 = 32'd591
; 
32'd14208: dataIn1 = 32'd625
; 
32'd14209: dataIn1 = 32'd629
; 
32'd14210: dataIn1 = 32'd686
; 
32'd14211: dataIn1 = 32'd718
; 
32'd14212: dataIn1 = 32'd734
; 
32'd14213: dataIn1 = 32'd770
; 
32'd14214: dataIn1 = 32'd565
; 
32'd14215: dataIn1 = 32'd568
; 
32'd14216: dataIn1 = 32'd654
; 
32'd14217: dataIn1 = 32'd687
; 
32'd14218: dataIn1 = 32'd695
; 
32'd14219: dataIn1 = 32'd763
; 
32'd14220: dataIn1 = 32'd802
; 
32'd14221: dataIn1 = 32'd601
; 
32'd14222: dataIn1 = 32'd624
; 
32'd14223: dataIn1 = 32'd651
; 
32'd14224: dataIn1 = 32'd688
; 
32'd14225: dataIn1 = 32'd713
; 
32'd14226: dataIn1 = 32'd721
; 
32'd14227: dataIn1 = 32'd723
; 
32'd14228: dataIn1 = 32'd764
; 
32'd14229: dataIn1 = 32'd607
; 
32'd14230: dataIn1 = 32'd626
; 
32'd14231: dataIn1 = 32'd649
; 
32'd14232: dataIn1 = 32'd689
; 
32'd14233: dataIn1 = 32'd693
; 
32'd14234: dataIn1 = 32'd737
; 
32'd14235: dataIn1 = 32'd748
; 
32'd14236: dataIn1 = 32'd765
; 
32'd14237: dataIn1 = 32'd769
; 
32'd14238: dataIn1 = 32'd782
; 
32'd14239: dataIn1 = 32'd803
; 
32'd14240: dataIn1 = 32'd610
; 
32'd14241: dataIn1 = 32'd643
; 
32'd14242: dataIn1 = 32'd647
; 
32'd14243: dataIn1 = 32'd690
; 
32'd14244: dataIn1 = 32'd717
; 
32'd14245: dataIn1 = 32'd732
; 
32'd14246: dataIn1 = 32'd746
; 
32'd14247: dataIn1 = 32'd568
; 
32'd14248: dataIn1 = 32'd648
; 
32'd14249: dataIn1 = 32'd653
; 
32'd14250: dataIn1 = 32'd691
; 
32'd14251: dataIn1 = 32'd720
; 
32'd14252: dataIn1 = 32'd552
; 
32'd14253: dataIn1 = 32'd625
; 
32'd14254: dataIn1 = 32'd647
; 
32'd14255: dataIn1 = 32'd692
; 
32'd14256: dataIn1 = 32'd718
; 
32'd14257: dataIn1 = 32'd794
; 
32'd14258: dataIn1 = 32'd801
; 
32'd14259: dataIn1 = 32'd557
; 
32'd14260: dataIn1 = 32'd677
; 
32'd14261: dataIn1 = 32'd689
; 
32'd14262: dataIn1 = 32'd693
; 
32'd14263: dataIn1 = 32'd740
; 
32'd14264: dataIn1 = 32'd757
; 
32'd14265: dataIn1 = 32'd769
; 
32'd14266: dataIn1 = 32'd804
; 
32'd14267: dataIn1 = 32'd565
; 
32'd14268: dataIn1 = 32'd659
; 
32'd14269: dataIn1 = 32'd665
; 
32'd14270: dataIn1 = 32'd694
; 
32'd14271: dataIn1 = 32'd763
; 
32'd14272: dataIn1 = 32'd774
; 
32'd14273: dataIn1 = 32'd568
; 
32'd14274: dataIn1 = 32'd642
; 
32'd14275: dataIn1 = 32'd687
; 
32'd14276: dataIn1 = 32'd695
; 
32'd14277: dataIn1 = 32'd747
; 
32'd14278: dataIn1 = 32'd577
; 
32'd14279: dataIn1 = 32'd621
; 
32'd14280: dataIn1 = 32'd656
; 
32'd14281: dataIn1 = 32'd696
; 
32'd14282: dataIn1 = 32'd704
; 
32'd14283: dataIn1 = 32'd578
; 
32'd14284: dataIn1 = 32'd657
; 
32'd14285: dataIn1 = 32'd673
; 
32'd14286: dataIn1 = 32'd697
; 
32'd14287: dataIn1 = 32'd726
; 
32'd14288: dataIn1 = 32'd727
; 
32'd14289: dataIn1 = 32'd790
; 
32'd14290: dataIn1 = 32'd805
; 
32'd14291: dataIn1 = 32'd585
; 
32'd14292: dataIn1 = 32'd600
; 
32'd14293: dataIn1 = 32'd634
; 
32'd14294: dataIn1 = 32'd698
; 
32'd14295: dataIn1 = 32'd735
; 
32'd14296: dataIn1 = 32'd589
; 
32'd14297: dataIn1 = 32'd590
; 
32'd14298: dataIn1 = 32'd611
; 
32'd14299: dataIn1 = 32'd699
; 
32'd14300: dataIn1 = 32'd700
; 
32'd14301: dataIn1 = 32'd716
; 
32'd14302: dataIn1 = 32'd773
; 
32'd14303: dataIn1 = 32'd590
; 
32'd14304: dataIn1 = 32'd666
; 
32'd14305: dataIn1 = 32'd699
; 
32'd14306: dataIn1 = 32'd700
; 
32'd14307: dataIn1 = 32'd728
; 
32'd14308: dataIn1 = 32'd730
; 
32'd14309: dataIn1 = 32'd599
; 
32'd14310: dataIn1 = 32'd660
; 
32'd14311: dataIn1 = 32'd674
; 
32'd14312: dataIn1 = 32'd701
; 
32'd14313: dataIn1 = 32'd711
; 
32'd14314: dataIn1 = 32'd761
; 
32'd14315: dataIn1 = 32'd772
; 
32'd14316: dataIn1 = 32'd776
; 
32'd14317: dataIn1 = 32'd600
; 
32'd14318: dataIn1 = 32'd612
; 
32'd14319: dataIn1 = 32'd684
; 
32'd14320: dataIn1 = 32'd702
; 
32'd14321: dataIn1 = 32'd722
; 
32'd14322: dataIn1 = 32'd601
; 
32'd14323: dataIn1 = 32'd620
; 
32'd14324: dataIn1 = 32'd678
; 
32'd14325: dataIn1 = 32'd703
; 
32'd14326: dataIn1 = 32'd713
; 
32'd14327: dataIn1 = 32'd759
; 
32'd14328: dataIn1 = 32'd604
; 
32'd14329: dataIn1 = 32'd621
; 
32'd14330: dataIn1 = 32'd696
; 
32'd14331: dataIn1 = 32'd704
; 
32'd14332: dataIn1 = 32'd749
; 
32'd14333: dataIn1 = 32'd752
; 
32'd14334: dataIn1 = 32'd760
; 
32'd14335: dataIn1 = 32'd605
; 
32'd14336: dataIn1 = 32'd647
; 
32'd14337: dataIn1 = 32'd657
; 
32'd14338: dataIn1 = 32'd705
; 
32'd14339: dataIn1 = 32'd715
; 
32'd14340: dataIn1 = 32'd738
; 
32'd14341: dataIn1 = 32'd794
; 
32'd14342: dataIn1 = 32'd607
; 
32'd14343: dataIn1 = 32'd622
; 
32'd14344: dataIn1 = 32'd673
; 
32'd14345: dataIn1 = 32'd706
; 
32'd14346: dataIn1 = 32'd726
; 
32'd14347: dataIn1 = 32'd736
; 
32'd14348: dataIn1 = 32'd753
; 
32'd14349: dataIn1 = 32'd766
; 
32'd14350: dataIn1 = 32'd790
; 
32'd14351: dataIn1 = 32'd608
; 
32'd14352: dataIn1 = 32'd626
; 
32'd14353: dataIn1 = 32'd659
; 
32'd14354: dataIn1 = 32'd707
; 
32'd14355: dataIn1 = 32'd711
; 
32'd14356: dataIn1 = 32'd611
; 
32'd14357: dataIn1 = 32'd638
; 
32'd14358: dataIn1 = 32'd639
; 
32'd14359: dataIn1 = 32'd708
; 
32'd14360: dataIn1 = 32'd728
; 
32'd14361: dataIn1 = 32'd758
; 
32'd14362: dataIn1 = 32'd612
; 
32'd14363: dataIn1 = 32'd624
; 
32'd14364: dataIn1 = 32'd655
; 
32'd14365: dataIn1 = 32'd709
; 
32'd14366: dataIn1 = 32'd720
; 
32'd14367: dataIn1 = 32'd721
; 
32'd14368: dataIn1 = 32'd722
; 
32'd14369: dataIn1 = 32'd767
; 
32'd14370: dataIn1 = 32'd623
; 
32'd14371: dataIn1 = 32'd655
; 
32'd14372: dataIn1 = 32'd665
; 
32'd14373: dataIn1 = 32'd710
; 
32'd14374: dataIn1 = 32'd750
; 
32'd14375: dataIn1 = 32'd774
; 
32'd14376: dataIn1 = 32'd776
; 
32'd14377: dataIn1 = 32'd626
; 
32'd14378: dataIn1 = 32'd701
; 
32'd14379: dataIn1 = 32'd707
; 
32'd14380: dataIn1 = 32'd711
; 
32'd14381: dataIn1 = 32'd737
; 
32'd14382: dataIn1 = 32'd772
; 
32'd14383: dataIn1 = 32'd774
; 
32'd14384: dataIn1 = 32'd617
; 
32'd14385: dataIn1 = 32'd631
; 
32'd14386: dataIn1 = 32'd672
; 
32'd14387: dataIn1 = 32'd712
; 
32'd14388: dataIn1 = 32'd731
; 
32'd14389: dataIn1 = 32'd739
; 
32'd14390: dataIn1 = 32'd600
; 
32'd14391: dataIn1 = 32'd688
; 
32'd14392: dataIn1 = 32'd703
; 
32'd14393: dataIn1 = 32'd713
; 
32'd14394: dataIn1 = 32'd723
; 
32'd14395: dataIn1 = 32'd775
; 
32'd14396: dataIn1 = 32'd605
; 
32'd14397: dataIn1 = 32'd643
; 
32'd14398: dataIn1 = 32'd683
; 
32'd14399: dataIn1 = 32'd714
; 
32'd14400: dataIn1 = 32'd715
; 
32'd14401: dataIn1 = 32'd732
; 
32'd14402: dataIn1 = 32'd647
; 
32'd14403: dataIn1 = 32'd705
; 
32'd14404: dataIn1 = 32'd714
; 
32'd14405: dataIn1 = 32'd715
; 
32'd14406: dataIn1 = 32'd738
; 
32'd14407: dataIn1 = 32'd791
; 
32'd14408: dataIn1 = 32'd806
; 
32'd14409: dataIn1 = 32'd590
; 
32'd14410: dataIn1 = 32'd669
; 
32'd14411: dataIn1 = 32'd699
; 
32'd14412: dataIn1 = 32'd716
; 
32'd14413: dataIn1 = 32'd730
; 
32'd14414: dataIn1 = 32'd552
; 
32'd14415: dataIn1 = 32'd632
; 
32'd14416: dataIn1 = 32'd690
; 
32'd14417: dataIn1 = 32'd717
; 
32'd14418: dataIn1 = 32'd746
; 
32'd14419: dataIn1 = 32'd787
; 
32'd14420: dataIn1 = 32'd670
; 
32'd14421: dataIn1 = 32'd686
; 
32'd14422: dataIn1 = 32'd692
; 
32'd14423: dataIn1 = 32'd718
; 
32'd14424: dataIn1 = 32'd818
; 
32'd14425: dataIn1 = 32'd871
; 
32'd14426: dataIn1 = 32'd623
; 
32'd14427: dataIn1 = 32'd651
; 
32'd14428: dataIn1 = 32'd682
; 
32'd14429: dataIn1 = 32'd719
; 
32'd14430: dataIn1 = 32'd733
; 
32'd14431: dataIn1 = 32'd776
; 
32'd14432: dataIn1 = 32'd648
; 
32'd14433: dataIn1 = 32'd691
; 
32'd14434: dataIn1 = 32'd709
; 
32'd14435: dataIn1 = 32'd720
; 
32'd14436: dataIn1 = 32'd747
; 
32'd14437: dataIn1 = 32'd750
; 
32'd14438: dataIn1 = 32'd780
; 
32'd14439: dataIn1 = 32'd655
; 
32'd14440: dataIn1 = 32'd688
; 
32'd14441: dataIn1 = 32'd709
; 
32'd14442: dataIn1 = 32'd721
; 
32'd14443: dataIn1 = 32'd783
; 
32'd14444: dataIn1 = 32'd807
; 
32'd14445: dataIn1 = 32'd684
; 
32'd14446: dataIn1 = 32'd702
; 
32'd14447: dataIn1 = 32'd709
; 
32'd14448: dataIn1 = 32'd722
; 
32'd14449: dataIn1 = 32'd767
; 
32'd14450: dataIn1 = 32'd768
; 
32'd14451: dataIn1 = 32'd600
; 
32'd14452: dataIn1 = 32'd688
; 
32'd14453: dataIn1 = 32'd713
; 
32'd14454: dataIn1 = 32'd723
; 
32'd14455: dataIn1 = 32'd767
; 
32'd14456: dataIn1 = 32'd775
; 
32'd14457: dataIn1 = 32'd635
; 
32'd14458: dataIn1 = 32'd637
; 
32'd14459: dataIn1 = 32'd683
; 
32'd14460: dataIn1 = 32'd724
; 
32'd14461: dataIn1 = 32'd725
; 
32'd14462: dataIn1 = 32'd731
; 
32'd14463: dataIn1 = 32'd784
; 
32'd14464: dataIn1 = 32'd635
; 
32'd14465: dataIn1 = 32'd650
; 
32'd14466: dataIn1 = 32'd724
; 
32'd14467: dataIn1 = 32'd725
; 
32'd14468: dataIn1 = 32'd755
; 
32'd14469: dataIn1 = 32'd784
; 
32'd14470: dataIn1 = 32'd786
; 
32'd14471: dataIn1 = 32'd808
; 
32'd14472: dataIn1 = 32'd843
; 
32'd14473: dataIn1 = 32'd657
; 
32'd14474: dataIn1 = 32'd697
; 
32'd14475: dataIn1 = 32'd706
; 
32'd14476: dataIn1 = 32'd726
; 
32'd14477: dataIn1 = 32'd790
; 
32'd14478: dataIn1 = 32'd805
; 
32'd14479: dataIn1 = 32'd809
; 
32'd14480: dataIn1 = 32'd670
; 
32'd14481: dataIn1 = 32'd671
; 
32'd14482: dataIn1 = 32'd697
; 
32'd14483: dataIn1 = 32'd727
; 
32'd14484: dataIn1 = 32'd795
; 
32'd14485: dataIn1 = 32'd818
; 
32'd14486: dataIn1 = 32'd850
; 
32'd14487: dataIn1 = 32'd861
; 
32'd14488: dataIn1 = 32'd648
; 
32'd14489: dataIn1 = 32'd700
; 
32'd14490: dataIn1 = 32'd708
; 
32'd14491: dataIn1 = 32'd728
; 
32'd14492: dataIn1 = 32'd773
; 
32'd14493: dataIn1 = 32'd830
; 
32'd14494: dataIn1 = 32'd853
; 
32'd14495: dataIn1 = 32'd602
; 
32'd14496: dataIn1 = 32'd636
; 
32'd14497: dataIn1 = 32'd668
; 
32'd14498: dataIn1 = 32'd729
; 
32'd14499: dataIn1 = 32'd742
; 
32'd14500: dataIn1 = 32'd757
; 
32'd14501: dataIn1 = 32'd799
; 
32'd14502: dataIn1 = 32'd669
; 
32'd14503: dataIn1 = 32'd700
; 
32'd14504: dataIn1 = 32'd716
; 
32'd14505: dataIn1 = 32'd730
; 
32'd14506: dataIn1 = 32'd743
; 
32'd14507: dataIn1 = 32'd778
; 
32'd14508: dataIn1 = 32'd810
; 
32'd14509: dataIn1 = 32'd830
; 
32'd14510: dataIn1 = 32'd847
; 
32'd14511: dataIn1 = 32'd635
; 
32'd14512: dataIn1 = 32'd712
; 
32'd14513: dataIn1 = 32'd724
; 
32'd14514: dataIn1 = 32'd731
; 
32'd14515: dataIn1 = 32'd756
; 
32'd14516: dataIn1 = 32'd792
; 
32'd14517: dataIn1 = 32'd808
; 
32'd14518: dataIn1 = 32'd826
; 
32'd14519: dataIn1 = 32'd851
; 
32'd14520: dataIn1 = 32'd858
; 
32'd14521: dataIn1 = 32'd680
; 
32'd14522: dataIn1 = 32'd690
; 
32'd14523: dataIn1 = 32'd714
; 
32'd14524: dataIn1 = 32'd732
; 
32'd14525: dataIn1 = 32'd791
; 
32'd14526: dataIn1 = 32'd792
; 
32'd14527: dataIn1 = 32'd651
; 
32'd14528: dataIn1 = 32'd682
; 
32'd14529: dataIn1 = 32'd719
; 
32'd14530: dataIn1 = 32'd733
; 
32'd14531: dataIn1 = 32'd734
; 
32'd14532: dataIn1 = 32'd807
; 
32'd14533: dataIn1 = 32'd817
; 
32'd14534: dataIn1 = 32'd591
; 
32'd14535: dataIn1 = 32'd686
; 
32'd14536: dataIn1 = 32'd733
; 
32'd14537: dataIn1 = 32'd734
; 
32'd14538: dataIn1 = 32'd764
; 
32'd14539: dataIn1 = 32'd801
; 
32'd14540: dataIn1 = 32'd672
; 
32'd14541: dataIn1 = 32'd681
; 
32'd14542: dataIn1 = 32'd698
; 
32'd14543: dataIn1 = 32'd735
; 
32'd14544: dataIn1 = 32'd775
; 
32'd14545: dataIn1 = 32'd779
; 
32'd14546: dataIn1 = 32'd824
; 
32'd14547: dataIn1 = 32'd869
; 
32'd14548: dataIn1 = 32'd883
; 
32'd14549: dataIn1 = 32'd607
; 
32'd14550: dataIn1 = 32'd659
; 
32'd14551: dataIn1 = 32'd706
; 
32'd14552: dataIn1 = 32'd736
; 
32'd14553: dataIn1 = 32'd737
; 
32'd14554: dataIn1 = 32'd811
; 
32'd14555: dataIn1 = 32'd689
; 
32'd14556: dataIn1 = 32'd711
; 
32'd14557: dataIn1 = 32'd736
; 
32'd14558: dataIn1 = 32'd737
; 
32'd14559: dataIn1 = 32'd822
; 
32'd14560: dataIn1 = 32'd823
; 
32'd14561: dataIn1 = 32'd831
; 
32'd14562: dataIn1 = 32'd854
; 
32'd14563: dataIn1 = 32'd683
; 
32'd14564: dataIn1 = 32'd705
; 
32'd14565: dataIn1 = 32'd715
; 
32'd14566: dataIn1 = 32'd738
; 
32'd14567: dataIn1 = 32'd809
; 
32'd14568: dataIn1 = 32'd635
; 
32'd14569: dataIn1 = 32'd672
; 
32'd14570: dataIn1 = 32'd712
; 
32'd14571: dataIn1 = 32'd739
; 
32'd14572: dataIn1 = 32'd832
; 
32'd14573: dataIn1 = 32'd855
; 
32'd14574: dataIn1 = 32'd856
; 
32'd14575: dataIn1 = 32'd589
; 
32'd14576: dataIn1 = 32'd650
; 
32'd14577: dataIn1 = 32'd693
; 
32'd14578: dataIn1 = 32'd740
; 
32'd14579: dataIn1 = 32'd782
; 
32'd14580: dataIn1 = 32'd804
; 
32'd14581: dataIn1 = 32'd810
; 
32'd14582: dataIn1 = 32'd812
; 
32'd14583: dataIn1 = 32'd833
; 
32'd14584: dataIn1 = 32'd592
; 
32'd14585: dataIn1 = 32'd650
; 
32'd14586: dataIn1 = 32'd664
; 
32'd14587: dataIn1 = 32'd741
; 
32'd14588: dataIn1 = 32'd748
; 
32'd14589: dataIn1 = 32'd762
; 
32'd14590: dataIn1 = 32'd786
; 
32'd14591: dataIn1 = 32'd789
; 
32'd14592: dataIn1 = 32'd632
; 
32'd14593: dataIn1 = 32'd667
; 
32'd14594: dataIn1 = 32'd729
; 
32'd14595: dataIn1 = 32'd742
; 
32'd14596: dataIn1 = 32'd787
; 
32'd14597: dataIn1 = 32'd814
; 
32'd14598: dataIn1 = 32'd825
; 
32'd14599: dataIn1 = 32'd834
; 
32'd14600: dataIn1 = 32'd844
; 
32'd14601: dataIn1 = 32'd852
; 
32'd14602: dataIn1 = 32'd867
; 
32'd14603: dataIn1 = 32'd635
; 
32'd14604: dataIn1 = 32'd679
; 
32'd14605: dataIn1 = 32'd730
; 
32'd14606: dataIn1 = 32'd743
; 
32'd14607: dataIn1 = 32'd778
; 
32'd14608: dataIn1 = 32'd788
; 
32'd14609: dataIn1 = 32'd813
; 
32'd14610: dataIn1 = 32'd835
; 
32'd14611: dataIn1 = 32'd602
; 
32'd14612: dataIn1 = 32'd638
; 
32'd14613: dataIn1 = 32'd681
; 
32'd14614: dataIn1 = 32'd744
; 
32'd14615: dataIn1 = 32'd799
; 
32'd14616: dataIn1 = 32'd800
; 
32'd14617: dataIn1 = 32'd645
; 
32'd14618: dataIn1 = 32'd652
; 
32'd14619: dataIn1 = 32'd678
; 
32'd14620: dataIn1 = 32'd745
; 
32'd14621: dataIn1 = 32'd749
; 
32'd14622: dataIn1 = 32'd795
; 
32'd14623: dataIn1 = 32'd815
; 
32'd14624: dataIn1 = 32'd647
; 
32'd14625: dataIn1 = 32'd690
; 
32'd14626: dataIn1 = 32'd717
; 
32'd14627: dataIn1 = 32'd746
; 
32'd14628: dataIn1 = 32'd791
; 
32'd14629: dataIn1 = 32'd794
; 
32'd14630: dataIn1 = 32'd846
; 
32'd14631: dataIn1 = 32'd648
; 
32'd14632: dataIn1 = 32'd695
; 
32'd14633: dataIn1 = 32'd720
; 
32'd14634: dataIn1 = 32'd747
; 
32'd14635: dataIn1 = 32'd771
; 
32'd14636: dataIn1 = 32'd780
; 
32'd14637: dataIn1 = 32'd836
; 
32'd14638: dataIn1 = 32'd842
; 
32'd14639: dataIn1 = 32'd876
; 
32'd14640: dataIn1 = 32'd650
; 
32'd14641: dataIn1 = 32'd689
; 
32'd14642: dataIn1 = 32'd741
; 
32'd14643: dataIn1 = 32'd748
; 
32'd14644: dataIn1 = 32'd782
; 
32'd14645: dataIn1 = 32'd789
; 
32'd14646: dataIn1 = 32'd803
; 
32'd14647: dataIn1 = 32'd845
; 
32'd14648: dataIn1 = 32'd652
; 
32'd14649: dataIn1 = 32'd704
; 
32'd14650: dataIn1 = 32'd745
; 
32'd14651: dataIn1 = 32'd749
; 
32'd14652: dataIn1 = 32'd795
; 
32'd14653: dataIn1 = 32'd813
; 
32'd14654: dataIn1 = 32'd655
; 
32'd14655: dataIn1 = 32'd710
; 
32'd14656: dataIn1 = 32'd720
; 
32'd14657: dataIn1 = 32'd750
; 
32'd14658: dataIn1 = 32'd783
; 
32'd14659: dataIn1 = 32'd797
; 
32'd14660: dataIn1 = 32'd798
; 
32'd14661: dataIn1 = 32'd836
; 
32'd14662: dataIn1 = 32'd659
; 
32'd14663: dataIn1 = 32'd662
; 
32'd14664: dataIn1 = 32'd673
; 
32'd14665: dataIn1 = 32'd751
; 
32'd14666: dataIn1 = 32'd777
; 
32'd14667: dataIn1 = 32'd793
; 
32'd14668: dataIn1 = 32'd820
; 
32'd14669: dataIn1 = 32'd662
; 
32'd14670: dataIn1 = 32'd671
; 
32'd14671: dataIn1 = 32'd704
; 
32'd14672: dataIn1 = 32'd752
; 
32'd14673: dataIn1 = 32'd760
; 
32'd14674: dataIn1 = 32'd796
; 
32'd14675: dataIn1 = 32'd663
; 
32'd14676: dataIn1 = 32'd664
; 
32'd14677: dataIn1 = 32'd706
; 
32'd14678: dataIn1 = 32'd753
; 
32'd14679: dataIn1 = 32'd762
; 
32'd14680: dataIn1 = 32'd809
; 
32'd14681: dataIn1 = 32'd632
; 
32'd14682: dataIn1 = 32'd668
; 
32'd14683: dataIn1 = 32'd674
; 
32'd14684: dataIn1 = 32'd754
; 
32'd14685: dataIn1 = 32'd785
; 
32'd14686: dataIn1 = 32'd650
; 
32'd14687: dataIn1 = 32'd669
; 
32'd14688: dataIn1 = 32'd725
; 
32'd14689: dataIn1 = 32'd755
; 
32'd14690: dataIn1 = 32'd788
; 
32'd14691: dataIn1 = 32'd810
; 
32'd14692: dataIn1 = 32'd847
; 
32'd14693: dataIn1 = 32'd672
; 
32'd14694: dataIn1 = 32'd675
; 
32'd14695: dataIn1 = 32'd731
; 
32'd14696: dataIn1 = 32'd756
; 
32'd14697: dataIn1 = 32'd800
; 
32'd14698: dataIn1 = 32'd826
; 
32'd14699: dataIn1 = 32'd834
; 
32'd14700: dataIn1 = 32'd674
; 
32'd14701: dataIn1 = 32'd693
; 
32'd14702: dataIn1 = 32'd729
; 
32'd14703: dataIn1 = 32'd757
; 
32'd14704: dataIn1 = 32'd785
; 
32'd14705: dataIn1 = 32'd814
; 
32'd14706: dataIn1 = 32'd677
; 
32'd14707: dataIn1 = 32'd681
; 
32'd14708: dataIn1 = 32'd708
; 
32'd14709: dataIn1 = 32'd758
; 
32'd14710: dataIn1 = 32'd837
; 
32'd14711: dataIn1 = 32'd853
; 
32'd14712: dataIn1 = 32'd652
; 
32'd14713: dataIn1 = 32'd678
; 
32'd14714: dataIn1 = 32'd703
; 
32'd14715: dataIn1 = 32'd759
; 
32'd14716: dataIn1 = 32'd815
; 
32'd14717: dataIn1 = 32'd824
; 
32'd14718: dataIn1 = 32'd838
; 
32'd14719: dataIn1 = 32'd679
; 
32'd14720: dataIn1 = 32'd704
; 
32'd14721: dataIn1 = 32'd752
; 
32'd14722: dataIn1 = 32'd760
; 
32'd14723: dataIn1 = 32'd813
; 
32'd14724: dataIn1 = 32'd682
; 
32'd14725: dataIn1 = 32'd685
; 
32'd14726: dataIn1 = 32'd701
; 
32'd14727: dataIn1 = 32'd761
; 
32'd14728: dataIn1 = 32'd683
; 
32'd14729: dataIn1 = 32'd741
; 
32'd14730: dataIn1 = 32'd753
; 
32'd14731: dataIn1 = 32'd762
; 
32'd14732: dataIn1 = 32'd789
; 
32'd14733: dataIn1 = 32'd839
; 
32'd14734: dataIn1 = 32'd659
; 
32'd14735: dataIn1 = 32'd687
; 
32'd14736: dataIn1 = 32'd694
; 
32'd14737: dataIn1 = 32'd763
; 
32'd14738: dataIn1 = 32'd793
; 
32'd14739: dataIn1 = 32'd798
; 
32'd14740: dataIn1 = 32'd822
; 
32'd14741: dataIn1 = 32'd678
; 
32'd14742: dataIn1 = 32'd688
; 
32'd14743: dataIn1 = 32'd734
; 
32'd14744: dataIn1 = 32'd764
; 
32'd14745: dataIn1 = 32'd781
; 
32'd14746: dataIn1 = 32'd807
; 
32'd14747: dataIn1 = 32'd607
; 
32'd14748: dataIn1 = 32'd664
; 
32'd14749: dataIn1 = 32'd689
; 
32'd14750: dataIn1 = 32'd765
; 
32'd14751: dataIn1 = 32'd766
; 
32'd14752: dataIn1 = 32'd664
; 
32'd14753: dataIn1 = 32'd706
; 
32'd14754: dataIn1 = 32'd765
; 
32'd14755: dataIn1 = 32'd766
; 
32'd14756: dataIn1 = 32'd803
; 
32'd14757: dataIn1 = 32'd811
; 
32'd14758: dataIn1 = 32'd829
; 
32'd14759: dataIn1 = 32'd709
; 
32'd14760: dataIn1 = 32'd722
; 
32'd14761: dataIn1 = 32'd723
; 
32'd14762: dataIn1 = 32'd767
; 
32'd14763: dataIn1 = 32'd779
; 
32'd14764: dataIn1 = 32'd797
; 
32'd14765: dataIn1 = 32'd828
; 
32'd14766: dataIn1 = 32'd648
; 
32'd14767: dataIn1 = 32'd684
; 
32'd14768: dataIn1 = 32'd722
; 
32'd14769: dataIn1 = 32'd768
; 
32'd14770: dataIn1 = 32'd780
; 
32'd14771: dataIn1 = 32'd674
; 
32'd14772: dataIn1 = 32'd689
; 
32'd14773: dataIn1 = 32'd693
; 
32'd14774: dataIn1 = 32'd769
; 
32'd14775: dataIn1 = 32'd816
; 
32'd14776: dataIn1 = 32'd823
; 
32'd14777: dataIn1 = 32'd849
; 
32'd14778: dataIn1 = 32'd670
; 
32'd14779: dataIn1 = 32'd678
; 
32'd14780: dataIn1 = 32'd686
; 
32'd14781: dataIn1 = 32'd770
; 
32'd14782: dataIn1 = 32'd781
; 
32'd14783: dataIn1 = 32'd662
; 
32'd14784: dataIn1 = 32'd679
; 
32'd14785: dataIn1 = 32'd747
; 
32'd14786: dataIn1 = 32'd771
; 
32'd14787: dataIn1 = 32'd802
; 
32'd14788: dataIn1 = 32'd674
; 
32'd14789: dataIn1 = 32'd701
; 
32'd14790: dataIn1 = 32'd711
; 
32'd14791: dataIn1 = 32'd772
; 
32'd14792: dataIn1 = 32'd823
; 
32'd14793: dataIn1 = 32'd827
; 
32'd14794: dataIn1 = 32'd677
; 
32'd14795: dataIn1 = 32'd699
; 
32'd14796: dataIn1 = 32'd728
; 
32'd14797: dataIn1 = 32'd773
; 
32'd14798: dataIn1 = 32'd830
; 
32'd14799: dataIn1 = 32'd694
; 
32'd14800: dataIn1 = 32'd710
; 
32'd14801: dataIn1 = 32'd711
; 
32'd14802: dataIn1 = 32'd774
; 
32'd14803: dataIn1 = 32'd798
; 
32'd14804: dataIn1 = 32'd840
; 
32'd14805: dataIn1 = 32'd854
; 
32'd14806: dataIn1 = 32'd870
; 
32'd14807: dataIn1 = 32'd713
; 
32'd14808: dataIn1 = 32'd723
; 
32'd14809: dataIn1 = 32'd735
; 
32'd14810: dataIn1 = 32'd775
; 
32'd14811: dataIn1 = 32'd781
; 
32'd14812: dataIn1 = 32'd828
; 
32'd14813: dataIn1 = 32'd841
; 
32'd14814: dataIn1 = 32'd869
; 
32'd14815: dataIn1 = 32'd701
; 
32'd14816: dataIn1 = 32'd710
; 
32'd14817: dataIn1 = 32'd719
; 
32'd14818: dataIn1 = 32'd776
; 
32'd14819: dataIn1 = 32'd783
; 
32'd14820: dataIn1 = 32'd827
; 
32'd14821: dataIn1 = 32'd840
; 
32'd14822: dataIn1 = 32'd873
; 
32'd14823: dataIn1 = 32'd671
; 
32'd14824: dataIn1 = 32'd673
; 
32'd14825: dataIn1 = 32'd751
; 
32'd14826: dataIn1 = 32'd777
; 
32'd14827: dataIn1 = 32'd796
; 
32'd14828: dataIn1 = 32'd820
; 
32'd14829: dataIn1 = 32'd679
; 
32'd14830: dataIn1 = 32'd730
; 
32'd14831: dataIn1 = 32'd743
; 
32'd14832: dataIn1 = 32'd778
; 
32'd14833: dataIn1 = 32'd835
; 
32'd14834: dataIn1 = 32'd842
; 
32'd14835: dataIn1 = 32'd906
; 
32'd14836: dataIn1 = 32'd681
; 
32'd14837: dataIn1 = 32'd735
; 
32'd14838: dataIn1 = 32'd767
; 
32'd14839: dataIn1 = 32'd779
; 
32'd14840: dataIn1 = 32'd828
; 
32'd14841: dataIn1 = 32'd837
; 
32'd14842: dataIn1 = 32'd869
; 
32'd14843: dataIn1 = 32'd880
; 
32'd14844: dataIn1 = 32'd720
; 
32'd14845: dataIn1 = 32'd747
; 
32'd14846: dataIn1 = 32'd768
; 
32'd14847: dataIn1 = 32'd780
; 
32'd14848: dataIn1 = 32'd797
; 
32'd14849: dataIn1 = 32'd764
; 
32'd14850: dataIn1 = 32'd770
; 
32'd14851: dataIn1 = 32'd775
; 
32'd14852: dataIn1 = 32'd781
; 
32'd14853: dataIn1 = 32'd817
; 
32'd14854: dataIn1 = 32'd824
; 
32'd14855: dataIn1 = 32'd877
; 
32'd14856: dataIn1 = 32'd888
; 
32'd14857: dataIn1 = 32'd912
; 
32'd14858: dataIn1 = 32'd929
; 
32'd14859: dataIn1 = 32'd933
; 
32'd14860: dataIn1 = 32'd689
; 
32'd14861: dataIn1 = 32'd740
; 
32'd14862: dataIn1 = 32'd748
; 
32'd14863: dataIn1 = 32'd782
; 
32'd14864: dataIn1 = 32'd816
; 
32'd14865: dataIn1 = 32'd721
; 
32'd14866: dataIn1 = 32'd750
; 
32'd14867: dataIn1 = 32'd776
; 
32'd14868: dataIn1 = 32'd783
; 
32'd14869: dataIn1 = 32'd881
; 
32'd14870: dataIn1 = 32'd683
; 
32'd14871: dataIn1 = 32'd724
; 
32'd14872: dataIn1 = 32'd725
; 
32'd14873: dataIn1 = 32'd784
; 
32'd14874: dataIn1 = 32'd806
; 
32'd14875: dataIn1 = 32'd808
; 
32'd14876: dataIn1 = 32'd839
; 
32'd14877: dataIn1 = 32'd843
; 
32'd14878: dataIn1 = 32'd851
; 
32'd14879: dataIn1 = 32'd674
; 
32'd14880: dataIn1 = 32'd754
; 
32'd14881: dataIn1 = 32'd757
; 
32'd14882: dataIn1 = 32'd785
; 
32'd14883: dataIn1 = 32'd827
; 
32'd14884: dataIn1 = 32'd844
; 
32'd14885: dataIn1 = 32'd849
; 
32'd14886: dataIn1 = 32'd859
; 
32'd14887: dataIn1 = 32'd650
; 
32'd14888: dataIn1 = 32'd725
; 
32'd14889: dataIn1 = 32'd741
; 
32'd14890: dataIn1 = 32'd786
; 
32'd14891: dataIn1 = 32'd812
; 
32'd14892: dataIn1 = 32'd843
; 
32'd14893: dataIn1 = 32'd845
; 
32'd14894: dataIn1 = 32'd682
; 
32'd14895: dataIn1 = 32'd717
; 
32'd14896: dataIn1 = 32'd742
; 
32'd14897: dataIn1 = 32'd787
; 
32'd14898: dataIn1 = 32'd825
; 
32'd14899: dataIn1 = 32'd844
; 
32'd14900: dataIn1 = 32'd846
; 
32'd14901: dataIn1 = 32'd848
; 
32'd14902: dataIn1 = 32'd635
; 
32'd14903: dataIn1 = 32'd743
; 
32'd14904: dataIn1 = 32'd755
; 
32'd14905: dataIn1 = 32'd788
; 
32'd14906: dataIn1 = 32'd835
; 
32'd14907: dataIn1 = 32'd847
; 
32'd14908: dataIn1 = 32'd864
; 
32'd14909: dataIn1 = 32'd878
; 
32'd14910: dataIn1 = 32'd903
; 
32'd14911: dataIn1 = 32'd741
; 
32'd14912: dataIn1 = 32'd748
; 
32'd14913: dataIn1 = 32'd762
; 
32'd14914: dataIn1 = 32'd789
; 
32'd14915: dataIn1 = 32'd697
; 
32'd14916: dataIn1 = 32'd706
; 
32'd14917: dataIn1 = 32'd726
; 
32'd14918: dataIn1 = 32'd790
; 
32'd14919: dataIn1 = 32'd805
; 
32'd14920: dataIn1 = 32'd811
; 
32'd14921: dataIn1 = 32'd829
; 
32'd14922: dataIn1 = 32'd850
; 
32'd14923: dataIn1 = 32'd863
; 
32'd14924: dataIn1 = 32'd868
; 
32'd14925: dataIn1 = 32'd715
; 
32'd14926: dataIn1 = 32'd732
; 
32'd14927: dataIn1 = 32'd746
; 
32'd14928: dataIn1 = 32'd791
; 
32'd14929: dataIn1 = 32'd792
; 
32'd14930: dataIn1 = 32'd806
; 
32'd14931: dataIn1 = 32'd825
; 
32'd14932: dataIn1 = 32'd857
; 
32'd14933: dataIn1 = 32'd731
; 
32'd14934: dataIn1 = 32'd732
; 
32'd14935: dataIn1 = 32'd791
; 
32'd14936: dataIn1 = 32'd792
; 
32'd14937: dataIn1 = 32'd834
; 
32'd14938: dataIn1 = 32'd865
; 
32'd14939: dataIn1 = 32'd659
; 
32'd14940: dataIn1 = 32'd751
; 
32'd14941: dataIn1 = 32'd763
; 
32'd14942: dataIn1 = 32'd793
; 
32'd14943: dataIn1 = 32'd692
; 
32'd14944: dataIn1 = 32'd705
; 
32'd14945: dataIn1 = 32'd746
; 
32'd14946: dataIn1 = 32'd794
; 
32'd14947: dataIn1 = 32'd819
; 
32'd14948: dataIn1 = 32'd857
; 
32'd14949: dataIn1 = 32'd871
; 
32'd14950: dataIn1 = 32'd727
; 
32'd14951: dataIn1 = 32'd745
; 
32'd14952: dataIn1 = 32'd749
; 
32'd14953: dataIn1 = 32'd795
; 
32'd14954: dataIn1 = 32'd818
; 
32'd14955: dataIn1 = 32'd838
; 
32'd14956: dataIn1 = 32'd861
; 
32'd14957: dataIn1 = 32'd662
; 
32'd14958: dataIn1 = 32'd752
; 
32'd14959: dataIn1 = 32'd777
; 
32'd14960: dataIn1 = 32'd796
; 
32'd14961: dataIn1 = 32'd802
; 
32'd14962: dataIn1 = 32'd820
; 
32'd14963: dataIn1 = 32'd821
; 
32'd14964: dataIn1 = 32'd868
; 
32'd14965: dataIn1 = 32'd895
; 
32'd14966: dataIn1 = 32'd901
; 
32'd14967: dataIn1 = 32'd750
; 
32'd14968: dataIn1 = 32'd767
; 
32'd14969: dataIn1 = 32'd780
; 
32'd14970: dataIn1 = 32'd797
; 
32'd14971: dataIn1 = 32'd880
; 
32'd14972: dataIn1 = 32'd881
; 
32'd14973: dataIn1 = 32'd750
; 
32'd14974: dataIn1 = 32'd763
; 
32'd14975: dataIn1 = 32'd774
; 
32'd14976: dataIn1 = 32'd798
; 
32'd14977: dataIn1 = 32'd836
; 
32'd14978: dataIn1 = 32'd840
; 
32'd14979: dataIn1 = 32'd677
; 
32'd14980: dataIn1 = 32'd729
; 
32'd14981: dataIn1 = 32'd744
; 
32'd14982: dataIn1 = 32'd799
; 
32'd14983: dataIn1 = 32'd814
; 
32'd14984: dataIn1 = 32'd852
; 
32'd14985: dataIn1 = 32'd875
; 
32'd14986: dataIn1 = 32'd882
; 
32'd14987: dataIn1 = 32'd681
; 
32'd14988: dataIn1 = 32'd744
; 
32'd14989: dataIn1 = 32'd756
; 
32'd14990: dataIn1 = 32'd800
; 
32'd14991: dataIn1 = 32'd837
; 
32'd14992: dataIn1 = 32'd875
; 
32'd14993: dataIn1 = 32'd883
; 
32'd14994: dataIn1 = 32'd886
; 
32'd14995: dataIn1 = 32'd682
; 
32'd14996: dataIn1 = 32'd692
; 
32'd14997: dataIn1 = 32'd734
; 
32'd14998: dataIn1 = 32'd801
; 
32'd14999: dataIn1 = 32'd817
; 
32'd15000: dataIn1 = 32'd848
; 
32'd15001: dataIn1 = 32'd871
; 
32'd15002: dataIn1 = 32'd877
; 
32'd15003: dataIn1 = 32'd687
; 
32'd15004: dataIn1 = 32'd771
; 
32'd15005: dataIn1 = 32'd796
; 
32'd15006: dataIn1 = 32'd802
; 
32'd15007: dataIn1 = 32'd821
; 
32'd15008: dataIn1 = 32'd842
; 
32'd15009: dataIn1 = 32'd884
; 
32'd15010: dataIn1 = 32'd689
; 
32'd15011: dataIn1 = 32'd748
; 
32'd15012: dataIn1 = 32'd766
; 
32'd15013: dataIn1 = 32'd803
; 
32'd15014: dataIn1 = 32'd816
; 
32'd15015: dataIn1 = 32'd831
; 
32'd15016: dataIn1 = 32'd677
; 
32'd15017: dataIn1 = 32'd693
; 
32'd15018: dataIn1 = 32'd740
; 
32'd15019: dataIn1 = 32'd804
; 
32'd15020: dataIn1 = 32'd833
; 
32'd15021: dataIn1 = 32'd849
; 
32'd15022: dataIn1 = 32'd882
; 
32'd15023: dataIn1 = 32'd885
; 
32'd15024: dataIn1 = 32'd887
; 
32'd15025: dataIn1 = 32'd697
; 
32'd15026: dataIn1 = 32'd726
; 
32'd15027: dataIn1 = 32'd790
; 
32'd15028: dataIn1 = 32'd805
; 
32'd15029: dataIn1 = 32'd819
; 
32'd15030: dataIn1 = 32'd850
; 
32'd15031: dataIn1 = 32'd715
; 
32'd15032: dataIn1 = 32'd784
; 
32'd15033: dataIn1 = 32'd791
; 
32'd15034: dataIn1 = 32'd806
; 
32'd15035: dataIn1 = 32'd721
; 
32'd15036: dataIn1 = 32'd733
; 
32'd15037: dataIn1 = 32'd764
; 
32'd15038: dataIn1 = 32'd807
; 
32'd15039: dataIn1 = 32'd841
; 
32'd15040: dataIn1 = 32'd725
; 
32'd15041: dataIn1 = 32'd731
; 
32'd15042: dataIn1 = 32'd784
; 
32'd15043: dataIn1 = 32'd808
; 
32'd15044: dataIn1 = 32'd832
; 
32'd15045: dataIn1 = 32'd851
; 
32'd15046: dataIn1 = 32'd862
; 
32'd15047: dataIn1 = 32'd726
; 
32'd15048: dataIn1 = 32'd738
; 
32'd15049: dataIn1 = 32'd753
; 
32'd15050: dataIn1 = 32'd809
; 
32'd15051: dataIn1 = 32'd819
; 
32'd15052: dataIn1 = 32'd839
; 
32'd15053: dataIn1 = 32'd730
; 
32'd15054: dataIn1 = 32'd740
; 
32'd15055: dataIn1 = 32'd755
; 
32'd15056: dataIn1 = 32'd810
; 
32'd15057: dataIn1 = 32'd812
; 
32'd15058: dataIn1 = 32'd833
; 
32'd15059: dataIn1 = 32'd736
; 
32'd15060: dataIn1 = 32'd766
; 
32'd15061: dataIn1 = 32'd790
; 
32'd15062: dataIn1 = 32'd811
; 
32'd15063: dataIn1 = 32'd822
; 
32'd15064: dataIn1 = 32'd829
; 
32'd15065: dataIn1 = 32'd740
; 
32'd15066: dataIn1 = 32'd786
; 
32'd15067: dataIn1 = 32'd810
; 
32'd15068: dataIn1 = 32'd812
; 
32'd15069: dataIn1 = 32'd845
; 
32'd15070: dataIn1 = 32'd743
; 
32'd15071: dataIn1 = 32'd749
; 
32'd15072: dataIn1 = 32'd760
; 
32'd15073: dataIn1 = 32'd813
; 
32'd15074: dataIn1 = 32'd855
; 
32'd15075: dataIn1 = 32'd866
; 
32'd15076: dataIn1 = 32'd742
; 
32'd15077: dataIn1 = 32'd757
; 
32'd15078: dataIn1 = 32'd799
; 
32'd15079: dataIn1 = 32'd814
; 
32'd15080: dataIn1 = 32'd852
; 
32'd15081: dataIn1 = 32'd678
; 
32'd15082: dataIn1 = 32'd745
; 
32'd15083: dataIn1 = 32'd759
; 
32'd15084: dataIn1 = 32'd815
; 
32'd15085: dataIn1 = 32'd838
; 
32'd15086: dataIn1 = 32'd769
; 
32'd15087: dataIn1 = 32'd782
; 
32'd15088: dataIn1 = 32'd803
; 
32'd15089: dataIn1 = 32'd816
; 
32'd15090: dataIn1 = 32'd872
; 
32'd15091: dataIn1 = 32'd885
; 
32'd15092: dataIn1 = 32'd733
; 
32'd15093: dataIn1 = 32'd781
; 
32'd15094: dataIn1 = 32'd801
; 
32'd15095: dataIn1 = 32'd817
; 
32'd15096: dataIn1 = 32'd873
; 
32'd15097: dataIn1 = 32'd889
; 
32'd15098: dataIn1 = 32'd913
; 
32'd15099: dataIn1 = 32'd929
; 
32'd15100: dataIn1 = 32'd935
; 
32'd15101: dataIn1 = 32'd718
; 
32'd15102: dataIn1 = 32'd727
; 
32'd15103: dataIn1 = 32'd795
; 
32'd15104: dataIn1 = 32'd818
; 
32'd15105: dataIn1 = 32'd861
; 
32'd15106: dataIn1 = 32'd910
; 
32'd15107: dataIn1 = 32'd911
; 
32'd15108: dataIn1 = 32'd912
; 
32'd15109: dataIn1 = 32'd794
; 
32'd15110: dataIn1 = 32'd805
; 
32'd15111: dataIn1 = 32'd809
; 
32'd15112: dataIn1 = 32'd819
; 
32'd15113: dataIn1 = 32'd863
; 
32'd15114: dataIn1 = 32'd751
; 
32'd15115: dataIn1 = 32'd777
; 
32'd15116: dataIn1 = 32'd796
; 
32'd15117: dataIn1 = 32'd820
; 
32'd15118: dataIn1 = 32'd821
; 
32'd15119: dataIn1 = 32'd796
; 
32'd15120: dataIn1 = 32'd802
; 
32'd15121: dataIn1 = 32'd820
; 
32'd15122: dataIn1 = 32'd821
; 
32'd15123: dataIn1 = 32'd895
; 
32'd15124: dataIn1 = 32'd900
; 
32'd15125: dataIn1 = 32'd914
; 
32'd15126: dataIn1 = 32'd930
; 
32'd15127: dataIn1 = 32'd737
; 
32'd15128: dataIn1 = 32'd763
; 
32'd15129: dataIn1 = 32'd811
; 
32'd15130: dataIn1 = 32'd822
; 
32'd15131: dataIn1 = 32'd874
; 
32'd15132: dataIn1 = 32'd914
; 
32'd15133: dataIn1 = 32'd931
; 
32'd15134: dataIn1 = 32'd737
; 
32'd15135: dataIn1 = 32'd769
; 
32'd15136: dataIn1 = 32'd772
; 
32'd15137: dataIn1 = 32'd823
; 
32'd15138: dataIn1 = 32'd854
; 
32'd15139: dataIn1 = 32'd915
; 
32'd15140: dataIn1 = 32'd920
; 
32'd15141: dataIn1 = 32'd735
; 
32'd15142: dataIn1 = 32'd759
; 
32'd15143: dataIn1 = 32'd781
; 
32'd15144: dataIn1 = 32'd824
; 
32'd15145: dataIn1 = 32'd860
; 
32'd15146: dataIn1 = 32'd742
; 
32'd15147: dataIn1 = 32'd787
; 
32'd15148: dataIn1 = 32'd791
; 
32'd15149: dataIn1 = 32'd825
; 
32'd15150: dataIn1 = 32'd846
; 
32'd15151: dataIn1 = 32'd857
; 
32'd15152: dataIn1 = 32'd867
; 
32'd15153: dataIn1 = 32'd907
; 
32'd15154: dataIn1 = 32'd916
; 
32'd15155: dataIn1 = 32'd672
; 
32'd15156: dataIn1 = 32'd731
; 
32'd15157: dataIn1 = 32'd756
; 
32'd15158: dataIn1 = 32'd826
; 
32'd15159: dataIn1 = 32'd883
; 
32'd15160: dataIn1 = 32'd891
; 
32'd15161: dataIn1 = 32'd772
; 
32'd15162: dataIn1 = 32'd776
; 
32'd15163: dataIn1 = 32'd785
; 
32'd15164: dataIn1 = 32'd827
; 
32'd15165: dataIn1 = 32'd870
; 
32'd15166: dataIn1 = 32'd873
; 
32'd15167: dataIn1 = 32'd896
; 
32'd15168: dataIn1 = 32'd915
; 
32'd15169: dataIn1 = 32'd918
; 
32'd15170: dataIn1 = 32'd767
; 
32'd15171: dataIn1 = 32'd775
; 
32'd15172: dataIn1 = 32'd779
; 
32'd15173: dataIn1 = 32'd828
; 
32'd15174: dataIn1 = 32'd841
; 
32'd15175: dataIn1 = 32'd766
; 
32'd15176: dataIn1 = 32'd790
; 
32'd15177: dataIn1 = 32'd811
; 
32'd15178: dataIn1 = 32'd829
; 
32'd15179: dataIn1 = 32'd831
; 
32'd15180: dataIn1 = 32'd728
; 
32'd15181: dataIn1 = 32'd730
; 
32'd15182: dataIn1 = 32'd773
; 
32'd15183: dataIn1 = 32'd830
; 
32'd15184: dataIn1 = 32'd853
; 
32'd15185: dataIn1 = 32'd882
; 
32'd15186: dataIn1 = 32'd887
; 
32'd15187: dataIn1 = 32'd890
; 
32'd15188: dataIn1 = 32'd906
; 
32'd15189: dataIn1 = 32'd945
; 
32'd15190: dataIn1 = 32'd737
; 
32'd15191: dataIn1 = 32'd803
; 
32'd15192: dataIn1 = 32'd829
; 
32'd15193: dataIn1 = 32'd831
; 
32'd15194: dataIn1 = 32'd872
; 
32'd15195: dataIn1 = 32'd893
; 
32'd15196: dataIn1 = 32'd897
; 
32'd15197: dataIn1 = 32'd920
; 
32'd15198: dataIn1 = 32'd926
; 
32'd15199: dataIn1 = 32'd931
; 
32'd15200: dataIn1 = 32'd635
; 
32'd15201: dataIn1 = 32'd739
; 
32'd15202: dataIn1 = 32'd808
; 
32'd15203: dataIn1 = 32'd832
; 
32'd15204: dataIn1 = 32'd855
; 
32'd15205: dataIn1 = 32'd858
; 
32'd15206: dataIn1 = 32'd862
; 
32'd15207: dataIn1 = 32'd908
; 
32'd15208: dataIn1 = 32'd740
; 
32'd15209: dataIn1 = 32'd804
; 
32'd15210: dataIn1 = 32'd810
; 
32'd15211: dataIn1 = 32'd833
; 
32'd15212: dataIn1 = 32'd887
; 
32'd15213: dataIn1 = 32'd742
; 
32'd15214: dataIn1 = 32'd756
; 
32'd15215: dataIn1 = 32'd792
; 
32'd15216: dataIn1 = 32'd834
; 
32'd15217: dataIn1 = 32'd886
; 
32'd15218: dataIn1 = 32'd891
; 
32'd15219: dataIn1 = 32'd907
; 
32'd15220: dataIn1 = 32'd921
; 
32'd15221: dataIn1 = 32'd927
; 
32'd15222: dataIn1 = 32'd743
; 
32'd15223: dataIn1 = 32'd778
; 
32'd15224: dataIn1 = 32'd788
; 
32'd15225: dataIn1 = 32'd835
; 
32'd15226: dataIn1 = 32'd864
; 
32'd15227: dataIn1 = 32'd866
; 
32'd15228: dataIn1 = 32'd903
; 
32'd15229: dataIn1 = 32'd747
; 
32'd15230: dataIn1 = 32'd750
; 
32'd15231: dataIn1 = 32'd798
; 
32'd15232: dataIn1 = 32'd836
; 
32'd15233: dataIn1 = 32'd876
; 
32'd15234: dataIn1 = 32'd881
; 
32'd15235: dataIn1 = 32'd884
; 
32'd15236: dataIn1 = 32'd892
; 
32'd15237: dataIn1 = 32'd900
; 
32'd15238: dataIn1 = 32'd902
; 
32'd15239: dataIn1 = 32'd758
; 
32'd15240: dataIn1 = 32'd779
; 
32'd15241: dataIn1 = 32'd800
; 
32'd15242: dataIn1 = 32'd837
; 
32'd15243: dataIn1 = 32'd875
; 
32'd15244: dataIn1 = 32'd894
; 
32'd15245: dataIn1 = 32'd909
; 
32'd15246: dataIn1 = 32'd759
; 
32'd15247: dataIn1 = 32'd795
; 
32'd15248: dataIn1 = 32'd815
; 
32'd15249: dataIn1 = 32'd838
; 
32'd15250: dataIn1 = 32'd856
; 
32'd15251: dataIn1 = 32'd860
; 
32'd15252: dataIn1 = 32'd879
; 
32'd15253: dataIn1 = 32'd762
; 
32'd15254: dataIn1 = 32'd784
; 
32'd15255: dataIn1 = 32'd809
; 
32'd15256: dataIn1 = 32'd839
; 
32'd15257: dataIn1 = 32'd897
; 
32'd15258: dataIn1 = 32'd774
; 
32'd15259: dataIn1 = 32'd776
; 
32'd15260: dataIn1 = 32'd798
; 
32'd15261: dataIn1 = 32'd840
; 
32'd15262: dataIn1 = 32'd870
; 
32'd15263: dataIn1 = 32'd874
; 
32'd15264: dataIn1 = 32'd904
; 
32'd15265: dataIn1 = 32'd775
; 
32'd15266: dataIn1 = 32'd807
; 
32'd15267: dataIn1 = 32'd828
; 
32'd15268: dataIn1 = 32'd841
; 
32'd15269: dataIn1 = 32'd889
; 
32'd15270: dataIn1 = 32'd747
; 
32'd15271: dataIn1 = 32'd778
; 
32'd15272: dataIn1 = 32'd802
; 
32'd15273: dataIn1 = 32'd842
; 
32'd15274: dataIn1 = 32'd876
; 
32'd15275: dataIn1 = 32'd884
; 
32'd15276: dataIn1 = 32'd895
; 
32'd15277: dataIn1 = 32'd902
; 
32'd15278: dataIn1 = 32'd930
; 
32'd15279: dataIn1 = 32'd725
; 
32'd15280: dataIn1 = 32'd784
; 
32'd15281: dataIn1 = 32'd786
; 
32'd15282: dataIn1 = 32'd843
; 
32'd15283: dataIn1 = 32'd878
; 
32'd15284: dataIn1 = 32'd897
; 
32'd15285: dataIn1 = 32'd742
; 
32'd15286: dataIn1 = 32'd785
; 
32'd15287: dataIn1 = 32'd787
; 
32'd15288: dataIn1 = 32'd844
; 
32'd15289: dataIn1 = 32'd867
; 
32'd15290: dataIn1 = 32'd748
; 
32'd15291: dataIn1 = 32'd786
; 
32'd15292: dataIn1 = 32'd812
; 
32'd15293: dataIn1 = 32'd845
; 
32'd15294: dataIn1 = 32'd872
; 
32'd15295: dataIn1 = 32'd746
; 
32'd15296: dataIn1 = 32'd787
; 
32'd15297: dataIn1 = 32'd825
; 
32'd15298: dataIn1 = 32'd846
; 
32'd15299: dataIn1 = 32'd730
; 
32'd15300: dataIn1 = 32'd755
; 
32'd15301: dataIn1 = 32'd788
; 
32'd15302: dataIn1 = 32'd847
; 
32'd15303: dataIn1 = 32'd864
; 
32'd15304: dataIn1 = 32'd878
; 
32'd15305: dataIn1 = 32'd682
; 
32'd15306: dataIn1 = 32'd787
; 
32'd15307: dataIn1 = 32'd801
; 
32'd15308: dataIn1 = 32'd848
; 
32'd15309: dataIn1 = 32'd896
; 
32'd15310: dataIn1 = 32'd913
; 
32'd15311: dataIn1 = 32'd769
; 
32'd15312: dataIn1 = 32'd785
; 
32'd15313: dataIn1 = 32'd804
; 
32'd15314: dataIn1 = 32'd849
; 
32'd15315: dataIn1 = 32'd859
; 
32'd15316: dataIn1 = 32'd885
; 
32'd15317: dataIn1 = 32'd727
; 
32'd15318: dataIn1 = 32'd790
; 
32'd15319: dataIn1 = 32'd805
; 
32'd15320: dataIn1 = 32'd850
; 
32'd15321: dataIn1 = 32'd863
; 
32'd15322: dataIn1 = 32'd731
; 
32'd15323: dataIn1 = 32'd784
; 
32'd15324: dataIn1 = 32'd808
; 
32'd15325: dataIn1 = 32'd851
; 
32'd15326: dataIn1 = 32'd858
; 
32'd15327: dataIn1 = 32'd862
; 
32'd15328: dataIn1 = 32'd865
; 
32'd15329: dataIn1 = 32'd899
; 
32'd15330: dataIn1 = 32'd742
; 
32'd15331: dataIn1 = 32'd799
; 
32'd15332: dataIn1 = 32'd814
; 
32'd15333: dataIn1 = 32'd852
; 
32'd15334: dataIn1 = 32'd859
; 
32'd15335: dataIn1 = 32'd921
; 
32'd15336: dataIn1 = 32'd923
; 
32'd15337: dataIn1 = 32'd728
; 
32'd15338: dataIn1 = 32'd758
; 
32'd15339: dataIn1 = 32'd830
; 
32'd15340: dataIn1 = 32'd853
; 
32'd15341: dataIn1 = 32'd737
; 
32'd15342: dataIn1 = 32'd774
; 
32'd15343: dataIn1 = 32'd823
; 
32'd15344: dataIn1 = 32'd854
; 
32'd15345: dataIn1 = 32'd874
; 
32'd15346: dataIn1 = 32'd739
; 
32'd15347: dataIn1 = 32'd813
; 
32'd15348: dataIn1 = 32'd832
; 
32'd15349: dataIn1 = 32'd855
; 
32'd15350: dataIn1 = 32'd856
; 
32'd15351: dataIn1 = 32'd866
; 
32'd15352: dataIn1 = 32'd879
; 
32'd15353: dataIn1 = 32'd908
; 
32'd15354: dataIn1 = 32'd974
; 
32'd15355: dataIn1 = 32'd739
; 
32'd15356: dataIn1 = 32'd838
; 
32'd15357: dataIn1 = 32'd855
; 
32'd15358: dataIn1 = 32'd856
; 
32'd15359: dataIn1 = 32'd860
; 
32'd15360: dataIn1 = 32'd791
; 
32'd15361: dataIn1 = 32'd794
; 
32'd15362: dataIn1 = 32'd825
; 
32'd15363: dataIn1 = 32'd857
; 
32'd15364: dataIn1 = 32'd865
; 
32'd15365: dataIn1 = 32'd907
; 
32'd15366: dataIn1 = 32'd916
; 
32'd15367: dataIn1 = 32'd731
; 
32'd15368: dataIn1 = 32'd832
; 
32'd15369: dataIn1 = 32'd851
; 
32'd15370: dataIn1 = 32'd858
; 
32'd15371: dataIn1 = 32'd899
; 
32'd15372: dataIn1 = 32'd785
; 
32'd15373: dataIn1 = 32'd849
; 
32'd15374: dataIn1 = 32'd852
; 
32'd15375: dataIn1 = 32'd859
; 
32'd15376: dataIn1 = 32'd915
; 
32'd15377: dataIn1 = 32'd923
; 
32'd15378: dataIn1 = 32'd932
; 
32'd15379: dataIn1 = 32'd824
; 
32'd15380: dataIn1 = 32'd838
; 
32'd15381: dataIn1 = 32'd856
; 
32'd15382: dataIn1 = 32'd860
; 
32'd15383: dataIn1 = 32'd879
; 
32'd15384: dataIn1 = 32'd888
; 
32'd15385: dataIn1 = 32'd898
; 
32'd15386: dataIn1 = 32'd727
; 
32'd15387: dataIn1 = 32'd795
; 
32'd15388: dataIn1 = 32'd818
; 
32'd15389: dataIn1 = 32'd861
; 
32'd15390: dataIn1 = 32'd868
; 
32'd15391: dataIn1 = 32'd910
; 
32'd15392: dataIn1 = 32'd911
; 
32'd15393: dataIn1 = 32'd924
; 
32'd15394: dataIn1 = 32'd808
; 
32'd15395: dataIn1 = 32'd832
; 
32'd15396: dataIn1 = 32'd851
; 
32'd15397: dataIn1 = 32'd862
; 
32'd15398: dataIn1 = 32'd899
; 
32'd15399: dataIn1 = 32'd908
; 
32'd15400: dataIn1 = 32'd925
; 
32'd15401: dataIn1 = 32'd790
; 
32'd15402: dataIn1 = 32'd819
; 
32'd15403: dataIn1 = 32'd850
; 
32'd15404: dataIn1 = 32'd863
; 
32'd15405: dataIn1 = 32'd926
; 
32'd15406: dataIn1 = 32'd788
; 
32'd15407: dataIn1 = 32'd835
; 
32'd15408: dataIn1 = 32'd847
; 
32'd15409: dataIn1 = 32'd864
; 
32'd15410: dataIn1 = 32'd890
; 
32'd15411: dataIn1 = 32'd903
; 
32'd15412: dataIn1 = 32'd906
; 
32'd15413: dataIn1 = 32'd792
; 
32'd15414: dataIn1 = 32'd851
; 
32'd15415: dataIn1 = 32'd857
; 
32'd15416: dataIn1 = 32'd865
; 
32'd15417: dataIn1 = 32'd925
; 
32'd15418: dataIn1 = 32'd927
; 
32'd15419: dataIn1 = 32'd813
; 
32'd15420: dataIn1 = 32'd835
; 
32'd15421: dataIn1 = 32'd855
; 
32'd15422: dataIn1 = 32'd866
; 
32'd15423: dataIn1 = 32'd901
; 
32'd15424: dataIn1 = 32'd928
; 
32'd15425: dataIn1 = 32'd974
; 
32'd15426: dataIn1 = 32'd742
; 
32'd15427: dataIn1 = 32'd825
; 
32'd15428: dataIn1 = 32'd844
; 
32'd15429: dataIn1 = 32'd867
; 
32'd15430: dataIn1 = 32'd896
; 
32'd15431: dataIn1 = 32'd921
; 
32'd15432: dataIn1 = 32'd790
; 
32'd15433: dataIn1 = 32'd796
; 
32'd15434: dataIn1 = 32'd861
; 
32'd15435: dataIn1 = 32'd868
; 
32'd15436: dataIn1 = 32'd910
; 
32'd15437: dataIn1 = 32'd914
; 
32'd15438: dataIn1 = 32'd924
; 
32'd15439: dataIn1 = 32'd735
; 
32'd15440: dataIn1 = 32'd775
; 
32'd15441: dataIn1 = 32'd779
; 
32'd15442: dataIn1 = 32'd869
; 
32'd15443: dataIn1 = 32'd880
; 
32'd15444: dataIn1 = 32'd888
; 
32'd15445: dataIn1 = 32'd898
; 
32'd15446: dataIn1 = 32'd774
; 
32'd15447: dataIn1 = 32'd827
; 
32'd15448: dataIn1 = 32'd840
; 
32'd15449: dataIn1 = 32'd870
; 
32'd15450: dataIn1 = 32'd718
; 
32'd15451: dataIn1 = 32'd794
; 
32'd15452: dataIn1 = 32'd801
; 
32'd15453: dataIn1 = 32'd871
; 
32'd15454: dataIn1 = 32'd877
; 
32'd15455: dataIn1 = 32'd912
; 
32'd15456: dataIn1 = 32'd816
; 
32'd15457: dataIn1 = 32'd831
; 
32'd15458: dataIn1 = 32'd845
; 
32'd15459: dataIn1 = 32'd872
; 
32'd15460: dataIn1 = 32'd893
; 
32'd15461: dataIn1 = 32'd905
; 
32'd15462: dataIn1 = 32'd776
; 
32'd15463: dataIn1 = 32'd817
; 
32'd15464: dataIn1 = 32'd827
; 
32'd15465: dataIn1 = 32'd873
; 
32'd15466: dataIn1 = 32'd904
; 
32'd15467: dataIn1 = 32'd918
; 
32'd15468: dataIn1 = 32'd822
; 
32'd15469: dataIn1 = 32'd840
; 
32'd15470: dataIn1 = 32'd854
; 
32'd15471: dataIn1 = 32'd874
; 
32'd15472: dataIn1 = 32'd900
; 
32'd15473: dataIn1 = 32'd931
; 
32'd15474: dataIn1 = 32'd799
; 
32'd15475: dataIn1 = 32'd800
; 
32'd15476: dataIn1 = 32'd837
; 
32'd15477: dataIn1 = 32'd875
; 
32'd15478: dataIn1 = 32'd886
; 
32'd15479: dataIn1 = 32'd894
; 
32'd15480: dataIn1 = 32'd747
; 
32'd15481: dataIn1 = 32'd836
; 
32'd15482: dataIn1 = 32'd842
; 
32'd15483: dataIn1 = 32'd876
; 
32'd15484: dataIn1 = 32'd902
; 
32'd15485: dataIn1 = 32'd945
; 
32'd15486: dataIn1 = 32'd781
; 
32'd15487: dataIn1 = 32'd801
; 
32'd15488: dataIn1 = 32'd871
; 
32'd15489: dataIn1 = 32'd877
; 
32'd15490: dataIn1 = 32'd913
; 
32'd15491: dataIn1 = 32'd929
; 
32'd15492: dataIn1 = 32'd788
; 
32'd15493: dataIn1 = 32'd843
; 
32'd15494: dataIn1 = 32'd847
; 
32'd15495: dataIn1 = 32'd878
; 
32'd15496: dataIn1 = 32'd890
; 
32'd15497: dataIn1 = 32'd838
; 
32'd15498: dataIn1 = 32'd855
; 
32'd15499: dataIn1 = 32'd860
; 
32'd15500: dataIn1 = 32'd879
; 
32'd15501: dataIn1 = 32'd911
; 
32'd15502: dataIn1 = 32'd928
; 
32'd15503: dataIn1 = 32'd974
; 
32'd15504: dataIn1 = 32'd779
; 
32'd15505: dataIn1 = 32'd797
; 
32'd15506: dataIn1 = 32'd869
; 
32'd15507: dataIn1 = 32'd880
; 
32'd15508: dataIn1 = 32'd892
; 
32'd15509: dataIn1 = 32'd783
; 
32'd15510: dataIn1 = 32'd797
; 
32'd15511: dataIn1 = 32'd836
; 
32'd15512: dataIn1 = 32'd881
; 
32'd15513: dataIn1 = 32'd889
; 
32'd15514: dataIn1 = 32'd892
; 
32'd15515: dataIn1 = 32'd904
; 
32'd15516: dataIn1 = 32'd799
; 
32'd15517: dataIn1 = 32'd804
; 
32'd15518: dataIn1 = 32'd830
; 
32'd15519: dataIn1 = 32'd882
; 
32'd15520: dataIn1 = 32'd923
; 
32'd15521: dataIn1 = 32'd932
; 
32'd15522: dataIn1 = 32'd735
; 
32'd15523: dataIn1 = 32'd800
; 
32'd15524: dataIn1 = 32'd826
; 
32'd15525: dataIn1 = 32'd883
; 
32'd15526: dataIn1 = 32'd891
; 
32'd15527: dataIn1 = 32'd909
; 
32'd15528: dataIn1 = 32'd802
; 
32'd15529: dataIn1 = 32'd836
; 
32'd15530: dataIn1 = 32'd842
; 
32'd15531: dataIn1 = 32'd884
; 
32'd15532: dataIn1 = 32'd804
; 
32'd15533: dataIn1 = 32'd816
; 
32'd15534: dataIn1 = 32'd849
; 
32'd15535: dataIn1 = 32'd885
; 
32'd15536: dataIn1 = 32'd893
; 
32'd15537: dataIn1 = 32'd905
; 
32'd15538: dataIn1 = 32'd800
; 
32'd15539: dataIn1 = 32'd834
; 
32'd15540: dataIn1 = 32'd875
; 
32'd15541: dataIn1 = 32'd886
; 
32'd15542: dataIn1 = 32'd894
; 
32'd15543: dataIn1 = 32'd940
; 
32'd15544: dataIn1 = 32'd804
; 
32'd15545: dataIn1 = 32'd830
; 
32'd15546: dataIn1 = 32'd833
; 
32'd15547: dataIn1 = 32'd887
; 
32'd15548: dataIn1 = 32'd905
; 
32'd15549: dataIn1 = 32'd781
; 
32'd15550: dataIn1 = 32'd860
; 
32'd15551: dataIn1 = 32'd869
; 
32'd15552: dataIn1 = 32'd888
; 
32'd15553: dataIn1 = 32'd898
; 
32'd15554: dataIn1 = 32'd962
; 
32'd15555: dataIn1 = 32'd817
; 
32'd15556: dataIn1 = 32'd841
; 
32'd15557: dataIn1 = 32'd881
; 
32'd15558: dataIn1 = 32'd889
; 
32'd15559: dataIn1 = 32'd830
; 
32'd15560: dataIn1 = 32'd864
; 
32'd15561: dataIn1 = 32'd878
; 
32'd15562: dataIn1 = 32'd890
; 
32'd15563: dataIn1 = 32'd826
; 
32'd15564: dataIn1 = 32'd834
; 
32'd15565: dataIn1 = 32'd883
; 
32'd15566: dataIn1 = 32'd891
; 
32'd15567: dataIn1 = 32'd940
; 
32'd15568: dataIn1 = 32'd836
; 
32'd15569: dataIn1 = 32'd880
; 
32'd15570: dataIn1 = 32'd881
; 
32'd15571: dataIn1 = 32'd892
; 
32'd15572: dataIn1 = 32'd831
; 
32'd15573: dataIn1 = 32'd872
; 
32'd15574: dataIn1 = 32'd885
; 
32'd15575: dataIn1 = 32'd893
; 
32'd15576: dataIn1 = 32'd920
; 
32'd15577: dataIn1 = 32'd837
; 
32'd15578: dataIn1 = 32'd875
; 
32'd15579: dataIn1 = 32'd886
; 
32'd15580: dataIn1 = 32'd894
; 
32'd15581: dataIn1 = 32'd909
; 
32'd15582: dataIn1 = 32'd940
; 
32'd15583: dataIn1 = 32'd796
; 
32'd15584: dataIn1 = 32'd821
; 
32'd15585: dataIn1 = 32'd842
; 
32'd15586: dataIn1 = 32'd895
; 
32'd15587: dataIn1 = 32'd901
; 
32'd15588: dataIn1 = 32'd827
; 
32'd15589: dataIn1 = 32'd848
; 
32'd15590: dataIn1 = 32'd867
; 
32'd15591: dataIn1 = 32'd896
; 
32'd15592: dataIn1 = 32'd831
; 
32'd15593: dataIn1 = 32'd839
; 
32'd15594: dataIn1 = 32'd843
; 
32'd15595: dataIn1 = 32'd897
; 
32'd15596: dataIn1 = 32'd925
; 
32'd15597: dataIn1 = 32'd860
; 
32'd15598: dataIn1 = 32'd869
; 
32'd15599: dataIn1 = 32'd888
; 
32'd15600: dataIn1 = 32'd898
; 
32'd15601: dataIn1 = 32'd851
; 
32'd15602: dataIn1 = 32'd858
; 
32'd15603: dataIn1 = 32'd862
; 
32'd15604: dataIn1 = 32'd899
; 
32'd15605: dataIn1 = 32'd927
; 
32'd15606: dataIn1 = 32'd821
; 
32'd15607: dataIn1 = 32'd836
; 
32'd15608: dataIn1 = 32'd874
; 
32'd15609: dataIn1 = 32'd900
; 
32'd15610: dataIn1 = 32'd796
; 
32'd15611: dataIn1 = 32'd866
; 
32'd15612: dataIn1 = 32'd895
; 
32'd15613: dataIn1 = 32'd901
; 
32'd15614: dataIn1 = 32'd924
; 
32'd15615: dataIn1 = 32'd836
; 
32'd15616: dataIn1 = 32'd842
; 
32'd15617: dataIn1 = 32'd876
; 
32'd15618: dataIn1 = 32'd902
; 
32'd15619: dataIn1 = 32'd930
; 
32'd15620: dataIn1 = 32'd788
; 
32'd15621: dataIn1 = 32'd835
; 
32'd15622: dataIn1 = 32'd864
; 
32'd15623: dataIn1 = 32'd903
; 
32'd15624: dataIn1 = 32'd840
; 
32'd15625: dataIn1 = 32'd873
; 
32'd15626: dataIn1 = 32'd881
; 
32'd15627: dataIn1 = 32'd904
; 
32'd15628: dataIn1 = 32'd872
; 
32'd15629: dataIn1 = 32'd885
; 
32'd15630: dataIn1 = 32'd887
; 
32'd15631: dataIn1 = 32'd905
; 
32'd15632: dataIn1 = 32'd932
; 
32'd15633: dataIn1 = 32'd778
; 
32'd15634: dataIn1 = 32'd830
; 
32'd15635: dataIn1 = 32'd864
; 
32'd15636: dataIn1 = 32'd906
; 
32'd15637: dataIn1 = 32'd825
; 
32'd15638: dataIn1 = 32'd834
; 
32'd15639: dataIn1 = 32'd857
; 
32'd15640: dataIn1 = 32'd907
; 
32'd15641: dataIn1 = 32'd916
; 
32'd15642: dataIn1 = 32'd832
; 
32'd15643: dataIn1 = 32'd855
; 
32'd15644: dataIn1 = 32'd862
; 
32'd15645: dataIn1 = 32'd908
; 
32'd15646: dataIn1 = 32'd837
; 
32'd15647: dataIn1 = 32'd883
; 
32'd15648: dataIn1 = 32'd894
; 
32'd15649: dataIn1 = 32'd909
; 
32'd15650: dataIn1 = 32'd818
; 
32'd15651: dataIn1 = 32'd861
; 
32'd15652: dataIn1 = 32'd868
; 
32'd15653: dataIn1 = 32'd910
; 
32'd15654: dataIn1 = 32'd818
; 
32'd15655: dataIn1 = 32'd861
; 
32'd15656: dataIn1 = 32'd879
; 
32'd15657: dataIn1 = 32'd911
; 
32'd15658: dataIn1 = 32'd933
; 
32'd15659: dataIn1 = 32'd962
; 
32'd15660: dataIn1 = 32'd781
; 
32'd15661: dataIn1 = 32'd818
; 
32'd15662: dataIn1 = 32'd871
; 
32'd15663: dataIn1 = 32'd912
; 
32'd15664: dataIn1 = 32'd933
; 
32'd15665: dataIn1 = 32'd817
; 
32'd15666: dataIn1 = 32'd848
; 
32'd15667: dataIn1 = 32'd877
; 
32'd15668: dataIn1 = 32'd913
; 
32'd15669: dataIn1 = 32'd918
; 
32'd15670: dataIn1 = 32'd935
; 
32'd15671: dataIn1 = 32'd821
; 
32'd15672: dataIn1 = 32'd822
; 
32'd15673: dataIn1 = 32'd868
; 
32'd15674: dataIn1 = 32'd914
; 
32'd15675: dataIn1 = 32'd926
; 
32'd15676: dataIn1 = 32'd823
; 
32'd15677: dataIn1 = 32'd827
; 
32'd15678: dataIn1 = 32'd859
; 
32'd15679: dataIn1 = 32'd915
; 
32'd15680: dataIn1 = 32'd825
; 
32'd15681: dataIn1 = 32'd857
; 
32'd15682: dataIn1 = 32'd907
; 
32'd15683: dataIn1 = 32'd916
; 
32'd15684: dataIn1 = 32'd826
; 
32'd15685: dataIn1 = 32'd860
; 
32'd15686: dataIn1 = 32'd891
; 
32'd15687: dataIn1 = 32'd917
; 
32'd15688: dataIn1 = 32'd827
; 
32'd15689: dataIn1 = 32'd873
; 
32'd15690: dataIn1 = 32'd913
; 
32'd15691: dataIn1 = 32'd918
; 
32'd15692: dataIn1 = 32'd935
; 
32'd15693: dataIn1 = 32'd830
; 
32'd15694: dataIn1 = 32'd837
; 
32'd15695: dataIn1 = 32'd882
; 
32'd15696: dataIn1 = 32'd919
; 
32'd15697: dataIn1 = 32'd823
; 
32'd15698: dataIn1 = 32'd831
; 
32'd15699: dataIn1 = 32'd893
; 
32'd15700: dataIn1 = 32'd920
; 
32'd15701: dataIn1 = 32'd834
; 
32'd15702: dataIn1 = 32'd852
; 
32'd15703: dataIn1 = 32'd867
; 
32'd15704: dataIn1 = 32'd921
; 
32'd15705: dataIn1 = 32'd857
; 
32'd15706: dataIn1 = 32'd865
; 
32'd15707: dataIn1 = 32'd871
; 
32'd15708: dataIn1 = 32'd922
; 
32'd15709: dataIn1 = 32'd852
; 
32'd15710: dataIn1 = 32'd859
; 
32'd15711: dataIn1 = 32'd882
; 
32'd15712: dataIn1 = 32'd923
; 
32'd15713: dataIn1 = 32'd861
; 
32'd15714: dataIn1 = 32'd868
; 
32'd15715: dataIn1 = 32'd901
; 
32'd15716: dataIn1 = 32'd924
; 
32'd15717: dataIn1 = 32'd928
; 
32'd15718: dataIn1 = 32'd862
; 
32'd15719: dataIn1 = 32'd865
; 
32'd15720: dataIn1 = 32'd897
; 
32'd15721: dataIn1 = 32'd925
; 
32'd15722: dataIn1 = 32'd831
; 
32'd15723: dataIn1 = 32'd863
; 
32'd15724: dataIn1 = 32'd914
; 
32'd15725: dataIn1 = 32'd926
; 
32'd15726: dataIn1 = 32'd834
; 
32'd15727: dataIn1 = 32'd865
; 
32'd15728: dataIn1 = 32'd899
; 
32'd15729: dataIn1 = 32'd927
; 
32'd15730: dataIn1 = 32'd866
; 
32'd15731: dataIn1 = 32'd879
; 
32'd15732: dataIn1 = 32'd924
; 
32'd15733: dataIn1 = 32'd928
; 
32'd15734: dataIn1 = 32'd781
; 
32'd15735: dataIn1 = 32'd817
; 
32'd15736: dataIn1 = 32'd877
; 
32'd15737: dataIn1 = 32'd929
; 
32'd15738: dataIn1 = 32'd821
; 
32'd15739: dataIn1 = 32'd842
; 
32'd15740: dataIn1 = 32'd902
; 
32'd15741: dataIn1 = 32'd930
; 
32'd15742: dataIn1 = 32'd822
; 
32'd15743: dataIn1 = 32'd831
; 
32'd15744: dataIn1 = 32'd874
; 
32'd15745: dataIn1 = 32'd931
; 
32'd15746: dataIn1 = 32'd859
; 
32'd15747: dataIn1 = 32'd882
; 
32'd15748: dataIn1 = 32'd905
; 
32'd15749: dataIn1 = 32'd932
; 
32'd15750: dataIn1 = 32'd781
; 
32'd15751: dataIn1 = 32'd911
; 
32'd15752: dataIn1 = 32'd912
; 
32'd15753: dataIn1 = 32'd933
; 
32'd15754: dataIn1 = 32'd962
; 
32'd15755: dataIn1 = 32'd869
; 
32'd15756: dataIn1 = 32'd888
; 
32'd15757: dataIn1 = 32'd898
; 
32'd15758: dataIn1 = 32'd934
; 
32'd15759: dataIn1 = 32'd817
; 
32'd15760: dataIn1 = 32'd913
; 
32'd15761: dataIn1 = 32'd918
; 
32'd15762: dataIn1 = 32'd935
; 
32'd15763: dataIn1 = 32'd781
; 
32'd15764: dataIn1 = 32'd912
; 
32'd15765: dataIn1 = 32'd929
; 
32'd15766: dataIn1 = 32'd936
; 
32'd15767: dataIn1 = 32'd866
; 
32'd15768: dataIn1 = 32'd901
; 
32'd15769: dataIn1 = 32'd906
; 
32'd15770: dataIn1 = 32'd937
; 
32'd15771: dataIn1 = 32'd913
; 
32'd15772: dataIn1 = 32'd929
; 
32'd15773: dataIn1 = 32'd938
; 
32'd15774: dataIn1 = 32'd831
; 
32'd15775: dataIn1 = 32'd872
; 
32'd15776: dataIn1 = 32'd897
; 
32'd15777: dataIn1 = 32'd939
; 
32'd15778: dataIn1 = 32'd886
; 
32'd15779: dataIn1 = 32'd891
; 
32'd15780: dataIn1 = 32'd894
; 
32'd15781: dataIn1 = 32'd940
; 
32'd15782: dataIn1 = 32'd882
; 
32'd15783: dataIn1 = 32'd887
; 
32'd15784: dataIn1 = 32'd932
; 
32'd15785: dataIn1 = 32'd941
; 
32'd15786: dataIn1 = 32'd876
; 
32'd15787: dataIn1 = 32'd880
; 
32'd15788: dataIn1 = 32'd902
; 
32'd15789: dataIn1 = 32'd942
; 
32'd15790: dataIn1 = 32'd945
; 
32'd15791: dataIn1 = 32'd880
; 
32'd15792: dataIn1 = 32'd889
; 
32'd15793: dataIn1 = 32'd943
; 
32'd15794: dataIn1 = 32'd883
; 
32'd15795: dataIn1 = 32'd891
; 
32'd15796: dataIn1 = 32'd909
; 
32'd15797: dataIn1 = 32'd944
; 
32'd15798: dataIn1 = 32'd830
; 
32'd15799: dataIn1 = 32'd876
; 
32'd15800: dataIn1 = 32'd945
; 
32'd15801: dataIn1 = 32'd881
; 
32'd15802: dataIn1 = 32'd900
; 
32'd15803: dataIn1 = 32'd902
; 
32'd15804: dataIn1 = 32'd946
; 
32'd15805: dataIn1 = 32'd827
; 
32'd15806: dataIn1 = 32'd859
; 
32'd15807: dataIn1 = 32'd896
; 
32'd15808: dataIn1 = 32'd947
; 
32'd15809: dataIn1 = 32'd899
; 
32'd15810: dataIn1 = 32'd908
; 
32'd15811: dataIn1 = 32'd948
; 
32'd15812: dataIn1 = 32'd894
; 
32'd15813: dataIn1 = 32'd923
; 
32'd15814: dataIn1 = 32'd949
; 
32'd15815: dataIn1 = 32'd865
; 
32'd15816: dataIn1 = 32'd899
; 
32'd15817: dataIn1 = 32'd927
; 
32'd15818: dataIn1 = 32'd950
; 
32'd15819: dataIn1 = 32'd905
; 
32'd15820: dataIn1 = 32'd915
; 
32'd15821: dataIn1 = 32'd932
; 
32'd15822: dataIn1 = 32'd951
; 
32'd15823: dataIn1 = 32'd896
; 
32'd15824: dataIn1 = 32'd907
; 
32'd15825: dataIn1 = 32'd921
; 
32'd15826: dataIn1 = 32'd952
; 
32'd15827: dataIn1 = 32'd827
; 
32'd15828: dataIn1 = 32'd874
; 
32'd15829: dataIn1 = 32'd904
; 
32'd15830: dataIn1 = 32'd953
; 
32'd15831: dataIn1 = 32'd921
; 
32'd15832: dataIn1 = 32'd940
; 
32'd15833: dataIn1 = 32'd954
; 
32'd15834: dataIn1 = 32'd830
; 
32'd15835: dataIn1 = 32'd890
; 
32'd15836: dataIn1 = 32'd955
; 
32'd15837: dataIn1 = 32'd890
; 
32'd15838: dataIn1 = 32'd897
; 
32'd15839: dataIn1 = 32'd925
; 
32'd15840: dataIn1 = 32'd956
; 
32'd15841: dataIn1 = 32'd842
; 
32'd15842: dataIn1 = 32'd902
; 
32'd15843: dataIn1 = 32'd945
; 
32'd15844: dataIn1 = 32'd957
; 
32'd15845: dataIn1 = 32'd893
; 
32'd15846: dataIn1 = 32'd920
; 
32'd15847: dataIn1 = 32'd958
; 
32'd15848: dataIn1 = 32'd821
; 
32'd15849: dataIn1 = 32'd868
; 
32'd15850: dataIn1 = 32'd914
; 
32'd15851: dataIn1 = 32'd959
; 
32'd15852: dataIn1 = 32'd895
; 
32'd15853: dataIn1 = 32'd901
; 
32'd15854: dataIn1 = 32'd960
; 
32'd15855: dataIn1 = 32'd862
; 
32'd15856: dataIn1 = 32'd903
; 
32'd15857: dataIn1 = 32'd961
; 
32'd15858: dataIn1 = 32'd888
; 
32'd15859: dataIn1 = 32'd911
; 
32'd15860: dataIn1 = 32'd933
; 
32'd15861: dataIn1 = 32'd962
; 
32'd15862: dataIn1 = 32'd871
; 
32'd15863: dataIn1 = 32'd916
; 
32'd15864: dataIn1 = 32'd963
; 
32'd15865: dataIn1 = 32'd821
; 
32'd15866: dataIn1 = 32'd874
; 
32'd15867: dataIn1 = 32'd914
; 
32'd15868: dataIn1 = 32'd964
; 
32'd15869: dataIn1 = 32'd830
; 
32'd15870: dataIn1 = 32'd890
; 
32'd15871: dataIn1 = 32'd965
; 
32'd15872: dataIn1 = 32'd834
; 
32'd15873: dataIn1 = 32'd907
; 
32'd15874: dataIn1 = 32'd927
; 
32'd15875: dataIn1 = 32'd966
; 
32'd15876: dataIn1 = 32'd859
; 
32'd15877: dataIn1 = 32'd896
; 
32'd15878: dataIn1 = 32'd921
; 
32'd15879: dataIn1 = 32'd967
; 
32'd15880: dataIn1 = 32'd860
; 
32'd15881: dataIn1 = 32'd879
; 
32'd15882: dataIn1 = 32'd962
; 
32'd15883: dataIn1 = 32'd968
; 
32'd15884: dataIn1 = 32'd863
; 
32'd15885: dataIn1 = 32'd868
; 
32'd15886: dataIn1 = 32'd910
; 
32'd15887: dataIn1 = 32'd969
; 
32'd15888: dataIn1 = 32'd866
; 
32'd15889: dataIn1 = 32'd903
; 
32'd15890: dataIn1 = 32'd906
; 
32'd15891: dataIn1 = 32'd970
; 
32'd15892: dataIn1 = 32'd863
; 
32'd15893: dataIn1 = 32'd871
; 
32'd15894: dataIn1 = 32'd912
; 
32'd15895: dataIn1 = 32'd971
; 
32'd15896: dataIn1 = 32'd872
; 
32'd15897: dataIn1 = 32'd905
; 
32'd15898: dataIn1 = 32'd972
; 
32'd15899: dataIn1 = 32'd874
; 
32'd15900: dataIn1 = 32'd904
; 
32'd15901: dataIn1 = 32'd973
; 
32'd15902: dataIn1 = 32'd855
; 
32'd15903: dataIn1 = 32'd866
; 
32'd15904: dataIn1 = 32'd879
; 
32'd15905: dataIn1 = 32'd974
; 
32'd15906: dataIn1 = 32'd880
; 
32'd15907: dataIn1 = 32'd881
; 
32'd15908: dataIn1 = 32'd975
; 
32'd15909: dataIn1 = 32'd881
; 
32'd15910: dataIn1 = 32'd889
; 
32'd15911: dataIn1 = 32'd904
; 
32'd15912: dataIn1 = 32'd976
; 
32'd15913: dataIn1 = 32'd896
; 
32'd15914: dataIn1 = 32'd918
; 
32'd15915: dataIn1 = 32'd977
; 
32'd15916: dataIn1 = 32'd863
; 
32'd15917: dataIn1 = 32'd897
; 
32'd15918: dataIn1 = 32'd926
; 
32'd15919: dataIn1 = 32'd978
; 
32'd15920: dataIn1 = 32'd900
; 
32'd15921: dataIn1 = 32'd930
; 
32'd15922: dataIn1 = 32'd979
; 
32'd15923: dataIn1 = 32'd901
; 
32'd15924: dataIn1 = 32'd928
; 
32'd15925: dataIn1 = 32'd980
; 
32'd15926: dataIn1 = 32'd904
; 
32'd15927: dataIn1 = 32'd918
; 
32'd15928: dataIn1 = 32'd981
; 
32'd15929: dataIn1 = 32'd911
; 
32'd15930: dataIn1 = 32'd982
; 
32'd15931: dataIn1 = 32'd871
; 
32'd15932: dataIn1 = 32'd912
; 
32'd15933: dataIn1 = 32'd983
; 
32'd15934: dataIn1 = 32'd896
; 
32'd15935: dataIn1 = 32'd913
; 
32'd15936: dataIn1 = 32'd984
; 
32'd15937: dataIn1 = 32'd923
; 
32'd15938: dataIn1 = 32'd932
; 
32'd15939: dataIn1 = 32'd985
; 
32'd15940: dataIn1 = 32'd911
; 
32'd15941: dataIn1 = 32'd912
; 
32'd15942: dataIn1 = 32'd933
; 
32'd15943: dataIn1 = 32'd986
; 
32'd15944: dataIn1 = 32'd834
; 
32'd15945: dataIn1 = 32'd987
; 
32'd15946: dataIn1 = 32'd859
; 
32'd15947: dataIn1 = 32'd923
; 
32'd15948: dataIn1 = 32'd988
; 
32'd15949: dataIn1 = 32'd863
; 
32'd15950: dataIn1 = 32'd926
; 
32'd15951: dataIn1 = 32'd989
; 
32'd15952: dataIn1 = 32'd859
; 
32'd15953: dataIn1 = 32'd915
; 
32'd15954: dataIn1 = 32'd990
; 
32'd15955: dataIn1 = 32'd863
; 
32'd15956: dataIn1 = 32'd991
; 
default:  
	dataIn1 = 32'd99999; 
endcase 
case(addr2) 
32'd2: dataIn2 = 32'd0; 
32'd3: dataIn2 = 32'd1; 
32'd4: dataIn2 = 32'd0; 
32'd5: dataIn2 = 32'd0; 
32'd6: dataIn2 = 32'd1; 
32'd7: dataIn2 = 32'd1; 
32'd8: dataIn2 = 32'd1; 
32'd9: dataIn2 = 32'd0; 
32'd10: dataIn2 = 32'd1; 
32'd11: dataIn2 = 32'd1; 
32'd12: dataIn2 = 32'd1; 
32'd13: dataIn2 = 32'd0; 
32'd14: dataIn2 = 32'd0; 
32'd15: dataIn2 = 32'd0; 
32'd16: dataIn2 = 32'd0; 
32'd17: dataIn2 = 32'd1; 
32'd18: dataIn2 = 32'd1; 
32'd19: dataIn2 = 32'd0; 
32'd20: dataIn2 = 32'd1; 
32'd21: dataIn2 = 32'd0; 
32'd22: dataIn2 = 32'd0; 
32'd23: dataIn2 = 32'd0; 
32'd24: dataIn2 = 32'd1; 
32'd25: dataIn2 = 32'd1; 
32'd26: dataIn2 = 32'd1; 
32'd27: dataIn2 = 32'd1; 
32'd28: dataIn2 = 32'd1; 
32'd29: dataIn2 = 32'd1; 
32'd30: dataIn2 = 32'd1; 
32'd31: dataIn2 = 32'd0; 
32'd32: dataIn2 = 32'd1; 
32'd33: dataIn2 = 32'd1; 
32'd34: dataIn2 = 32'd0; 
32'd35: dataIn2 = 32'd0; 
32'd36: dataIn2 = 32'd0; 
32'd37: dataIn2 = 32'd0; 
32'd38: dataIn2 = 32'd0; 
32'd39: dataIn2 = 32'd0; 
32'd40: dataIn2 = 32'd0; 
32'd41: dataIn2 = 32'd0; 
32'd42: dataIn2 = 32'd0; 
32'd43: dataIn2 = 32'd0; 
32'd44: dataIn2 = 32'd0; 
32'd45: dataIn2 = 32'd0; 
32'd46: dataIn2 = 32'd1; 
32'd47: dataIn2 = 32'd0; 
32'd48: dataIn2 = 32'd0; 
32'd49: dataIn2 = 32'd0; 
32'd50: dataIn2 = 32'd0; 
32'd51: dataIn2 = 32'd1; 
32'd52: dataIn2 = 32'd0; 
32'd53: dataIn2 = 32'd0; 
32'd54: dataIn2 = 32'd1; 
32'd55: dataIn2 = 32'd1; 
32'd56: dataIn2 = 32'd1; 
32'd57: dataIn2 = 32'd1; 
32'd58: dataIn2 = 32'd1; 
32'd59: dataIn2 = 32'd1; 
32'd60: dataIn2 = 32'd0; 
32'd61: dataIn2 = 32'd0; 
32'd62: dataIn2 = 32'd0; 
32'd63: dataIn2 = 32'd1; 
32'd64: dataIn2 = 32'd1; 
32'd65: dataIn2 = 32'd0; 
32'd66: dataIn2 = 32'd0; 
32'd67: dataIn2 = 32'd0; 
32'd68: dataIn2 = 32'd0; 
32'd69: dataIn2 = 32'd0; 
32'd70: dataIn2 = 32'd0; 
32'd71: dataIn2 = 32'd0; 
32'd72: dataIn2 = 32'd0; 
32'd73: dataIn2 = 32'd0; 
32'd74: dataIn2 = 32'd1; 
32'd75: dataIn2 = 32'd1; 
32'd76: dataIn2 = 32'd1; 
32'd77: dataIn2 = 32'd0; 
32'd78: dataIn2 = 32'd0; 
32'd79: dataIn2 = 32'd0; 
32'd80: dataIn2 = 32'd0; 
32'd81: dataIn2 = 32'd0; 
32'd82: dataIn2 = 32'd0; 
32'd83: dataIn2 = 32'd0; 
32'd84: dataIn2 = 32'd0; 
32'd85: dataIn2 = 32'd0; 
32'd86: dataIn2 = 32'd1; 
32'd87: dataIn2 = 32'd0; 
32'd88: dataIn2 = 32'd0; 
32'd89: dataIn2 = 32'd1; 
32'd90: dataIn2 = 32'd1; 
32'd91: dataIn2 = 32'd1; 
32'd92: dataIn2 = 32'd1; 
32'd93: dataIn2 = 32'd1; 
32'd94: dataIn2 = 32'd0; 
32'd95: dataIn2 = 32'd0; 
32'd96: dataIn2 = 32'd0; 
32'd97: dataIn2 = 32'd1; 
32'd98: dataIn2 = 32'd0; 
32'd99: dataIn2 = 32'd0; 
32'd100: dataIn2 = 32'd0; 
32'd101: dataIn2 = 32'd1; 
32'd102: dataIn2 = 32'd0; 
32'd103: dataIn2 = 32'd1; 
32'd104: dataIn2 = 32'd1; 
32'd105: dataIn2 = 32'd1; 
32'd106: dataIn2 = 32'd0; 
32'd107: dataIn2 = 32'd0; 
32'd108: dataIn2 = 32'd0; 
32'd109: dataIn2 = 32'd0; 
32'd110: dataIn2 = 32'd0; 
32'd111: dataIn2 = 32'd0; 
32'd112: dataIn2 = 32'd1; 
32'd113: dataIn2 = 32'd0; 
32'd114: dataIn2 = 32'd1; 
32'd115: dataIn2 = 32'd0; 
32'd116: dataIn2 = 32'd0; 
32'd117: dataIn2 = 32'd1; 
32'd118: dataIn2 = 32'd0; 
32'd119: dataIn2 = 32'd0; 
32'd120: dataIn2 = 32'd0; 
32'd121: dataIn2 = 32'd1; 
32'd122: dataIn2 = 32'd1; 
32'd123: dataIn2 = 32'd0; 
32'd124: dataIn2 = 32'd0; 
32'd125: dataIn2 = 32'd0; 
32'd126: dataIn2 = 32'd1; 
32'd127: dataIn2 = 32'd1; 
32'd128: dataIn2 = 32'd1; 
32'd129: dataIn2 = 32'd0; 
32'd130: dataIn2 = 32'd0; 
32'd131: dataIn2 = 32'd0; 
32'd132: dataIn2 = 32'd0; 
32'd133: dataIn2 = 32'd1; 
32'd134: dataIn2 = 32'd1; 
32'd135: dataIn2 = 32'd1; 
32'd136: dataIn2 = 32'd1; 
32'd137: dataIn2 = 32'd1; 
32'd138: dataIn2 = 32'd1; 
32'd139: dataIn2 = 32'd0; 
32'd140: dataIn2 = 32'd0; 
32'd141: dataIn2 = 32'd0; 
32'd142: dataIn2 = 32'd0; 
32'd143: dataIn2 = 32'd1; 
32'd144: dataIn2 = 32'd1; 
32'd145: dataIn2 = 32'd1; 
32'd146: dataIn2 = 32'd0; 
32'd147: dataIn2 = 32'd1; 
32'd148: dataIn2 = 32'd1; 
32'd149: dataIn2 = 32'd0; 
32'd150: dataIn2 = 32'd1; 
32'd151: dataIn2 = 32'd1; 
32'd152: dataIn2 = 32'd0; 
32'd153: dataIn2 = 32'd1; 
32'd154: dataIn2 = 32'd1; 
32'd155: dataIn2 = 32'd1; 
32'd156: dataIn2 = 32'd0; 
32'd157: dataIn2 = 32'd1; 
32'd158: dataIn2 = 32'd0; 
32'd159: dataIn2 = 32'd0; 
32'd160: dataIn2 = 32'd0; 
32'd161: dataIn2 = 32'd1; 
32'd162: dataIn2 = 32'd0; 
32'd163: dataIn2 = 32'd0; 
32'd164: dataIn2 = 32'd1; 
32'd165: dataIn2 = 32'd0; 
32'd166: dataIn2 = 32'd1; 
32'd167: dataIn2 = 32'd0; 
32'd168: dataIn2 = 32'd0; 
32'd169: dataIn2 = 32'd1; 
32'd170: dataIn2 = 32'd1; 
32'd171: dataIn2 = 32'd1; 
32'd172: dataIn2 = 32'd1; 
32'd173: dataIn2 = 32'd1; 
32'd174: dataIn2 = 32'd1; 
32'd175: dataIn2 = 32'd0; 
32'd176: dataIn2 = 32'd0; 
32'd177: dataIn2 = 32'd1; 
32'd178: dataIn2 = 32'd0; 
32'd179: dataIn2 = 32'd0; 
32'd180: dataIn2 = 32'd0; 
32'd181: dataIn2 = 32'd1; 
32'd182: dataIn2 = 32'd1; 
32'd183: dataIn2 = 32'd0; 
32'd184: dataIn2 = 32'd0; 
32'd185: dataIn2 = 32'd1; 
32'd186: dataIn2 = 32'd1; 
32'd187: dataIn2 = 32'd1; 
32'd188: dataIn2 = 32'd0; 
32'd189: dataIn2 = 32'd1; 
32'd190: dataIn2 = 32'd1; 
32'd191: dataIn2 = 32'd0; 
32'd192: dataIn2 = 32'd1; 
32'd193: dataIn2 = 32'd1; 
32'd194: dataIn2 = 32'd0; 
32'd195: dataIn2 = 32'd0; 
32'd196: dataIn2 = 32'd1; 
32'd197: dataIn2 = 32'd0; 
32'd198: dataIn2 = 32'd0; 
32'd199: dataIn2 = 32'd0; 
32'd200: dataIn2 = 32'd0; 
32'd201: dataIn2 = 32'd1; 
32'd202: dataIn2 = 32'd0; 
32'd203: dataIn2 = 32'd0; 
32'd204: dataIn2 = 32'd0; 
32'd205: dataIn2 = 32'd1; 
32'd206: dataIn2 = 32'd1; 
32'd207: dataIn2 = 32'd0; 
32'd208: dataIn2 = 32'd1; 
32'd209: dataIn2 = 32'd0; 
32'd210: dataIn2 = 32'd1; 
32'd211: dataIn2 = 32'd0; 
32'd212: dataIn2 = 32'd1; 
32'd213: dataIn2 = 32'd1; 
32'd214: dataIn2 = 32'd0; 
32'd215: dataIn2 = 32'd0; 
32'd216: dataIn2 = 32'd0; 
32'd217: dataIn2 = 32'd0; 
32'd218: dataIn2 = 32'd1; 
32'd219: dataIn2 = 32'd1; 
32'd220: dataIn2 = 32'd1; 
32'd221: dataIn2 = 32'd1; 
32'd222: dataIn2 = 32'd0; 
32'd223: dataIn2 = 32'd1; 
32'd224: dataIn2 = 32'd1; 
32'd225: dataIn2 = 32'd0; 
32'd226: dataIn2 = 32'd0; 
32'd227: dataIn2 = 32'd1; 
32'd228: dataIn2 = 32'd1; 
32'd229: dataIn2 = 32'd0; 
32'd230: dataIn2 = 32'd0; 
32'd231: dataIn2 = 32'd1; 
32'd232: dataIn2 = 32'd1; 
32'd233: dataIn2 = 32'd0; 
32'd234: dataIn2 = 32'd0; 
32'd235: dataIn2 = 32'd1; 
32'd236: dataIn2 = 32'd0; 
32'd237: dataIn2 = 32'd1; 
32'd238: dataIn2 = 32'd0; 
32'd239: dataIn2 = 32'd1; 
32'd240: dataIn2 = 32'd0; 
32'd241: dataIn2 = 32'd0; 
32'd242: dataIn2 = 32'd1; 
32'd243: dataIn2 = 32'd1; 
32'd244: dataIn2 = 32'd1; 
32'd245: dataIn2 = 32'd1; 
32'd246: dataIn2 = 32'd0; 
32'd247: dataIn2 = 32'd0; 
32'd248: dataIn2 = 32'd1; 
32'd249: dataIn2 = 32'd0; 
32'd250: dataIn2 = 32'd1; 
32'd251: dataIn2 = 32'd0; 
32'd252: dataIn2 = 32'd1; 
32'd253: dataIn2 = 32'd1; 
32'd254: dataIn2 = 32'd1; 
32'd255: dataIn2 = 32'd0; 
32'd256: dataIn2 = 32'd0; 
32'd257: dataIn2 = 32'd0; 
32'd258: dataIn2 = 32'd1; 
32'd259: dataIn2 = 32'd0; 
32'd260: dataIn2 = 32'd0; 
32'd261: dataIn2 = 32'd0; 
32'd262: dataIn2 = 32'd0; 
32'd263: dataIn2 = 32'd1; 
32'd264: dataIn2 = 32'd1; 
32'd265: dataIn2 = 32'd1; 
32'd266: dataIn2 = 32'd0; 
32'd267: dataIn2 = 32'd1; 
32'd268: dataIn2 = 32'd0; 
32'd269: dataIn2 = 32'd0; 
32'd270: dataIn2 = 32'd0; 
32'd271: dataIn2 = 32'd1; 
32'd272: dataIn2 = 32'd1; 
32'd273: dataIn2 = 32'd0; 
32'd274: dataIn2 = 32'd1; 
32'd275: dataIn2 = 32'd1; 
32'd276: dataIn2 = 32'd0; 
32'd277: dataIn2 = 32'd0; 
32'd278: dataIn2 = 32'd1; 
32'd279: dataIn2 = 32'd0; 
32'd280: dataIn2 = 32'd1; 
32'd281: dataIn2 = 32'd0; 
32'd282: dataIn2 = 32'd1; 
32'd283: dataIn2 = 32'd0; 
32'd284: dataIn2 = 32'd1; 
32'd285: dataIn2 = 32'd0; 
32'd286: dataIn2 = 32'd1; 
32'd287: dataIn2 = 32'd1; 
32'd288: dataIn2 = 32'd0; 
32'd289: dataIn2 = 32'd1; 
32'd290: dataIn2 = 32'd0; 
32'd291: dataIn2 = 32'd1; 
32'd292: dataIn2 = 32'd1; 
32'd293: dataIn2 = 32'd0; 
32'd294: dataIn2 = 32'd0; 
32'd295: dataIn2 = 32'd1; 
32'd296: dataIn2 = 32'd1; 
32'd297: dataIn2 = 32'd1; 
32'd298: dataIn2 = 32'd1; 
32'd299: dataIn2 = 32'd1; 
32'd300: dataIn2 = 32'd0; 
32'd301: dataIn2 = 32'd1; 
32'd302: dataIn2 = 32'd1; 
32'd303: dataIn2 = 32'd0; 
32'd304: dataIn2 = 32'd1; 
32'd305: dataIn2 = 32'd0; 
32'd306: dataIn2 = 32'd1; 
32'd307: dataIn2 = 32'd0; 
32'd308: dataIn2 = 32'd0; 
32'd309: dataIn2 = 32'd1; 
32'd310: dataIn2 = 32'd0; 
32'd311: dataIn2 = 32'd1; 
32'd312: dataIn2 = 32'd0; 
32'd313: dataIn2 = 32'd1; 
32'd314: dataIn2 = 32'd1; 
32'd315: dataIn2 = 32'd0; 
32'd316: dataIn2 = 32'd1; 
32'd317: dataIn2 = 32'd1; 
32'd318: dataIn2 = 32'd1; 
32'd319: dataIn2 = 32'd0; 
32'd320: dataIn2 = 32'd0; 
32'd321: dataIn2 = 32'd1; 
32'd322: dataIn2 = 32'd0; 
32'd323: dataIn2 = 32'd1; 
32'd324: dataIn2 = 32'd0; 
32'd325: dataIn2 = 32'd0; 
32'd326: dataIn2 = 32'd1; 
32'd327: dataIn2 = 32'd0; 
32'd328: dataIn2 = 32'd0; 
32'd329: dataIn2 = 32'd1; 
32'd330: dataIn2 = 32'd1; 
32'd331: dataIn2 = 32'd1; 
32'd332: dataIn2 = 32'd1; 
32'd333: dataIn2 = 32'd1; 
32'd334: dataIn2 = 32'd1; 
32'd335: dataIn2 = 32'd0; 
32'd336: dataIn2 = 32'd0; 
32'd337: dataIn2 = 32'd1; 
32'd338: dataIn2 = 32'd0; 
32'd339: dataIn2 = 32'd0; 
32'd340: dataIn2 = 32'd0; 
32'd341: dataIn2 = 32'd0; 
32'd342: dataIn2 = 32'd1; 
32'd343: dataIn2 = 32'd1; 
32'd344: dataIn2 = 32'd1; 
32'd345: dataIn2 = 32'd1; 
32'd346: dataIn2 = 32'd1; 
32'd347: dataIn2 = 32'd0; 
32'd348: dataIn2 = 32'd0; 
32'd349: dataIn2 = 32'd0; 
32'd350: dataIn2 = 32'd1; 
32'd351: dataIn2 = 32'd0; 
32'd352: dataIn2 = 32'd0; 
32'd353: dataIn2 = 32'd0; 
32'd354: dataIn2 = 32'd0; 
32'd355: dataIn2 = 32'd0; 
32'd356: dataIn2 = 32'd0; 
32'd357: dataIn2 = 32'd0; 
32'd358: dataIn2 = 32'd1; 
32'd359: dataIn2 = 32'd1; 
32'd360: dataIn2 = 32'd1; 
32'd361: dataIn2 = 32'd1; 
32'd362: dataIn2 = 32'd0; 
32'd363: dataIn2 = 32'd0; 
32'd364: dataIn2 = 32'd1; 
32'd365: dataIn2 = 32'd1; 
32'd366: dataIn2 = 32'd1; 
32'd367: dataIn2 = 32'd0; 
32'd368: dataIn2 = 32'd0; 
32'd369: dataIn2 = 32'd1; 
32'd370: dataIn2 = 32'd0; 
32'd371: dataIn2 = 32'd1; 
32'd372: dataIn2 = 32'd0; 
32'd373: dataIn2 = 32'd1; 
32'd374: dataIn2 = 32'd0; 
32'd375: dataIn2 = 32'd0; 
32'd376: dataIn2 = 32'd0; 
32'd377: dataIn2 = 32'd0; 
32'd378: dataIn2 = 32'd1; 
32'd379: dataIn2 = 32'd1; 
32'd380: dataIn2 = 32'd0; 
32'd381: dataIn2 = 32'd1; 
32'd382: dataIn2 = 32'd1; 
32'd383: dataIn2 = 32'd1; 
32'd384: dataIn2 = 32'd1; 
32'd385: dataIn2 = 32'd1; 
32'd386: dataIn2 = 32'd0; 
32'd387: dataIn2 = 32'd0; 
32'd388: dataIn2 = 32'd1; 
32'd389: dataIn2 = 32'd0; 
32'd390: dataIn2 = 32'd1; 
32'd391: dataIn2 = 32'd0; 
32'd392: dataIn2 = 32'd1; 
32'd393: dataIn2 = 32'd0; 
32'd394: dataIn2 = 32'd0; 
32'd395: dataIn2 = 32'd1; 
32'd396: dataIn2 = 32'd1; 
32'd397: dataIn2 = 32'd1; 
32'd398: dataIn2 = 32'd0; 
32'd399: dataIn2 = 32'd0; 
32'd400: dataIn2 = 32'd0; 
32'd401: dataIn2 = 32'd0; 
32'd402: dataIn2 = 32'd1; 
32'd403: dataIn2 = 32'd0; 
32'd404: dataIn2 = 32'd1; 
32'd405: dataIn2 = 32'd1; 
32'd406: dataIn2 = 32'd1; 
32'd407: dataIn2 = 32'd0; 
32'd408: dataIn2 = 32'd1; 
32'd409: dataIn2 = 32'd0; 
32'd410: dataIn2 = 32'd1; 
32'd411: dataIn2 = 32'd0; 
32'd412: dataIn2 = 32'd0; 
32'd413: dataIn2 = 32'd1; 
32'd414: dataIn2 = 32'd0; 
32'd415: dataIn2 = 32'd0; 
32'd416: dataIn2 = 32'd1; 
32'd417: dataIn2 = 32'd1; 
32'd418: dataIn2 = 32'd0; 
32'd419: dataIn2 = 32'd1; 
32'd420: dataIn2 = 32'd0; 
32'd421: dataIn2 = 32'd0; 
32'd422: dataIn2 = 32'd1; 
32'd423: dataIn2 = 32'd1; 
32'd424: dataIn2 = 32'd1; 
32'd425: dataIn2 = 32'd0; 
32'd426: dataIn2 = 32'd0; 
32'd427: dataIn2 = 32'd0; 
32'd428: dataIn2 = 32'd1; 
32'd429: dataIn2 = 32'd1; 
32'd430: dataIn2 = 32'd1; 
32'd431: dataIn2 = 32'd1; 
32'd432: dataIn2 = 32'd0; 
32'd433: dataIn2 = 32'd1; 
32'd434: dataIn2 = 32'd0; 
32'd435: dataIn2 = 32'd0; 
32'd436: dataIn2 = 32'd0; 
32'd437: dataIn2 = 32'd0; 
32'd438: dataIn2 = 32'd1; 
32'd439: dataIn2 = 32'd1; 
32'd440: dataIn2 = 32'd1; 
32'd441: dataIn2 = 32'd1; 
32'd442: dataIn2 = 32'd0; 
32'd443: dataIn2 = 32'd0; 
32'd444: dataIn2 = 32'd1; 
32'd445: dataIn2 = 32'd0; 
32'd446: dataIn2 = 32'd1; 
32'd447: dataIn2 = 32'd0; 
32'd448: dataIn2 = 32'd1; 
32'd449: dataIn2 = 32'd1; 
32'd450: dataIn2 = 32'd1; 
32'd451: dataIn2 = 32'd0; 
32'd452: dataIn2 = 32'd1; 
32'd453: dataIn2 = 32'd1; 
32'd454: dataIn2 = 32'd0; 
32'd455: dataIn2 = 32'd1; 
32'd456: dataIn2 = 32'd1; 
32'd457: dataIn2 = 32'd0; 
32'd458: dataIn2 = 32'd1; 
32'd459: dataIn2 = 32'd1; 
32'd460: dataIn2 = 32'd0; 
32'd461: dataIn2 = 32'd0; 
32'd462: dataIn2 = 32'd0; 
32'd463: dataIn2 = 32'd0; 
32'd464: dataIn2 = 32'd1; 
32'd465: dataIn2 = 32'd1; 
32'd466: dataIn2 = 32'd1; 
32'd467: dataIn2 = 32'd0; 
32'd468: dataIn2 = 32'd0; 
32'd469: dataIn2 = 32'd1; 
32'd470: dataIn2 = 32'd0; 
32'd471: dataIn2 = 32'd0; 
32'd472: dataIn2 = 32'd1; 
32'd473: dataIn2 = 32'd1; 
32'd474: dataIn2 = 32'd0; 
32'd475: dataIn2 = 32'd1; 
32'd476: dataIn2 = 32'd0; 
32'd477: dataIn2 = 32'd1; 
32'd478: dataIn2 = 32'd1; 
32'd479: dataIn2 = 32'd0; 
32'd480: dataIn2 = 32'd1; 
32'd481: dataIn2 = 32'd0; 
32'd482: dataIn2 = 32'd1; 
32'd483: dataIn2 = 32'd1; 
32'd484: dataIn2 = 32'd1; 
32'd485: dataIn2 = 32'd0; 
32'd486: dataIn2 = 32'd1; 
32'd487: dataIn2 = 32'd0; 
32'd488: dataIn2 = 32'd1; 
32'd489: dataIn2 = 32'd1; 
32'd490: dataIn2 = 32'd1; 
32'd491: dataIn2 = 32'd1; 
32'd492: dataIn2 = 32'd0; 
32'd493: dataIn2 = 32'd0; 
32'd494: dataIn2 = 32'd0; 
32'd495: dataIn2 = 32'd1; 
32'd496: dataIn2 = 32'd0; 
32'd497: dataIn2 = 32'd0; 
32'd498: dataIn2 = 32'd0; 
32'd499: dataIn2 = 32'd0; 
32'd500: dataIn2 = 32'd0; 
32'd501: dataIn2 = 32'd0; 
32'd502: dataIn2 = 32'd1; 
32'd503: dataIn2 = 32'd1; 
32'd504: dataIn2 = 32'd0; 
32'd505: dataIn2 = 32'd1; 
32'd506: dataIn2 = 32'd1; 
32'd507: dataIn2 = 32'd0; 
32'd508: dataIn2 = 32'd1; 
32'd509: dataIn2 = 32'd1; 
32'd510: dataIn2 = 32'd0; 
32'd511: dataIn2 = 32'd0; 
32'd512: dataIn2 = 32'd1; 
32'd513: dataIn2 = 32'd0; 
32'd514: dataIn2 = 32'd0; 
32'd515: dataIn2 = 32'd0; 
32'd516: dataIn2 = 32'd0; 
32'd517: dataIn2 = 32'd1; 
32'd518: dataIn2 = 32'd1; 
32'd519: dataIn2 = 32'd0; 
32'd520: dataIn2 = 32'd0; 
32'd521: dataIn2 = 32'd1; 
32'd522: dataIn2 = 32'd0; 
32'd523: dataIn2 = 32'd1; 
32'd524: dataIn2 = 32'd1; 
32'd525: dataIn2 = 32'd0; 
32'd526: dataIn2 = 32'd1; 
32'd527: dataIn2 = 32'd1; 
32'd528: dataIn2 = 32'd0; 
32'd529: dataIn2 = 32'd1; 
32'd530: dataIn2 = 32'd1; 
32'd531: dataIn2 = 32'd1; 
32'd532: dataIn2 = 32'd1; 
32'd533: dataIn2 = 32'd0; 
32'd534: dataIn2 = 32'd0; 
32'd535: dataIn2 = 32'd0; 
32'd536: dataIn2 = 32'd1; 
32'd537: dataIn2 = 32'd1; 
32'd538: dataIn2 = 32'd1; 
32'd539: dataIn2 = 32'd1; 
32'd540: dataIn2 = 32'd0; 
32'd541: dataIn2 = 32'd1; 
32'd542: dataIn2 = 32'd0; 
32'd543: dataIn2 = 32'd0; 
32'd544: dataIn2 = 32'd1; 
32'd545: dataIn2 = 32'd1; 
32'd546: dataIn2 = 32'd0; 
32'd547: dataIn2 = 32'd0; 
32'd548: dataIn2 = 32'd0; 
32'd549: dataIn2 = 32'd0; 
32'd550: dataIn2 = 32'd1; 
32'd551: dataIn2 = 32'd1; 
32'd552: dataIn2 = 32'd1; 
32'd553: dataIn2 = 32'd0; 
32'd554: dataIn2 = 32'd0; 
32'd555: dataIn2 = 32'd1; 
32'd556: dataIn2 = 32'd1; 
32'd557: dataIn2 = 32'd0; 
32'd558: dataIn2 = 32'd1; 
32'd559: dataIn2 = 32'd0; 
32'd560: dataIn2 = 32'd0; 
32'd561: dataIn2 = 32'd1; 
32'd562: dataIn2 = 32'd1; 
32'd563: dataIn2 = 32'd1; 
32'd564: dataIn2 = 32'd1; 
32'd565: dataIn2 = 32'd0; 
32'd566: dataIn2 = 32'd1; 
32'd567: dataIn2 = 32'd1; 
32'd568: dataIn2 = 32'd0; 
32'd569: dataIn2 = 32'd0; 
32'd570: dataIn2 = 32'd0; 
32'd571: dataIn2 = 32'd1; 
32'd572: dataIn2 = 32'd1; 
32'd573: dataIn2 = 32'd1; 
32'd574: dataIn2 = 32'd1; 
32'd575: dataIn2 = 32'd0; 
32'd576: dataIn2 = 32'd0; 
32'd577: dataIn2 = 32'd1; 
32'd578: dataIn2 = 32'd1; 
32'd579: dataIn2 = 32'd0; 
32'd580: dataIn2 = 32'd1; 
32'd581: dataIn2 = 32'd1; 
32'd582: dataIn2 = 32'd0; 
32'd583: dataIn2 = 32'd1; 
32'd584: dataIn2 = 32'd0; 
32'd585: dataIn2 = 32'd0; 
32'd586: dataIn2 = 32'd1; 
32'd587: dataIn2 = 32'd1; 
32'd588: dataIn2 = 32'd0; 
32'd589: dataIn2 = 32'd0; 
32'd590: dataIn2 = 32'd1; 
32'd591: dataIn2 = 32'd0; 
32'd592: dataIn2 = 32'd0; 
32'd593: dataIn2 = 32'd0; 
32'd594: dataIn2 = 32'd1; 
32'd595: dataIn2 = 32'd1; 
32'd596: dataIn2 = 32'd0; 
32'd597: dataIn2 = 32'd1; 
32'd598: dataIn2 = 32'd0; 
32'd599: dataIn2 = 32'd1; 
32'd600: dataIn2 = 32'd1; 
32'd601: dataIn2 = 32'd0; 
32'd602: dataIn2 = 32'd1; 
32'd603: dataIn2 = 32'd1; 
32'd604: dataIn2 = 32'd0; 
32'd605: dataIn2 = 32'd0; 
32'd606: dataIn2 = 32'd1; 
32'd607: dataIn2 = 32'd1; 
32'd608: dataIn2 = 32'd1; 
32'd609: dataIn2 = 32'd1; 
32'd610: dataIn2 = 32'd1; 
32'd611: dataIn2 = 32'd1; 
32'd612: dataIn2 = 32'd1; 
32'd613: dataIn2 = 32'd1; 
32'd614: dataIn2 = 32'd1; 
32'd615: dataIn2 = 32'd0; 
32'd616: dataIn2 = 32'd0; 
32'd617: dataIn2 = 32'd0; 
32'd618: dataIn2 = 32'd1; 
32'd619: dataIn2 = 32'd1; 
32'd620: dataIn2 = 32'd0; 
32'd621: dataIn2 = 32'd0; 
32'd622: dataIn2 = 32'd0; 
32'd623: dataIn2 = 32'd0; 
32'd624: dataIn2 = 32'd1; 
32'd625: dataIn2 = 32'd1; 
32'd626: dataIn2 = 32'd0; 
32'd627: dataIn2 = 32'd0; 
32'd628: dataIn2 = 32'd1; 
32'd629: dataIn2 = 32'd0; 
32'd630: dataIn2 = 32'd1; 
32'd631: dataIn2 = 32'd0; 
32'd632: dataIn2 = 32'd1; 
32'd633: dataIn2 = 32'd1; 
32'd634: dataIn2 = 32'd0; 
32'd635: dataIn2 = 32'd1; 
32'd636: dataIn2 = 32'd0; 
32'd637: dataIn2 = 32'd0; 
32'd638: dataIn2 = 32'd0; 
32'd639: dataIn2 = 32'd0; 
32'd640: dataIn2 = 32'd0; 
32'd641: dataIn2 = 32'd0; 
32'd642: dataIn2 = 32'd0; 
32'd643: dataIn2 = 32'd1; 
32'd644: dataIn2 = 32'd0; 
32'd645: dataIn2 = 32'd0; 
32'd646: dataIn2 = 32'd1; 
32'd647: dataIn2 = 32'd0; 
32'd648: dataIn2 = 32'd1; 
32'd649: dataIn2 = 32'd0; 
32'd650: dataIn2 = 32'd0; 
32'd651: dataIn2 = 32'd1; 
32'd652: dataIn2 = 32'd0; 
32'd653: dataIn2 = 32'd0; 
32'd654: dataIn2 = 32'd0; 
32'd655: dataIn2 = 32'd1; 
32'd656: dataIn2 = 32'd0; 
32'd657: dataIn2 = 32'd0; 
32'd658: dataIn2 = 32'd0; 
32'd659: dataIn2 = 32'd0; 
32'd660: dataIn2 = 32'd0; 
32'd661: dataIn2 = 32'd1; 
32'd662: dataIn2 = 32'd0; 
32'd663: dataIn2 = 32'd1; 
32'd664: dataIn2 = 32'd0; 
32'd665: dataIn2 = 32'd0; 
32'd666: dataIn2 = 32'd0; 
32'd667: dataIn2 = 32'd0; 
32'd668: dataIn2 = 32'd0; 
32'd669: dataIn2 = 32'd1; 
32'd670: dataIn2 = 32'd0; 
32'd671: dataIn2 = 32'd0; 
32'd672: dataIn2 = 32'd1; 
32'd673: dataIn2 = 32'd1; 
32'd674: dataIn2 = 32'd1; 
32'd675: dataIn2 = 32'd1; 
32'd676: dataIn2 = 32'd0; 
32'd677: dataIn2 = 32'd1; 
32'd678: dataIn2 = 32'd1; 
32'd679: dataIn2 = 32'd0; 
32'd680: dataIn2 = 32'd0; 
32'd681: dataIn2 = 32'd1; 
32'd682: dataIn2 = 32'd0; 
32'd683: dataIn2 = 32'd1; 
32'd684: dataIn2 = 32'd1; 
32'd685: dataIn2 = 32'd0; 
32'd686: dataIn2 = 32'd1; 
32'd687: dataIn2 = 32'd0; 
32'd688: dataIn2 = 32'd1; 
32'd689: dataIn2 = 32'd1; 
32'd690: dataIn2 = 32'd1; 
32'd691: dataIn2 = 32'd0; 
32'd692: dataIn2 = 32'd0; 
32'd693: dataIn2 = 32'd0; 
32'd694: dataIn2 = 32'd0; 
32'd695: dataIn2 = 32'd0; 
32'd696: dataIn2 = 32'd1; 
32'd697: dataIn2 = 32'd0; 
32'd698: dataIn2 = 32'd1; 
32'd699: dataIn2 = 32'd1; 
32'd700: dataIn2 = 32'd0; 
32'd701: dataIn2 = 32'd0; 
32'd702: dataIn2 = 32'd0; 
32'd703: dataIn2 = 32'd1; 
32'd704: dataIn2 = 32'd0; 
32'd705: dataIn2 = 32'd0; 
32'd706: dataIn2 = 32'd0; 
32'd707: dataIn2 = 32'd0; 
32'd708: dataIn2 = 32'd0; 
32'd709: dataIn2 = 32'd0; 
32'd710: dataIn2 = 32'd1; 
32'd711: dataIn2 = 32'd0; 
32'd712: dataIn2 = 32'd1; 
32'd713: dataIn2 = 32'd1; 
32'd714: dataIn2 = 32'd0; 
32'd715: dataIn2 = 32'd1; 
32'd716: dataIn2 = 32'd1; 
32'd717: dataIn2 = 32'd1; 
32'd718: dataIn2 = 32'd0; 
32'd719: dataIn2 = 32'd1; 
32'd720: dataIn2 = 32'd0; 
32'd721: dataIn2 = 32'd0; 
32'd722: dataIn2 = 32'd0; 
32'd723: dataIn2 = 32'd1; 
32'd724: dataIn2 = 32'd0; 
32'd725: dataIn2 = 32'd1; 
32'd726: dataIn2 = 32'd1; 
32'd727: dataIn2 = 32'd0; 
32'd728: dataIn2 = 32'd0; 
32'd729: dataIn2 = 32'd0; 
32'd730: dataIn2 = 32'd1; 
32'd731: dataIn2 = 32'd0; 
32'd732: dataIn2 = 32'd1; 
32'd733: dataIn2 = 32'd0; 
32'd734: dataIn2 = 32'd1; 
32'd735: dataIn2 = 32'd0; 
32'd736: dataIn2 = 32'd0; 
32'd737: dataIn2 = 32'd1; 
32'd738: dataIn2 = 32'd1; 
32'd739: dataIn2 = 32'd0; 
32'd740: dataIn2 = 32'd1; 
32'd741: dataIn2 = 32'd1; 
32'd742: dataIn2 = 32'd1; 
32'd743: dataIn2 = 32'd1; 
32'd744: dataIn2 = 32'd1; 
32'd745: dataIn2 = 32'd1; 
32'd746: dataIn2 = 32'd1; 
32'd747: dataIn2 = 32'd1; 
32'd748: dataIn2 = 32'd0; 
32'd749: dataIn2 = 32'd0; 
32'd750: dataIn2 = 32'd0; 
32'd751: dataIn2 = 32'd0; 
32'd752: dataIn2 = 32'd0; 
32'd753: dataIn2 = 32'd1; 
32'd754: dataIn2 = 32'd0; 
32'd755: dataIn2 = 32'd1; 
32'd756: dataIn2 = 32'd0; 
32'd757: dataIn2 = 32'd1; 
32'd758: dataIn2 = 32'd0; 
32'd759: dataIn2 = 32'd1; 
32'd760: dataIn2 = 32'd1; 
32'd761: dataIn2 = 32'd0; 
32'd762: dataIn2 = 32'd0; 
32'd763: dataIn2 = 32'd1; 
32'd764: dataIn2 = 32'd0; 
32'd765: dataIn2 = 32'd1; 
32'd766: dataIn2 = 32'd1; 
32'd767: dataIn2 = 32'd0; 
32'd768: dataIn2 = 32'd0; 
32'd769: dataIn2 = 32'd0; 
32'd770: dataIn2 = 32'd0; 
32'd771: dataIn2 = 32'd1; 
32'd772: dataIn2 = 32'd1; 
32'd773: dataIn2 = 32'd0; 
32'd774: dataIn2 = 32'd1; 
32'd775: dataIn2 = 32'd1; 
32'd776: dataIn2 = 32'd0; 
32'd777: dataIn2 = 32'd0; 
32'd778: dataIn2 = 32'd0; 
32'd779: dataIn2 = 32'd0; 
32'd780: dataIn2 = 32'd0; 
32'd781: dataIn2 = 32'd0; 
32'd782: dataIn2 = 32'd0; 
32'd783: dataIn2 = 32'd0; 
32'd784: dataIn2 = 32'd0; 
32'd785: dataIn2 = 32'd0; 
32'd786: dataIn2 = 32'd1; 
32'd787: dataIn2 = 32'd0; 
32'd788: dataIn2 = 32'd0; 
32'd789: dataIn2 = 32'd0; 
32'd790: dataIn2 = 32'd1; 
32'd791: dataIn2 = 32'd1; 
32'd792: dataIn2 = 32'd1; 
32'd793: dataIn2 = 32'd0; 
32'd794: dataIn2 = 32'd1; 
32'd795: dataIn2 = 32'd0; 
32'd796: dataIn2 = 32'd1; 
32'd797: dataIn2 = 32'd1; 
32'd798: dataIn2 = 32'd0; 
32'd799: dataIn2 = 32'd1; 
32'd800: dataIn2 = 32'd0; 
32'd801: dataIn2 = 32'd1; 
32'd802: dataIn2 = 32'd0; 
32'd803: dataIn2 = 32'd1; 
32'd804: dataIn2 = 32'd1; 
32'd805: dataIn2 = 32'd0; 
32'd806: dataIn2 = 32'd0; 
32'd807: dataIn2 = 32'd1; 
32'd808: dataIn2 = 32'd0; 
32'd809: dataIn2 = 32'd0; 
32'd810: dataIn2 = 32'd0; 
32'd811: dataIn2 = 32'd1; 
32'd812: dataIn2 = 32'd1; 
32'd813: dataIn2 = 32'd1; 
32'd814: dataIn2 = 32'd1; 
32'd815: dataIn2 = 32'd0; 
32'd816: dataIn2 = 32'd1; 
32'd817: dataIn2 = 32'd0; 
32'd818: dataIn2 = 32'd0; 
32'd819: dataIn2 = 32'd1; 
32'd820: dataIn2 = 32'd0; 
32'd821: dataIn2 = 32'd1; 
32'd822: dataIn2 = 32'd1; 
32'd823: dataIn2 = 32'd0; 
32'd824: dataIn2 = 32'd1; 
32'd825: dataIn2 = 32'd1; 
32'd826: dataIn2 = 32'd1; 
32'd827: dataIn2 = 32'd0; 
32'd828: dataIn2 = 32'd0; 
32'd829: dataIn2 = 32'd0; 
32'd830: dataIn2 = 32'd0; 
32'd831: dataIn2 = 32'd1; 
32'd832: dataIn2 = 32'd1; 
32'd833: dataIn2 = 32'd0; 
32'd834: dataIn2 = 32'd0; 
32'd835: dataIn2 = 32'd0; 
32'd836: dataIn2 = 32'd1; 
32'd837: dataIn2 = 32'd1; 
32'd838: dataIn2 = 32'd0; 
32'd839: dataIn2 = 32'd0; 
32'd840: dataIn2 = 32'd0; 
32'd841: dataIn2 = 32'd0; 
32'd842: dataIn2 = 32'd1; 
32'd843: dataIn2 = 32'd0; 
32'd844: dataIn2 = 32'd1; 
32'd845: dataIn2 = 32'd0; 
32'd846: dataIn2 = 32'd0; 
32'd847: dataIn2 = 32'd1; 
32'd848: dataIn2 = 32'd1; 
32'd849: dataIn2 = 32'd0; 
32'd850: dataIn2 = 32'd1; 
32'd851: dataIn2 = 32'd1; 
32'd852: dataIn2 = 32'd1; 
32'd853: dataIn2 = 32'd1; 
32'd854: dataIn2 = 32'd1; 
32'd855: dataIn2 = 32'd1; 
32'd856: dataIn2 = 32'd0; 
32'd857: dataIn2 = 32'd0; 
32'd858: dataIn2 = 32'd1; 
32'd859: dataIn2 = 32'd0; 
32'd860: dataIn2 = 32'd1; 
32'd861: dataIn2 = 32'd0; 
32'd862: dataIn2 = 32'd1; 
32'd863: dataIn2 = 32'd0; 
32'd864: dataIn2 = 32'd0; 
32'd865: dataIn2 = 32'd1; 
32'd866: dataIn2 = 32'd0; 
32'd867: dataIn2 = 32'd1; 
32'd868: dataIn2 = 32'd0; 
32'd869: dataIn2 = 32'd1; 
32'd870: dataIn2 = 32'd0; 
32'd871: dataIn2 = 32'd0; 
32'd872: dataIn2 = 32'd0; 
32'd873: dataIn2 = 32'd0; 
32'd874: dataIn2 = 32'd0; 
32'd875: dataIn2 = 32'd0; 
32'd876: dataIn2 = 32'd0; 
32'd877: dataIn2 = 32'd1; 
32'd878: dataIn2 = 32'd0; 
32'd879: dataIn2 = 32'd0; 
32'd880: dataIn2 = 32'd0; 
32'd881: dataIn2 = 32'd1; 
32'd882: dataIn2 = 32'd0; 
32'd883: dataIn2 = 32'd0; 
32'd884: dataIn2 = 32'd0; 
32'd885: dataIn2 = 32'd0; 
32'd886: dataIn2 = 32'd0; 
32'd887: dataIn2 = 32'd1; 
32'd888: dataIn2 = 32'd1; 
32'd889: dataIn2 = 32'd0; 
32'd890: dataIn2 = 32'd1; 
32'd891: dataIn2 = 32'd1; 
32'd892: dataIn2 = 32'd1; 
32'd893: dataIn2 = 32'd0; 
32'd894: dataIn2 = 32'd0; 
32'd895: dataIn2 = 32'd1; 
32'd896: dataIn2 = 32'd0; 
32'd897: dataIn2 = 32'd0; 
32'd898: dataIn2 = 32'd1; 
32'd899: dataIn2 = 32'd1; 
32'd900: dataIn2 = 32'd0; 
32'd901: dataIn2 = 32'd1; 
32'd902: dataIn2 = 32'd1; 
32'd903: dataIn2 = 32'd1; 
32'd904: dataIn2 = 32'd1; 
32'd905: dataIn2 = 32'd1; 
32'd906: dataIn2 = 32'd1; 
32'd907: dataIn2 = 32'd1; 
32'd908: dataIn2 = 32'd0; 
32'd909: dataIn2 = 32'd0; 
32'd910: dataIn2 = 32'd0; 
32'd911: dataIn2 = 32'd1; 
32'd912: dataIn2 = 32'd1; 
32'd913: dataIn2 = 32'd0; 
32'd914: dataIn2 = 32'd1; 
32'd915: dataIn2 = 32'd0; 
32'd916: dataIn2 = 32'd0; 
32'd917: dataIn2 = 32'd1; 
32'd918: dataIn2 = 32'd0; 
32'd919: dataIn2 = 32'd0; 
32'd920: dataIn2 = 32'd1; 
32'd921: dataIn2 = 32'd1; 
32'd922: dataIn2 = 32'd1; 
32'd923: dataIn2 = 32'd0; 
32'd924: dataIn2 = 32'd0; 
32'd925: dataIn2 = 32'd1; 
32'd926: dataIn2 = 32'd0; 
32'd927: dataIn2 = 32'd1; 
32'd928: dataIn2 = 32'd0; 
32'd929: dataIn2 = 32'd1; 
32'd930: dataIn2 = 32'd1; 
32'd931: dataIn2 = 32'd0; 
32'd932: dataIn2 = 32'd1; 
32'd933: dataIn2 = 32'd0; 
32'd934: dataIn2 = 32'd1; 
32'd935: dataIn2 = 32'd0; 
32'd936: dataIn2 = 32'd0; 
32'd937: dataIn2 = 32'd0; 
32'd938: dataIn2 = 32'd1; 
32'd939: dataIn2 = 32'd1; 
32'd940: dataIn2 = 32'd0; 
32'd941: dataIn2 = 32'd0; 
32'd942: dataIn2 = 32'd0; 
32'd943: dataIn2 = 32'd1; 
32'd944: dataIn2 = 32'd0; 
32'd945: dataIn2 = 32'd0; 
32'd946: dataIn2 = 32'd0; 
32'd947: dataIn2 = 32'd1; 
32'd948: dataIn2 = 32'd0; 
32'd949: dataIn2 = 32'd1; 
32'd950: dataIn2 = 32'd0; 
32'd951: dataIn2 = 32'd0; 
32'd952: dataIn2 = 32'd1; 
32'd953: dataIn2 = 32'd0; 
32'd954: dataIn2 = 32'd1; 
32'd955: dataIn2 = 32'd1; 
32'd956: dataIn2 = 32'd1; 
32'd957: dataIn2 = 32'd0; 
32'd958: dataIn2 = 32'd1; 
32'd959: dataIn2 = 32'd0; 
32'd960: dataIn2 = 32'd0; 
32'd961: dataIn2 = 32'd1; 
32'd962: dataIn2 = 32'd1; 
32'd963: dataIn2 = 32'd1; 
32'd964: dataIn2 = 32'd0; 
32'd965: dataIn2 = 32'd0; 
32'd966: dataIn2 = 32'd0; 
32'd967: dataIn2 = 32'd0; 
32'd968: dataIn2 = 32'd0; 
32'd969: dataIn2 = 32'd1; 
32'd970: dataIn2 = 32'd1; 
32'd971: dataIn2 = 32'd0; 
32'd972: dataIn2 = 32'd1; 
32'd973: dataIn2 = 32'd1; 
32'd974: dataIn2 = 32'd1; 
32'd975: dataIn2 = 32'd1; 
32'd976: dataIn2 = 32'd0; 
32'd977: dataIn2 = 32'd0; 
32'd978: dataIn2 = 32'd0; 
32'd979: dataIn2 = 32'd1; 
32'd980: dataIn2 = 32'd1; 
32'd981: dataIn2 = 32'd1; 
32'd982: dataIn2 = 32'd0; 
32'd983: dataIn2 = 32'd1; 
32'd984: dataIn2 = 32'd1; 
32'd985: dataIn2 = 32'd0; 
32'd986: dataIn2 = 32'd1; 
32'd987: dataIn2 = 32'd0; 
32'd988: dataIn2 = 32'd0; 
32'd989: dataIn2 = 32'd1; 
32'd990: dataIn2 = 32'd1; 
32'd991: dataIn2 = 32'd0; 
32'd992: dataIn2 = 32'd1; 
default: 
	dataIn2 = 32'd99999; 
endcase 
end 
always begin 
#10 Clk = ~Clk; 
end 
//========== VCD ============ 
`ifdef VCD 
initial 
begin 
	$dumpfile("jpwh.vcd");  
	$dumpvars; 
end 
`endif 
//===========RTLVCD ========== 
`ifdef RTLVCD 
initial 
begin 
	$dumpfile("hht_rtl.vcd"); 
	$dumpvars; 
end 
`endif 
endmodule 
