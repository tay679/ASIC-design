//11738x11738 
// Code your testbench here 
// or browse Examples 
// Verilog test bench for HHT with buffer 
`timescale 1ns/1ps 
module testbench; 
  parameter V_SIZE = 9; 
  parameter COL_SIZE = 79566 ; 
reg Clk,Rst,WR,mem_init; 
reg [31:0] dataIn1,dataIn2,csize; 
reg [31:0]v_values_base; 
wire [31:0]addr1,addr2; 
wire [4:0] regaddr1,regaddr2; 
reg[31:0] cpu_addr;
wire hht;
wire [31:0]val[0:8]; 
reg [31:0]wdata_col_base; 
wire [31:0] dataOut; 
reg fe_init; 
reg wn,rn,RD; 
wire [4:0]adata; 
wire [31:0] rdata; 
 // Instantiate memory module 
//  memmodel m1 (addr,dataIn,dataOut,WR,Clk,Rst); 
//  mem_buffer m1 (dataOut, full, empty, Clk, Rst, wn, rn, dataIn); 
control t1 (Clk,wdata_col_base,v_values_base,addr1,addr2,dataIn1,dataIn2,Rst,RD,csize,cpu_addr,hht,regaddr1,regaddr2,rdata,adata); ;  
//frontend t1 (Clk,Rst,fe_init,wdata_col_base,data_req,dataIn,init, 
//{m_cols[0],m_cols[1],m_cols[2],m_cols[3],m_cols[4]}, 
//done,wn); 
initial begin 
Clk = 1'b0; 
  RD = 1'b1; 
 #15; 
Rst = 1'b0; 
cpu_addr = 32'd126;
  v_values_base = 32'd2; 
  wdata_col_base = 32'd117400 ; 
  csize = COL_SIZE; 
 fe_init = 1'b1; 
#15 Rst = 1'b1; 
// RD = 1'b0; 
// RD = 1'b1; 
 #17100000; 
$finish; 
end 
always @(*) begin 
//$display("%b,%b",t1.fe1.count,t1.fe1.vdata_req); 
case(addr1)  
32'd117400: dataIn1 = 32'd1
; 
32'd117401: dataIn1 = 32'd959
; 
32'd117402: dataIn1 = 32'd1264
; 
32'd117403: dataIn1 = 32'd1265
; 
32'd117404: dataIn1 = 32'd1267
; 
32'd117405: dataIn1 = 32'd1469
; 
32'd117406: dataIn1 = 32'd1859
; 
32'd117407: dataIn1 = 32'd2
; 
32'd117408: dataIn1 = 32'd3426
; 
32'd117409: dataIn1 = 32'd3427
; 
32'd117410: dataIn1 = 32'd3452
; 
32'd117411: dataIn1 = 32'd3453
; 
32'd117412: dataIn1 = 32'd3483
; 
32'd117413: dataIn1 = 32'd3487
; 
32'd117414: dataIn1 = 32'd3
; 
32'd117415: dataIn1 = 32'd4636
; 
32'd117416: dataIn1 = 32'd4638
; 
32'd117417: dataIn1 = 32'd9689
; 
32'd117418: dataIn1 = 32'd9690
; 
32'd117419: dataIn1 = 32'd9757
; 
32'd117420: dataIn1 = 32'd4
; 
32'd117421: dataIn1 = 32'd4644
; 
32'd117422: dataIn1 = 32'd4646
; 
32'd117423: dataIn1 = 32'd4817
; 
32'd117424: dataIn1 = 32'd4836
; 
32'd117425: dataIn1 = 32'd5861
; 
32'd117426: dataIn1 = 32'd6140
; 
32'd117427: dataIn1 = 32'd8902
; 
32'd117428: dataIn1 = 32'd5
; 
32'd117429: dataIn1 = 32'd5740
; 
32'd117430: dataIn1 = 32'd5741
; 
32'd117431: dataIn1 = 32'd5826
; 
32'd117432: dataIn1 = 32'd6055
; 
32'd117433: dataIn1 = 32'd8924
; 
32'd117434: dataIn1 = 32'd8925
; 
32'd117435: dataIn1 = 32'd6
; 
32'd117436: dataIn1 = 32'd5938
; 
32'd117437: dataIn1 = 32'd5940
; 
32'd117438: dataIn1 = 32'd5995
; 
32'd117439: dataIn1 = 32'd6065
; 
32'd117440: dataIn1 = 32'd8962
; 
32'd117441: dataIn1 = 32'd8963
; 
32'd117442: dataIn1 = 32'd7
; 
32'd117443: dataIn1 = 32'd7605
; 
32'd117444: dataIn1 = 32'd7606
; 
32'd117445: dataIn1 = 32'd7712
; 
32'd117446: dataIn1 = 32'd7713
; 
32'd117447: dataIn1 = 32'd9605
; 
32'd117448: dataIn1 = 32'd9607
; 
32'd117449: dataIn1 = 32'd8
; 
32'd117450: dataIn1 = 32'd4716
; 
32'd117451: dataIn1 = 32'd4717
; 
32'd117452: dataIn1 = 32'd7858
; 
32'd117453: dataIn1 = 32'd7859
; 
32'd117454: dataIn1 = 32'd7965
; 
32'd117455: dataIn1 = 32'd7966
; 
32'd117456: dataIn1 = 32'd9
; 
32'd117457: dataIn1 = 32'd4734
; 
32'd117458: dataIn1 = 32'd4735
; 
32'd117459: dataIn1 = 32'd8111
; 
32'd117460: dataIn1 = 32'd8112
; 
32'd117461: dataIn1 = 32'd8218
; 
32'd117462: dataIn1 = 32'd8219
; 
32'd117463: dataIn1 = 32'd10
; 
32'd117464: dataIn1 = 32'd4752
; 
32'd117465: dataIn1 = 32'd4753
; 
32'd117466: dataIn1 = 32'd8363
; 
32'd117467: dataIn1 = 32'd8364
; 
32'd117468: dataIn1 = 32'd8470
; 
32'd117469: dataIn1 = 32'd8471
; 
32'd117470: dataIn1 = 32'd11
; 
32'd117471: dataIn1 = 32'd4770
; 
32'd117472: dataIn1 = 32'd4771
; 
32'd117473: dataIn1 = 32'd8616
; 
32'd117474: dataIn1 = 32'd8617
; 
32'd117475: dataIn1 = 32'd8723
; 
32'd117476: dataIn1 = 32'd8724
; 
32'd117477: dataIn1 = 32'd12
; 
32'd117478: dataIn1 = 32'd4788
; 
32'd117479: dataIn1 = 32'd4789
; 
32'd117480: dataIn1 = 32'd8868
; 
32'd117481: dataIn1 = 32'd8869
; 
32'd117482: dataIn1 = 32'd9448
; 
32'd117483: dataIn1 = 32'd13
; 
32'd117484: dataIn1 = 32'd3467
; 
32'd117485: dataIn1 = 32'd9313
; 
32'd117486: dataIn1 = 32'd9314
; 
32'd117487: dataIn1 = 32'd14
; 
32'd117488: dataIn1 = 32'd3434
; 
32'd117489: dataIn1 = 32'd3457
; 
32'd117490: dataIn1 = 32'd5431
; 
32'd117491: dataIn1 = 32'd5432
; 
32'd117492: dataIn1 = 32'd5513
; 
32'd117493: dataIn1 = 32'd6730
; 
32'd117494: dataIn1 = 32'd6734
; 
32'd117495: dataIn1 = 32'd15
; 
32'd117496: dataIn1 = 32'd2323
; 
32'd117497: dataIn1 = 32'd2324
; 
32'd117498: dataIn1 = 32'd2737
; 
32'd117499: dataIn1 = 32'd2741
; 
32'd117500: dataIn1 = 32'd3433
; 
32'd117501: dataIn1 = 32'd3436
; 
32'd117502: dataIn1 = 32'd3978
; 
32'd117503: dataIn1 = 32'd16
; 
32'd117504: dataIn1 = 32'd2701
; 
32'd117505: dataIn1 = 32'd2702
; 
32'd117506: dataIn1 = 32'd2742
; 
32'd117507: dataIn1 = 32'd2746
; 
32'd117508: dataIn1 = 32'd3435
; 
32'd117509: dataIn1 = 32'd3437
; 
32'd117510: dataIn1 = 32'd17
; 
32'd117511: dataIn1 = 32'd2748
; 
32'd117512: dataIn1 = 32'd3419
; 
32'd117513: dataIn1 = 32'd5433
; 
32'd117514: dataIn1 = 32'd5434
; 
32'd117515: dataIn1 = 32'd5514
; 
32'd117516: dataIn1 = 32'd5515
; 
32'd117517: dataIn1 = 32'd9328
; 
32'd117518: dataIn1 = 32'd18
; 
32'd117519: dataIn1 = 32'd2107
; 
32'd117520: dataIn1 = 32'd2108
; 
32'd117521: dataIn1 = 32'd5435
; 
32'd117522: dataIn1 = 32'd5436
; 
32'd117523: dataIn1 = 32'd5516
; 
32'd117524: dataIn1 = 32'd5517
; 
32'd117525: dataIn1 = 32'd9330
; 
32'd117526: dataIn1 = 32'd19
; 
32'd117527: dataIn1 = 32'd2109
; 
32'd117528: dataIn1 = 32'd2111
; 
32'd117529: dataIn1 = 32'd5437
; 
32'd117530: dataIn1 = 32'd5438
; 
32'd117531: dataIn1 = 32'd5518
; 
32'd117532: dataIn1 = 32'd5519
; 
32'd117533: dataIn1 = 32'd6736
; 
32'd117534: dataIn1 = 32'd20
; 
32'd117535: dataIn1 = 32'd5521
; 
32'd117536: dataIn1 = 32'd9452
; 
32'd117537: dataIn1 = 32'd9674
; 
32'd117538: dataIn1 = 32'd9675
; 
32'd117539: dataIn1 = 32'd9755
; 
32'd117540: dataIn1 = 32'd9825
; 
32'd117541: dataIn1 = 32'd10129
; 
32'd117542: dataIn1 = 32'd21
; 
32'd117543: dataIn1 = 32'd2117
; 
32'd117544: dataIn1 = 32'd5441
; 
32'd117545: dataIn1 = 32'd5442
; 
32'd117546: dataIn1 = 32'd5522
; 
32'd117547: dataIn1 = 32'd5523
; 
32'd117548: dataIn1 = 32'd9333
; 
32'd117549: dataIn1 = 32'd10225
; 
32'd117550: dataIn1 = 32'd22
; 
32'd117551: dataIn1 = 32'd2118
; 
32'd117552: dataIn1 = 32'd2120
; 
32'd117553: dataIn1 = 32'd5443
; 
32'd117554: dataIn1 = 32'd5444
; 
32'd117555: dataIn1 = 32'd5524
; 
32'd117556: dataIn1 = 32'd6731
; 
32'd117557: dataIn1 = 32'd9335
; 
32'd117558: dataIn1 = 32'd23
; 
32'd117559: dataIn1 = 32'd2121
; 
32'd117560: dataIn1 = 32'd9316
; 
32'd117561: dataIn1 = 32'd9317
; 
32'd117562: dataIn1 = 32'd24
; 
32'd117563: dataIn1 = 32'd2123
; 
32'd117564: dataIn1 = 32'd2124
; 
32'd117565: dataIn1 = 32'd2126
; 
32'd117566: dataIn1 = 32'd3457
; 
32'd117567: dataIn1 = 32'd3467
; 
32'd117568: dataIn1 = 32'd25
; 
32'd117569: dataIn1 = 32'd2125
; 
32'd117570: dataIn1 = 32'd2126
; 
32'd117571: dataIn1 = 32'd2128
; 
32'd117572: dataIn1 = 32'd2130
; 
32'd117573: dataIn1 = 32'd3433
; 
32'd117574: dataIn1 = 32'd3434
; 
32'd117575: dataIn1 = 32'd26
; 
32'd117576: dataIn1 = 32'd2129
; 
32'd117577: dataIn1 = 32'd2130
; 
32'd117578: dataIn1 = 32'd2132
; 
32'd117579: dataIn1 = 32'd2134
; 
32'd117580: dataIn1 = 32'd3435
; 
32'd117581: dataIn1 = 32'd3436
; 
32'd117582: dataIn1 = 32'd27
; 
32'd117583: dataIn1 = 32'd2133
; 
32'd117584: dataIn1 = 32'd2134
; 
32'd117585: dataIn1 = 32'd2136
; 
32'd117586: dataIn1 = 32'd2138
; 
32'd117587: dataIn1 = 32'd3419
; 
32'd117588: dataIn1 = 32'd3437
; 
32'd117589: dataIn1 = 32'd28
; 
32'd117590: dataIn1 = 32'd2106
; 
32'd117591: dataIn1 = 32'd2108
; 
32'd117592: dataIn1 = 32'd2137
; 
32'd117593: dataIn1 = 32'd2138
; 
32'd117594: dataIn1 = 32'd2140
; 
32'd117595: dataIn1 = 32'd2748
; 
32'd117596: dataIn1 = 32'd29
; 
32'd117597: dataIn1 = 32'd2106
; 
32'd117598: dataIn1 = 32'd2107
; 
32'd117599: dataIn1 = 32'd2109
; 
32'd117600: dataIn1 = 32'd2110
; 
32'd117601: dataIn1 = 32'd2141
; 
32'd117602: dataIn1 = 32'd2143
; 
32'd117603: dataIn1 = 32'd30
; 
32'd117604: dataIn1 = 32'd2110
; 
32'd117605: dataIn1 = 32'd2111
; 
32'd117606: dataIn1 = 32'd2112
; 
32'd117607: dataIn1 = 32'd2113
; 
32'd117608: dataIn1 = 32'd2144
; 
32'd117609: dataIn1 = 32'd2146
; 
32'd117610: dataIn1 = 32'd9450
; 
32'd117611: dataIn1 = 32'd10155
; 
32'd117612: dataIn1 = 32'd31
; 
32'd117613: dataIn1 = 32'd2116
; 
32'd117614: dataIn1 = 32'd9454
; 
32'd117615: dataIn1 = 32'd9455
; 
32'd117616: dataIn1 = 32'd9457
; 
32'd117617: dataIn1 = 32'd9462
; 
32'd117618: dataIn1 = 32'd9818
; 
32'd117619: dataIn1 = 32'd9829
; 
32'd117620: dataIn1 = 32'd10153
; 
32'd117621: dataIn1 = 32'd32
; 
32'd117622: dataIn1 = 32'd2116
; 
32'd117623: dataIn1 = 32'd2117
; 
32'd117624: dataIn1 = 32'd2118
; 
32'd117625: dataIn1 = 32'd2119
; 
32'd117626: dataIn1 = 32'd2150
; 
32'd117627: dataIn1 = 32'd2152
; 
32'd117628: dataIn1 = 32'd33
; 
32'd117629: dataIn1 = 32'd2119
; 
32'd117630: dataIn1 = 32'd2120
; 
32'd117631: dataIn1 = 32'd2121
; 
32'd117632: dataIn1 = 32'd2153
; 
32'd117633: dataIn1 = 32'd2155
; 
32'd117634: dataIn1 = 32'd34
; 
32'd117635: dataIn1 = 32'd2122
; 
32'd117636: dataIn1 = 32'd2124
; 
32'd117637: dataIn1 = 32'd2157
; 
32'd117638: dataIn1 = 32'd35
; 
32'd117639: dataIn1 = 32'd2122
; 
32'd117640: dataIn1 = 32'd2123
; 
32'd117641: dataIn1 = 32'd2125
; 
32'd117642: dataIn1 = 32'd2127
; 
32'd117643: dataIn1 = 32'd2156
; 
32'd117644: dataIn1 = 32'd2159
; 
32'd117645: dataIn1 = 32'd36
; 
32'd117646: dataIn1 = 32'd2127
; 
32'd117647: dataIn1 = 32'd2128
; 
32'd117648: dataIn1 = 32'd2129
; 
32'd117649: dataIn1 = 32'd2131
; 
32'd117650: dataIn1 = 32'd2160
; 
32'd117651: dataIn1 = 32'd2162
; 
32'd117652: dataIn1 = 32'd37
; 
32'd117653: dataIn1 = 32'd2131
; 
32'd117654: dataIn1 = 32'd2132
; 
32'd117655: dataIn1 = 32'd2133
; 
32'd117656: dataIn1 = 32'd2135
; 
32'd117657: dataIn1 = 32'd2163
; 
32'd117658: dataIn1 = 32'd2165
; 
32'd117659: dataIn1 = 32'd38
; 
32'd117660: dataIn1 = 32'd2135
; 
32'd117661: dataIn1 = 32'd2136
; 
32'd117662: dataIn1 = 32'd2137
; 
32'd117663: dataIn1 = 32'd2139
; 
32'd117664: dataIn1 = 32'd2166
; 
32'd117665: dataIn1 = 32'd2168
; 
32'd117666: dataIn1 = 32'd39
; 
32'd117667: dataIn1 = 32'd2139
; 
32'd117668: dataIn1 = 32'd2140
; 
32'd117669: dataIn1 = 32'd2141
; 
32'd117670: dataIn1 = 32'd2142
; 
32'd117671: dataIn1 = 32'd2169
; 
32'd117672: dataIn1 = 32'd2171
; 
32'd117673: dataIn1 = 32'd40
; 
32'd117674: dataIn1 = 32'd2142
; 
32'd117675: dataIn1 = 32'd2143
; 
32'd117676: dataIn1 = 32'd2144
; 
32'd117677: dataIn1 = 32'd2145
; 
32'd117678: dataIn1 = 32'd2172
; 
32'd117679: dataIn1 = 32'd2174
; 
32'd117680: dataIn1 = 32'd41
; 
32'd117681: dataIn1 = 32'd2145
; 
32'd117682: dataIn1 = 32'd9463
; 
32'd117683: dataIn1 = 32'd9464
; 
32'd117684: dataIn1 = 32'd9467
; 
32'd117685: dataIn1 = 32'd9781
; 
32'd117686: dataIn1 = 32'd9838
; 
32'd117687: dataIn1 = 32'd9845
; 
32'd117688: dataIn1 = 32'd10157
; 
32'd117689: dataIn1 = 32'd42
; 
32'd117690: dataIn1 = 32'd2150
; 
32'd117691: dataIn1 = 32'd3595
; 
32'd117692: dataIn1 = 32'd3596
; 
32'd117693: dataIn1 = 32'd3603
; 
32'd117694: dataIn1 = 32'd9477
; 
32'd117695: dataIn1 = 32'd9769
; 
32'd117696: dataIn1 = 32'd43
; 
32'd117697: dataIn1 = 32'd2152
; 
32'd117698: dataIn1 = 32'd2153
; 
32'd117699: dataIn1 = 32'd2154
; 
32'd117700: dataIn1 = 32'd3605
; 
32'd117701: dataIn1 = 32'd3606
; 
32'd117702: dataIn1 = 32'd5308
; 
32'd117703: dataIn1 = 32'd44
; 
32'd117704: dataIn1 = 32'd2154
; 
32'd117705: dataIn1 = 32'd2155
; 
32'd117706: dataIn1 = 32'd2184
; 
32'd117707: dataIn1 = 32'd45
; 
32'd117708: dataIn1 = 32'd2156
; 
32'd117709: dataIn1 = 32'd2157
; 
32'd117710: dataIn1 = 32'd2158
; 
32'd117711: dataIn1 = 32'd2186
; 
32'd117712: dataIn1 = 32'd2187
; 
32'd117713: dataIn1 = 32'd46
; 
32'd117714: dataIn1 = 32'd2158
; 
32'd117715: dataIn1 = 32'd2159
; 
32'd117716: dataIn1 = 32'd2160
; 
32'd117717: dataIn1 = 32'd2161
; 
32'd117718: dataIn1 = 32'd2188
; 
32'd117719: dataIn1 = 32'd2190
; 
32'd117720: dataIn1 = 32'd47
; 
32'd117721: dataIn1 = 32'd2161
; 
32'd117722: dataIn1 = 32'd2162
; 
32'd117723: dataIn1 = 32'd2163
; 
32'd117724: dataIn1 = 32'd2164
; 
32'd117725: dataIn1 = 32'd2191
; 
32'd117726: dataIn1 = 32'd2193
; 
32'd117727: dataIn1 = 32'd48
; 
32'd117728: dataIn1 = 32'd2164
; 
32'd117729: dataIn1 = 32'd2165
; 
32'd117730: dataIn1 = 32'd2166
; 
32'd117731: dataIn1 = 32'd2167
; 
32'd117732: dataIn1 = 32'd2194
; 
32'd117733: dataIn1 = 32'd2196
; 
32'd117734: dataIn1 = 32'd49
; 
32'd117735: dataIn1 = 32'd2167
; 
32'd117736: dataIn1 = 32'd2168
; 
32'd117737: dataIn1 = 32'd2169
; 
32'd117738: dataIn1 = 32'd2170
; 
32'd117739: dataIn1 = 32'd2197
; 
32'd117740: dataIn1 = 32'd2199
; 
32'd117741: dataIn1 = 32'd50
; 
32'd117742: dataIn1 = 32'd2170
; 
32'd117743: dataIn1 = 32'd2171
; 
32'd117744: dataIn1 = 32'd2172
; 
32'd117745: dataIn1 = 32'd2173
; 
32'd117746: dataIn1 = 32'd2200
; 
32'd117747: dataIn1 = 32'd2202
; 
32'd117748: dataIn1 = 32'd3611
; 
32'd117749: dataIn1 = 32'd51
; 
32'd117750: dataIn1 = 32'd2173
; 
32'd117751: dataIn1 = 32'd2174
; 
32'd117752: dataIn1 = 32'd3623
; 
32'd117753: dataIn1 = 32'd3624
; 
32'd117754: dataIn1 = 32'd3631
; 
32'd117755: dataIn1 = 32'd9780
; 
32'd117756: dataIn1 = 32'd52
; 
32'd117757: dataIn1 = 32'd3591
; 
32'd117758: dataIn1 = 32'd3597
; 
32'd117759: dataIn1 = 32'd3637
; 
32'd117760: dataIn1 = 32'd10158
; 
32'd117761: dataIn1 = 32'd10159
; 
32'd117762: dataIn1 = 32'd10226
; 
32'd117763: dataIn1 = 32'd53
; 
32'd117764: dataIn1 = 32'd3598
; 
32'd117765: dataIn1 = 32'd3599
; 
32'd117766: dataIn1 = 32'd3604
; 
32'd117767: dataIn1 = 32'd3610
; 
32'd117768: dataIn1 = 32'd3645
; 
32'd117769: dataIn1 = 32'd3649
; 
32'd117770: dataIn1 = 32'd54
; 
32'd117771: dataIn1 = 32'd2182
; 
32'd117772: dataIn1 = 32'd2183
; 
32'd117773: dataIn1 = 32'd2184
; 
32'd117774: dataIn1 = 32'd2212
; 
32'd117775: dataIn1 = 32'd2214
; 
32'd117776: dataIn1 = 32'd3609
; 
32'd117777: dataIn1 = 32'd5309
; 
32'd117778: dataIn1 = 32'd55
; 
32'd117779: dataIn1 = 32'd2185
; 
32'd117780: dataIn1 = 32'd2187
; 
32'd117781: dataIn1 = 32'd2216
; 
32'd117782: dataIn1 = 32'd3657
; 
32'd117783: dataIn1 = 32'd56
; 
32'd117784: dataIn1 = 32'd2185
; 
32'd117785: dataIn1 = 32'd2186
; 
32'd117786: dataIn1 = 32'd2188
; 
32'd117787: dataIn1 = 32'd2189
; 
32'd117788: dataIn1 = 32'd2215
; 
32'd117789: dataIn1 = 32'd2218
; 
32'd117790: dataIn1 = 32'd9782
; 
32'd117791: dataIn1 = 32'd57
; 
32'd117792: dataIn1 = 32'd2189
; 
32'd117793: dataIn1 = 32'd2190
; 
32'd117794: dataIn1 = 32'd2191
; 
32'd117795: dataIn1 = 32'd2192
; 
32'd117796: dataIn1 = 32'd2219
; 
32'd117797: dataIn1 = 32'd2221
; 
32'd117798: dataIn1 = 32'd9784
; 
32'd117799: dataIn1 = 32'd58
; 
32'd117800: dataIn1 = 32'd2192
; 
32'd117801: dataIn1 = 32'd2193
; 
32'd117802: dataIn1 = 32'd2194
; 
32'd117803: dataIn1 = 32'd2195
; 
32'd117804: dataIn1 = 32'd2222
; 
32'd117805: dataIn1 = 32'd2224
; 
32'd117806: dataIn1 = 32'd3664
; 
32'd117807: dataIn1 = 32'd59
; 
32'd117808: dataIn1 = 32'd2195
; 
32'd117809: dataIn1 = 32'd2196
; 
32'd117810: dataIn1 = 32'd2197
; 
32'd117811: dataIn1 = 32'd3675
; 
32'd117812: dataIn1 = 32'd3676
; 
32'd117813: dataIn1 = 32'd3683
; 
32'd117814: dataIn1 = 32'd60
; 
32'd117815: dataIn1 = 32'd2199
; 
32'd117816: dataIn1 = 32'd3614
; 
32'd117817: dataIn1 = 32'd3615
; 
32'd117818: dataIn1 = 32'd3685
; 
32'd117819: dataIn1 = 32'd3686
; 
32'd117820: dataIn1 = 32'd3690
; 
32'd117821: dataIn1 = 32'd61
; 
32'd117822: dataIn1 = 32'd3616
; 
32'd117823: dataIn1 = 32'd9549
; 
32'd117824: dataIn1 = 32'd9550
; 
32'd117825: dataIn1 = 32'd9552
; 
32'd117826: dataIn1 = 32'd9556
; 
32'd117827: dataIn1 = 32'd10012
; 
32'd117828: dataIn1 = 32'd10021
; 
32'd117829: dataIn1 = 32'd10196
; 
32'd117830: dataIn1 = 32'd62
; 
32'd117831: dataIn1 = 32'd3626
; 
32'd117832: dataIn1 = 32'd3627
; 
32'd117833: dataIn1 = 32'd3632
; 
32'd117834: dataIn1 = 32'd3638
; 
32'd117835: dataIn1 = 32'd3710
; 
32'd117836: dataIn1 = 32'd3714
; 
32'd117837: dataIn1 = 32'd10166
; 
32'd117838: dataIn1 = 32'd63
; 
32'd117839: dataIn1 = 32'd3639
; 
32'd117840: dataIn1 = 32'd3640
; 
32'd117841: dataIn1 = 32'd3644
; 
32'd117842: dataIn1 = 32'd3650
; 
32'd117843: dataIn1 = 32'd3722
; 
32'd117844: dataIn1 = 32'd3726
; 
32'd117845: dataIn1 = 32'd64
; 
32'd117846: dataIn1 = 32'd2213
; 
32'd117847: dataIn1 = 32'd3651
; 
32'd117848: dataIn1 = 32'd3652
; 
32'd117849: dataIn1 = 32'd3655
; 
32'd117850: dataIn1 = 32'd3731
; 
32'd117851: dataIn1 = 32'd5312
; 
32'd117852: dataIn1 = 32'd65
; 
32'd117853: dataIn1 = 32'd2213
; 
32'd117854: dataIn1 = 32'd2214
; 
32'd117855: dataIn1 = 32'd5455
; 
32'd117856: dataIn1 = 32'd66
; 
32'd117857: dataIn1 = 32'd3656
; 
32'd117858: dataIn1 = 32'd3658
; 
32'd117859: dataIn1 = 32'd9559
; 
32'd117860: dataIn1 = 32'd9560
; 
32'd117861: dataIn1 = 32'd9567
; 
32'd117862: dataIn1 = 32'd10027
; 
32'd117863: dataIn1 = 32'd67
; 
32'd117864: dataIn1 = 32'd10062
; 
32'd117865: dataIn1 = 32'd10063
; 
32'd117866: dataIn1 = 32'd10065
; 
32'd117867: dataIn1 = 32'd10075
; 
32'd117868: dataIn1 = 32'd10205
; 
32'd117869: dataIn1 = 32'd10208
; 
32'd117870: dataIn1 = 32'd68
; 
32'd117871: dataIn1 = 32'd10094
; 
32'd117872: dataIn1 = 32'd10095
; 
32'd117873: dataIn1 = 32'd10097
; 
32'd117874: dataIn1 = 32'd10107
; 
32'd117875: dataIn1 = 32'd10213
; 
32'd117876: dataIn1 = 32'd10216
; 
32'd117877: dataIn1 = 32'd69
; 
32'd117878: dataIn1 = 32'd9920
; 
32'd117879: dataIn1 = 32'd9921
; 
32'd117880: dataIn1 = 32'd9923
; 
32'd117881: dataIn1 = 32'd9942
; 
32'd117882: dataIn1 = 32'd10173
; 
32'd117883: dataIn1 = 32'd10180
; 
32'd117884: dataIn1 = 32'd70
; 
32'd117885: dataIn1 = 32'd3784
; 
32'd117886: dataIn1 = 32'd3788
; 
32'd117887: dataIn1 = 32'd9519
; 
32'd117888: dataIn1 = 32'd9520
; 
32'd117889: dataIn1 = 32'd9526
; 
32'd117890: dataIn1 = 32'd9960
; 
32'd117891: dataIn1 = 32'd10183
; 
32'd117892: dataIn1 = 32'd71
; 
32'd117893: dataIn1 = 32'd3692
; 
32'd117894: dataIn1 = 32'd3693
; 
32'd117895: dataIn1 = 32'd3697
; 
32'd117896: dataIn1 = 32'd3703
; 
32'd117897: dataIn1 = 32'd3796
; 
32'd117898: dataIn1 = 32'd3800
; 
32'd117899: dataIn1 = 32'd10235
; 
32'd117900: dataIn1 = 32'd72
; 
32'd117901: dataIn1 = 32'd3704
; 
32'd117902: dataIn1 = 32'd3705
; 
32'd117903: dataIn1 = 32'd3709
; 
32'd117904: dataIn1 = 32'd3715
; 
32'd117905: dataIn1 = 32'd3808
; 
32'd117906: dataIn1 = 32'd3812
; 
32'd117907: dataIn1 = 32'd73
; 
32'd117908: dataIn1 = 32'd2264
; 
32'd117909: dataIn1 = 32'd3716
; 
32'd117910: dataIn1 = 32'd3717
; 
32'd117911: dataIn1 = 32'd3721
; 
32'd117912: dataIn1 = 32'd3727
; 
32'd117913: dataIn1 = 32'd3820
; 
32'd117914: dataIn1 = 32'd74
; 
32'd117915: dataIn1 = 32'd85
; 
32'd117916: dataIn1 = 32'd2238
; 
32'd117917: dataIn1 = 32'd2239
; 
32'd117918: dataIn1 = 32'd2240
; 
32'd117919: dataIn1 = 32'd2265
; 
32'd117920: dataIn1 = 32'd3725
; 
32'd117921: dataIn1 = 32'd3729
; 
32'd117922: dataIn1 = 32'd5311
; 
32'd117923: dataIn1 = 32'd75
; 
32'd117924: dataIn1 = 32'd85
; 
32'd117925: dataIn1 = 32'd86
; 
32'd117926: dataIn1 = 32'd5311
; 
32'd117927: dataIn1 = 32'd5312
; 
32'd117928: dataIn1 = 32'd5455
; 
32'd117929: dataIn1 = 32'd76
; 
32'd117930: dataIn1 = 32'd3737
; 
32'd117931: dataIn1 = 32'd3738
; 
32'd117932: dataIn1 = 32'd3824
; 
32'd117933: dataIn1 = 32'd77
; 
32'd117934: dataIn1 = 32'd3739
; 
32'd117935: dataIn1 = 32'd3740
; 
32'd117936: dataIn1 = 32'd3745
; 
32'd117937: dataIn1 = 32'd3752
; 
32'd117938: dataIn1 = 32'd3825
; 
32'd117939: dataIn1 = 32'd3827
; 
32'd117940: dataIn1 = 32'd78
; 
32'd117941: dataIn1 = 32'd3753
; 
32'd117942: dataIn1 = 32'd3754
; 
32'd117943: dataIn1 = 32'd3759
; 
32'd117944: dataIn1 = 32'd3765
; 
32'd117945: dataIn1 = 32'd3835
; 
32'd117946: dataIn1 = 32'd3837
; 
32'd117947: dataIn1 = 32'd79
; 
32'd117948: dataIn1 = 32'd3766
; 
32'd117949: dataIn1 = 32'd3767
; 
32'd117950: dataIn1 = 32'd3771
; 
32'd117951: dataIn1 = 32'd3777
; 
32'd117952: dataIn1 = 32'd3847
; 
32'd117953: dataIn1 = 32'd3849
; 
32'd117954: dataIn1 = 32'd80
; 
32'd117955: dataIn1 = 32'd3778
; 
32'd117956: dataIn1 = 32'd3779
; 
32'd117957: dataIn1 = 32'd3783
; 
32'd117958: dataIn1 = 32'd3789
; 
32'd117959: dataIn1 = 32'd3853
; 
32'd117960: dataIn1 = 32'd3855
; 
32'd117961: dataIn1 = 32'd81
; 
32'd117962: dataIn1 = 32'd3790
; 
32'd117963: dataIn1 = 32'd3791
; 
32'd117964: dataIn1 = 32'd3795
; 
32'd117965: dataIn1 = 32'd3801
; 
32'd117966: dataIn1 = 32'd3859
; 
32'd117967: dataIn1 = 32'd3861
; 
32'd117968: dataIn1 = 32'd82
; 
32'd117969: dataIn1 = 32'd2282
; 
32'd117970: dataIn1 = 32'd2284
; 
32'd117971: dataIn1 = 32'd3802
; 
32'd117972: dataIn1 = 32'd3803
; 
32'd117973: dataIn1 = 32'd3807
; 
32'd117974: dataIn1 = 32'd3813
; 
32'd117975: dataIn1 = 32'd83
; 
32'd117976: dataIn1 = 32'd94
; 
32'd117977: dataIn1 = 32'd2263
; 
32'd117978: dataIn1 = 32'd2285
; 
32'd117979: dataIn1 = 32'd3814
; 
32'd117980: dataIn1 = 32'd3815
; 
32'd117981: dataIn1 = 32'd3819
; 
32'd117982: dataIn1 = 32'd84
; 
32'd117983: dataIn1 = 32'd85
; 
32'd117984: dataIn1 = 32'd94
; 
32'd117985: dataIn1 = 32'd95
; 
32'd117986: dataIn1 = 32'd2263
; 
32'd117987: dataIn1 = 32'd2264
; 
32'd117988: dataIn1 = 32'd2265
; 
32'd117989: dataIn1 = 32'd74
; 
32'd117990: dataIn1 = 32'd75
; 
32'd117991: dataIn1 = 32'd84
; 
32'd117992: dataIn1 = 32'd85
; 
32'd117993: dataIn1 = 32'd86
; 
32'd117994: dataIn1 = 32'd95
; 
32'd117995: dataIn1 = 32'd96
; 
32'd117996: dataIn1 = 32'd2265
; 
32'd117997: dataIn1 = 32'd5311
; 
32'd117998: dataIn1 = 32'd75
; 
32'd117999: dataIn1 = 32'd85
; 
32'd118000: dataIn1 = 32'd86
; 
32'd118001: dataIn1 = 32'd96
; 
32'd118002: dataIn1 = 32'd87
; 
32'd118003: dataIn1 = 32'd2266
; 
32'd118004: dataIn1 = 32'd2267
; 
32'd118005: dataIn1 = 32'd2268
; 
32'd118006: dataIn1 = 32'd3822
; 
32'd118007: dataIn1 = 32'd5313
; 
32'd118008: dataIn1 = 32'd5315
; 
32'd118009: dataIn1 = 32'd10288
; 
32'd118010: dataIn1 = 32'd88
; 
32'd118011: dataIn1 = 32'd3828
; 
32'd118012: dataIn1 = 32'd3829
; 
32'd118013: dataIn1 = 32'd3834
; 
32'd118014: dataIn1 = 32'd3839
; 
32'd118015: dataIn1 = 32'd5314
; 
32'd118016: dataIn1 = 32'd5317
; 
32'd118017: dataIn1 = 32'd89
; 
32'd118018: dataIn1 = 32'd100
; 
32'd118019: dataIn1 = 32'd2274
; 
32'd118020: dataIn1 = 32'd3840
; 
32'd118021: dataIn1 = 32'd3841
; 
32'd118022: dataIn1 = 32'd3846
; 
32'd118023: dataIn1 = 32'd5316
; 
32'd118024: dataIn1 = 32'd90
; 
32'd118025: dataIn1 = 32'd100
; 
32'd118026: dataIn1 = 32'd101
; 
32'd118027: dataIn1 = 32'd2274
; 
32'd118028: dataIn1 = 32'd2275
; 
32'd118029: dataIn1 = 32'd2276
; 
32'd118030: dataIn1 = 32'd2277
; 
32'd118031: dataIn1 = 32'd3851
; 
32'd118032: dataIn1 = 32'd91
; 
32'd118033: dataIn1 = 32'd101
; 
32'd118034: dataIn1 = 32'd102
; 
32'd118035: dataIn1 = 32'd2277
; 
32'd118036: dataIn1 = 32'd2278
; 
32'd118037: dataIn1 = 32'd2279
; 
32'd118038: dataIn1 = 32'd2280
; 
32'd118039: dataIn1 = 32'd3857
; 
32'd118040: dataIn1 = 32'd92
; 
32'd118041: dataIn1 = 32'd102
; 
32'd118042: dataIn1 = 32'd103
; 
32'd118043: dataIn1 = 32'd2280
; 
32'd118044: dataIn1 = 32'd2281
; 
32'd118045: dataIn1 = 32'd2282
; 
32'd118046: dataIn1 = 32'd2283
; 
32'd118047: dataIn1 = 32'd93
; 
32'd118048: dataIn1 = 32'd94
; 
32'd118049: dataIn1 = 32'd103
; 
32'd118050: dataIn1 = 32'd104
; 
32'd118051: dataIn1 = 32'd2283
; 
32'd118052: dataIn1 = 32'd2284
; 
32'd118053: dataIn1 = 32'd2285
; 
32'd118054: dataIn1 = 32'd83
; 
32'd118055: dataIn1 = 32'd84
; 
32'd118056: dataIn1 = 32'd93
; 
32'd118057: dataIn1 = 32'd94
; 
32'd118058: dataIn1 = 32'd95
; 
32'd118059: dataIn1 = 32'd104
; 
32'd118060: dataIn1 = 32'd105
; 
32'd118061: dataIn1 = 32'd2263
; 
32'd118062: dataIn1 = 32'd2285
; 
32'd118063: dataIn1 = 32'd84
; 
32'd118064: dataIn1 = 32'd85
; 
32'd118065: dataIn1 = 32'd94
; 
32'd118066: dataIn1 = 32'd95
; 
32'd118067: dataIn1 = 32'd96
; 
32'd118068: dataIn1 = 32'd105
; 
32'd118069: dataIn1 = 32'd106
; 
32'd118070: dataIn1 = 32'd85
; 
32'd118071: dataIn1 = 32'd86
; 
32'd118072: dataIn1 = 32'd95
; 
32'd118073: dataIn1 = 32'd96
; 
32'd118074: dataIn1 = 32'd106
; 
32'd118075: dataIn1 = 32'd107
; 
32'd118076: dataIn1 = 32'd97
; 
32'd118077: dataIn1 = 32'd98
; 
32'd118078: dataIn1 = 32'd5315
; 
32'd118079: dataIn1 = 32'd10288
; 
32'd118080: dataIn1 = 32'd97
; 
32'd118081: dataIn1 = 32'd98
; 
32'd118082: dataIn1 = 32'd5314
; 
32'd118083: dataIn1 = 32'd5315
; 
32'd118084: dataIn1 = 32'd5456
; 
32'd118085: dataIn1 = 32'd99
; 
32'd118086: dataIn1 = 32'd5316
; 
32'd118087: dataIn1 = 32'd5317
; 
32'd118088: dataIn1 = 32'd5456
; 
32'd118089: dataIn1 = 32'd10289
; 
32'd118090: dataIn1 = 32'd89
; 
32'd118091: dataIn1 = 32'd90
; 
32'd118092: dataIn1 = 32'd100
; 
32'd118093: dataIn1 = 32'd101
; 
32'd118094: dataIn1 = 32'd2274
; 
32'd118095: dataIn1 = 32'd5316
; 
32'd118096: dataIn1 = 32'd10289
; 
32'd118097: dataIn1 = 32'd90
; 
32'd118098: dataIn1 = 32'd91
; 
32'd118099: dataIn1 = 32'd100
; 
32'd118100: dataIn1 = 32'd101
; 
32'd118101: dataIn1 = 32'd102
; 
32'd118102: dataIn1 = 32'd2277
; 
32'd118103: dataIn1 = 32'd91
; 
32'd118104: dataIn1 = 32'd92
; 
32'd118105: dataIn1 = 32'd101
; 
32'd118106: dataIn1 = 32'd102
; 
32'd118107: dataIn1 = 32'd103
; 
32'd118108: dataIn1 = 32'd2280
; 
32'd118109: dataIn1 = 32'd92
; 
32'd118110: dataIn1 = 32'd93
; 
32'd118111: dataIn1 = 32'd102
; 
32'd118112: dataIn1 = 32'd103
; 
32'd118113: dataIn1 = 32'd104
; 
32'd118114: dataIn1 = 32'd2283
; 
32'd118115: dataIn1 = 32'd93
; 
32'd118116: dataIn1 = 32'd94
; 
32'd118117: dataIn1 = 32'd103
; 
32'd118118: dataIn1 = 32'd104
; 
32'd118119: dataIn1 = 32'd105
; 
32'd118120: dataIn1 = 32'd94
; 
32'd118121: dataIn1 = 32'd95
; 
32'd118122: dataIn1 = 32'd104
; 
32'd118123: dataIn1 = 32'd105
; 
32'd118124: dataIn1 = 32'd106
; 
32'd118125: dataIn1 = 32'd95
; 
32'd118126: dataIn1 = 32'd96
; 
32'd118127: dataIn1 = 32'd105
; 
32'd118128: dataIn1 = 32'd106
; 
32'd118129: dataIn1 = 32'd107
; 
32'd118130: dataIn1 = 32'd96
; 
32'd118131: dataIn1 = 32'd106
; 
32'd118132: dataIn1 = 32'd107
; 
32'd118133: dataIn1 = 32'd108
; 
32'd118134: dataIn1 = 32'd1720
; 
32'd118135: dataIn1 = 32'd1721
; 
32'd118136: dataIn1 = 32'd1722
; 
32'd118137: dataIn1 = 32'd5527
; 
32'd118138: dataIn1 = 32'd5528
; 
32'd118139: dataIn1 = 32'd5529
; 
32'd118140: dataIn1 = 32'd109
; 
32'd118141: dataIn1 = 32'd5328
; 
32'd118142: dataIn1 = 32'd5329
; 
32'd118143: dataIn1 = 32'd5460
; 
32'd118144: dataIn1 = 32'd5461
; 
32'd118145: dataIn1 = 32'd5536
; 
32'd118146: dataIn1 = 32'd5537
; 
32'd118147: dataIn1 = 32'd110
; 
32'd118148: dataIn1 = 32'd5336
; 
32'd118149: dataIn1 = 32'd5337
; 
32'd118150: dataIn1 = 32'd5464
; 
32'd118151: dataIn1 = 32'd5465
; 
32'd118152: dataIn1 = 32'd5544
; 
32'd118153: dataIn1 = 32'd5545
; 
32'd118154: dataIn1 = 32'd111
; 
32'd118155: dataIn1 = 32'd5344
; 
32'd118156: dataIn1 = 32'd5345
; 
32'd118157: dataIn1 = 32'd5468
; 
32'd118158: dataIn1 = 32'd5469
; 
32'd118159: dataIn1 = 32'd5552
; 
32'd118160: dataIn1 = 32'd5553
; 
32'd118161: dataIn1 = 32'd112
; 
32'd118162: dataIn1 = 32'd5352
; 
32'd118163: dataIn1 = 32'd5353
; 
32'd118164: dataIn1 = 32'd5472
; 
32'd118165: dataIn1 = 32'd5473
; 
32'd118166: dataIn1 = 32'd5560
; 
32'd118167: dataIn1 = 32'd5561
; 
32'd118168: dataIn1 = 32'd113
; 
32'd118169: dataIn1 = 32'd5360
; 
32'd118170: dataIn1 = 32'd5361
; 
32'd118171: dataIn1 = 32'd5476
; 
32'd118172: dataIn1 = 32'd5477
; 
32'd118173: dataIn1 = 32'd5568
; 
32'd118174: dataIn1 = 32'd5569
; 
32'd118175: dataIn1 = 32'd114
; 
32'd118176: dataIn1 = 32'd5368
; 
32'd118177: dataIn1 = 32'd5369
; 
32'd118178: dataIn1 = 32'd5480
; 
32'd118179: dataIn1 = 32'd5481
; 
32'd118180: dataIn1 = 32'd5576
; 
32'd118181: dataIn1 = 32'd5577
; 
32'd118182: dataIn1 = 32'd115
; 
32'd118183: dataIn1 = 32'd5376
; 
32'd118184: dataIn1 = 32'd5377
; 
32'd118185: dataIn1 = 32'd5484
; 
32'd118186: dataIn1 = 32'd5485
; 
32'd118187: dataIn1 = 32'd5584
; 
32'd118188: dataIn1 = 32'd5585
; 
32'd118189: dataIn1 = 32'd116
; 
32'd118190: dataIn1 = 32'd5384
; 
32'd118191: dataIn1 = 32'd5385
; 
32'd118192: dataIn1 = 32'd5488
; 
32'd118193: dataIn1 = 32'd5489
; 
32'd118194: dataIn1 = 32'd5592
; 
32'd118195: dataIn1 = 32'd5593
; 
32'd118196: dataIn1 = 32'd117
; 
32'd118197: dataIn1 = 32'd5392
; 
32'd118198: dataIn1 = 32'd5393
; 
32'd118199: dataIn1 = 32'd5492
; 
32'd118200: dataIn1 = 32'd5493
; 
32'd118201: dataIn1 = 32'd5600
; 
32'd118202: dataIn1 = 32'd5601
; 
32'd118203: dataIn1 = 32'd118
; 
32'd118204: dataIn1 = 32'd5400
; 
32'd118205: dataIn1 = 32'd5401
; 
32'd118206: dataIn1 = 32'd5496
; 
32'd118207: dataIn1 = 32'd5497
; 
32'd118208: dataIn1 = 32'd5608
; 
32'd118209: dataIn1 = 32'd5609
; 
32'd118210: dataIn1 = 32'd119
; 
32'd118211: dataIn1 = 32'd5408
; 
32'd118212: dataIn1 = 32'd5409
; 
32'd118213: dataIn1 = 32'd5500
; 
32'd118214: dataIn1 = 32'd5501
; 
32'd118215: dataIn1 = 32'd5616
; 
32'd118216: dataIn1 = 32'd5617
; 
32'd118217: dataIn1 = 32'd120
; 
32'd118218: dataIn1 = 32'd5416
; 
32'd118219: dataIn1 = 32'd5417
; 
32'd118220: dataIn1 = 32'd5504
; 
32'd118221: dataIn1 = 32'd5505
; 
32'd118222: dataIn1 = 32'd5624
; 
32'd118223: dataIn1 = 32'd5625
; 
32'd118224: dataIn1 = 32'd121
; 
32'd118225: dataIn1 = 32'd5424
; 
32'd118226: dataIn1 = 32'd5425
; 
32'd118227: dataIn1 = 32'd5508
; 
32'd118228: dataIn1 = 32'd5632
; 
32'd118229: dataIn1 = 32'd122
; 
32'd118230: dataIn1 = 32'd965
; 
32'd118231: dataIn1 = 32'd966
; 
32'd118232: dataIn1 = 32'd1035
; 
32'd118233: dataIn1 = 32'd1036
; 
32'd118234: dataIn1 = 32'd2031
; 
32'd118235: dataIn1 = 32'd2033
; 
32'd118236: dataIn1 = 32'd3480
; 
32'd118237: dataIn1 = 32'd3484
; 
32'd118238: dataIn1 = 32'd123
; 
32'd118239: dataIn1 = 32'd963
; 
32'd118240: dataIn1 = 32'd1034
; 
32'd118241: dataIn1 = 32'd2032
; 
32'd118242: dataIn1 = 32'd3496
; 
32'd118243: dataIn1 = 32'd124
; 
32'd118244: dataIn1 = 32'd4640
; 
32'd118245: dataIn1 = 32'd4641
; 
32'd118246: dataIn1 = 32'd9677
; 
32'd118247: dataIn1 = 32'd9679
; 
32'd118248: dataIn1 = 32'd9704
; 
32'd118249: dataIn1 = 32'd9724
; 
32'd118250: dataIn1 = 32'd125
; 
32'd118251: dataIn1 = 32'd971
; 
32'd118252: dataIn1 = 32'd972
; 
32'd118253: dataIn1 = 32'd1037
; 
32'd118254: dataIn1 = 32'd1038
; 
32'd118255: dataIn1 = 32'd2040
; 
32'd118256: dataIn1 = 32'd3455
; 
32'd118257: dataIn1 = 32'd3465
; 
32'd118258: dataIn1 = 32'd126
; 
32'd118259: dataIn1 = 32'd3864
; 
32'd118260: dataIn1 = 32'd3865
; 
32'd118261: dataIn1 = 32'd3866
; 
32'd118262: dataIn1 = 32'd4610
; 
32'd118263: dataIn1 = 32'd5951
; 
32'd118264: dataIn1 = 32'd5952
; 
32'd118265: dataIn1 = 32'd127
; 
32'd118266: dataIn1 = 32'd5666
; 
32'd118267: dataIn1 = 32'd5667
; 
32'd118268: dataIn1 = 32'd5787
; 
32'd118269: dataIn1 = 32'd5944
; 
32'd118270: dataIn1 = 32'd6892
; 
32'd118271: dataIn1 = 32'd6893
; 
32'd118272: dataIn1 = 32'd128
; 
32'd118273: dataIn1 = 32'd3891
; 
32'd118274: dataIn1 = 32'd3892
; 
32'd118275: dataIn1 = 32'd3925
; 
32'd118276: dataIn1 = 32'd3926
; 
32'd118277: dataIn1 = 32'd4603
; 
32'd118278: dataIn1 = 32'd5427
; 
32'd118279: dataIn1 = 32'd129
; 
32'd118280: dataIn1 = 32'd2526
; 
32'd118281: dataIn1 = 32'd2528
; 
32'd118282: dataIn1 = 32'd5721
; 
32'd118283: dataIn1 = 32'd5722
; 
32'd118284: dataIn1 = 32'd5936
; 
32'd118285: dataIn1 = 32'd5937
; 
32'd118286: dataIn1 = 32'd130
; 
32'd118287: dataIn1 = 32'd5902
; 
32'd118288: dataIn1 = 32'd5903
; 
32'd118289: dataIn1 = 32'd5972
; 
32'd118290: dataIn1 = 32'd6033
; 
32'd118291: dataIn1 = 32'd7237
; 
32'd118292: dataIn1 = 32'd7238
; 
32'd118293: dataIn1 = 32'd131
; 
32'd118294: dataIn1 = 32'd4604
; 
32'd118295: dataIn1 = 32'd4605
; 
32'd118296: dataIn1 = 32'd4621
; 
32'd118297: dataIn1 = 32'd4635
; 
32'd118298: dataIn1 = 32'd5980
; 
32'd118299: dataIn1 = 32'd5982
; 
32'd118300: dataIn1 = 32'd132
; 
32'd118301: dataIn1 = 32'd984
; 
32'd118302: dataIn1 = 32'd985
; 
32'd118303: dataIn1 = 32'd1043
; 
32'd118304: dataIn1 = 32'd1044
; 
32'd118305: dataIn1 = 32'd2052
; 
32'd118306: dataIn1 = 32'd3431
; 
32'd118307: dataIn1 = 32'd3432
; 
32'd118308: dataIn1 = 32'd133
; 
32'd118309: dataIn1 = 32'd7404
; 
32'd118310: dataIn1 = 32'd7405
; 
32'd118311: dataIn1 = 32'd7489
; 
32'd118312: dataIn1 = 32'd7576
; 
32'd118313: dataIn1 = 32'd9603
; 
32'd118314: dataIn1 = 32'd9604
; 
32'd118315: dataIn1 = 32'd134
; 
32'd118316: dataIn1 = 32'd990
; 
32'd118317: dataIn1 = 32'd991
; 
32'd118318: dataIn1 = 32'd1045
; 
32'd118319: dataIn1 = 32'd1046
; 
32'd118320: dataIn1 = 32'd2059
; 
32'd118321: dataIn1 = 32'd3473
; 
32'd118322: dataIn1 = 32'd3477
; 
32'd118323: dataIn1 = 32'd135
; 
32'd118324: dataIn1 = 32'd992
; 
32'd118325: dataIn1 = 32'd993
; 
32'd118326: dataIn1 = 32'd1047
; 
32'd118327: dataIn1 = 32'd1048
; 
32'd118328: dataIn1 = 32'd2060
; 
32'd118329: dataIn1 = 32'd3489
; 
32'd118330: dataIn1 = 32'd3493
; 
32'd118331: dataIn1 = 32'd136
; 
32'd118332: dataIn1 = 32'd7655
; 
32'd118333: dataIn1 = 32'd7656
; 
32'd118334: dataIn1 = 32'd7742
; 
32'd118335: dataIn1 = 32'd7829
; 
32'd118336: dataIn1 = 32'd9609
; 
32'd118337: dataIn1 = 32'd9610
; 
32'd118338: dataIn1 = 32'd137
; 
32'd118339: dataIn1 = 32'd998
; 
32'd118340: dataIn1 = 32'd999
; 
32'd118341: dataIn1 = 32'd1049
; 
32'd118342: dataIn1 = 32'd1050
; 
32'd118343: dataIn1 = 32'd2067
; 
32'd118344: dataIn1 = 32'd3503
; 
32'd118345: dataIn1 = 32'd3505
; 
32'd118346: dataIn1 = 32'd138
; 
32'd118347: dataIn1 = 32'd1000
; 
32'd118348: dataIn1 = 32'd1001
; 
32'd118349: dataIn1 = 32'd1051
; 
32'd118350: dataIn1 = 32'd1052
; 
32'd118351: dataIn1 = 32'd2068
; 
32'd118352: dataIn1 = 32'd3511
; 
32'd118353: dataIn1 = 32'd3513
; 
32'd118354: dataIn1 = 32'd139
; 
32'd118355: dataIn1 = 32'd4723
; 
32'd118356: dataIn1 = 32'd4724
; 
32'd118357: dataIn1 = 32'd7908
; 
32'd118358: dataIn1 = 32'd7909
; 
32'd118359: dataIn1 = 32'd7995
; 
32'd118360: dataIn1 = 32'd8082
; 
32'd118361: dataIn1 = 32'd140
; 
32'd118362: dataIn1 = 32'd1006
; 
32'd118363: dataIn1 = 32'd1007
; 
32'd118364: dataIn1 = 32'd1053
; 
32'd118365: dataIn1 = 32'd1054
; 
32'd118366: dataIn1 = 32'd2075
; 
32'd118367: dataIn1 = 32'd3519
; 
32'd118368: dataIn1 = 32'd3521
; 
32'd118369: dataIn1 = 32'd141
; 
32'd118370: dataIn1 = 32'd1008
; 
32'd118371: dataIn1 = 32'd1009
; 
32'd118372: dataIn1 = 32'd1055
; 
32'd118373: dataIn1 = 32'd1056
; 
32'd118374: dataIn1 = 32'd2076
; 
32'd118375: dataIn1 = 32'd3527
; 
32'd118376: dataIn1 = 32'd3529
; 
32'd118377: dataIn1 = 32'd142
; 
32'd118378: dataIn1 = 32'd4741
; 
32'd118379: dataIn1 = 32'd4742
; 
32'd118380: dataIn1 = 32'd8161
; 
32'd118381: dataIn1 = 32'd8162
; 
32'd118382: dataIn1 = 32'd8248
; 
32'd118383: dataIn1 = 32'd8334
; 
32'd118384: dataIn1 = 32'd143
; 
32'd118385: dataIn1 = 32'd1014
; 
32'd118386: dataIn1 = 32'd1015
; 
32'd118387: dataIn1 = 32'd1057
; 
32'd118388: dataIn1 = 32'd1058
; 
32'd118389: dataIn1 = 32'd2083
; 
32'd118390: dataIn1 = 32'd3535
; 
32'd118391: dataIn1 = 32'd3537
; 
32'd118392: dataIn1 = 32'd144
; 
32'd118393: dataIn1 = 32'd1016
; 
32'd118394: dataIn1 = 32'd1017
; 
32'd118395: dataIn1 = 32'd1059
; 
32'd118396: dataIn1 = 32'd1060
; 
32'd118397: dataIn1 = 32'd2084
; 
32'd118398: dataIn1 = 32'd3543
; 
32'd118399: dataIn1 = 32'd3545
; 
32'd118400: dataIn1 = 32'd145
; 
32'd118401: dataIn1 = 32'd4759
; 
32'd118402: dataIn1 = 32'd4760
; 
32'd118403: dataIn1 = 32'd8413
; 
32'd118404: dataIn1 = 32'd8414
; 
32'd118405: dataIn1 = 32'd8500
; 
32'd118406: dataIn1 = 32'd8587
; 
32'd118407: dataIn1 = 32'd146
; 
32'd118408: dataIn1 = 32'd1022
; 
32'd118409: dataIn1 = 32'd1023
; 
32'd118410: dataIn1 = 32'd1061
; 
32'd118411: dataIn1 = 32'd1062
; 
32'd118412: dataIn1 = 32'd2091
; 
32'd118413: dataIn1 = 32'd3551
; 
32'd118414: dataIn1 = 32'd3553
; 
32'd118415: dataIn1 = 32'd147
; 
32'd118416: dataIn1 = 32'd1024
; 
32'd118417: dataIn1 = 32'd1025
; 
32'd118418: dataIn1 = 32'd1063
; 
32'd118419: dataIn1 = 32'd1064
; 
32'd118420: dataIn1 = 32'd2092
; 
32'd118421: dataIn1 = 32'd3559
; 
32'd118422: dataIn1 = 32'd3561
; 
32'd118423: dataIn1 = 32'd148
; 
32'd118424: dataIn1 = 32'd4777
; 
32'd118425: dataIn1 = 32'd4778
; 
32'd118426: dataIn1 = 32'd8666
; 
32'd118427: dataIn1 = 32'd8667
; 
32'd118428: dataIn1 = 32'd8753
; 
32'd118429: dataIn1 = 32'd8839
; 
32'd118430: dataIn1 = 32'd149
; 
32'd118431: dataIn1 = 32'd1030
; 
32'd118432: dataIn1 = 32'd1031
; 
32'd118433: dataIn1 = 32'd1065
; 
32'd118434: dataIn1 = 32'd1066
; 
32'd118435: dataIn1 = 32'd2096
; 
32'd118436: dataIn1 = 32'd2099
; 
32'd118437: dataIn1 = 32'd3567
; 
32'd118438: dataIn1 = 32'd3569
; 
32'd118439: dataIn1 = 32'd150
; 
32'd118440: dataIn1 = 32'd1033
; 
32'd118441: dataIn1 = 32'd1067
; 
32'd118442: dataIn1 = 32'd2100
; 
32'd118443: dataIn1 = 32'd3575
; 
32'd118444: dataIn1 = 32'd151
; 
32'd118445: dataIn1 = 32'd3422
; 
32'd118446: dataIn1 = 32'd3423
; 
32'd118447: dataIn1 = 32'd3450
; 
32'd118448: dataIn1 = 32'd3451
; 
32'd118449: dataIn1 = 32'd3463
; 
32'd118450: dataIn1 = 32'd3471
; 
32'd118451: dataIn1 = 32'd152
; 
32'd118452: dataIn1 = 32'd565
; 
32'd118453: dataIn1 = 32'd566
; 
32'd118454: dataIn1 = 32'd571
; 
32'd118455: dataIn1 = 32'd3499
; 
32'd118456: dataIn1 = 32'd3502
; 
32'd118457: dataIn1 = 32'd5457
; 
32'd118458: dataIn1 = 32'd153
; 
32'd118459: dataIn1 = 32'd5324
; 
32'd118460: dataIn1 = 32'd5325
; 
32'd118461: dataIn1 = 32'd5458
; 
32'd118462: dataIn1 = 32'd5459
; 
32'd118463: dataIn1 = 32'd5532
; 
32'd118464: dataIn1 = 32'd5533
; 
32'd118465: dataIn1 = 32'd154
; 
32'd118466: dataIn1 = 32'd2770
; 
32'd118467: dataIn1 = 32'd2771
; 
32'd118468: dataIn1 = 32'd3052
; 
32'd118469: dataIn1 = 32'd3932
; 
32'd118470: dataIn1 = 32'd3933
; 
32'd118471: dataIn1 = 32'd3960
; 
32'd118472: dataIn1 = 32'd155
; 
32'd118473: dataIn1 = 32'd2780
; 
32'd118474: dataIn1 = 32'd2781
; 
32'd118475: dataIn1 = 32'd3047
; 
32'd118476: dataIn1 = 32'd3061
; 
32'd118477: dataIn1 = 32'd4008
; 
32'd118478: dataIn1 = 32'd4009
; 
32'd118479: dataIn1 = 32'd156
; 
32'd118480: dataIn1 = 32'd2486
; 
32'd118481: dataIn1 = 32'd2487
; 
32'd118482: dataIn1 = 32'd2521
; 
32'd118483: dataIn1 = 32'd3420
; 
32'd118484: dataIn1 = 32'd3454
; 
32'd118485: dataIn1 = 32'd10265
; 
32'd118486: dataIn1 = 32'd157
; 
32'd118487: dataIn1 = 32'd2785
; 
32'd118488: dataIn1 = 32'd2786
; 
32'd118489: dataIn1 = 32'd3065
; 
32'd118490: dataIn1 = 32'd3072
; 
32'd118491: dataIn1 = 32'd4029
; 
32'd118492: dataIn1 = 32'd4030
; 
32'd118493: dataIn1 = 32'd158
; 
32'd118494: dataIn1 = 32'd5332
; 
32'd118495: dataIn1 = 32'd5333
; 
32'd118496: dataIn1 = 32'd5462
; 
32'd118497: dataIn1 = 32'd5463
; 
32'd118498: dataIn1 = 32'd5540
; 
32'd118499: dataIn1 = 32'd5541
; 
32'd118500: dataIn1 = 32'd159
; 
32'd118501: dataIn1 = 32'd2810
; 
32'd118502: dataIn1 = 32'd2811
; 
32'd118503: dataIn1 = 32'd3082
; 
32'd118504: dataIn1 = 32'd3107
; 
32'd118505: dataIn1 = 32'd4056
; 
32'd118506: dataIn1 = 32'd4057
; 
32'd118507: dataIn1 = 32'd160
; 
32'd118508: dataIn1 = 32'd5340
; 
32'd118509: dataIn1 = 32'd5341
; 
32'd118510: dataIn1 = 32'd5466
; 
32'd118511: dataIn1 = 32'd5467
; 
32'd118512: dataIn1 = 32'd5548
; 
32'd118513: dataIn1 = 32'd5549
; 
32'd118514: dataIn1 = 32'd161
; 
32'd118515: dataIn1 = 32'd2805
; 
32'd118516: dataIn1 = 32'd2806
; 
32'd118517: dataIn1 = 32'd3094
; 
32'd118518: dataIn1 = 32'd3102
; 
32'd118519: dataIn1 = 32'd4078
; 
32'd118520: dataIn1 = 32'd4079
; 
32'd118521: dataIn1 = 32'd162
; 
32'd118522: dataIn1 = 32'd2820
; 
32'd118523: dataIn1 = 32'd2821
; 
32'd118524: dataIn1 = 32'd3089
; 
32'd118525: dataIn1 = 32'd3117
; 
32'd118526: dataIn1 = 32'd4104
; 
32'd118527: dataIn1 = 32'd4105
; 
32'd118528: dataIn1 = 32'd163
; 
32'd118529: dataIn1 = 32'd2825
; 
32'd118530: dataIn1 = 32'd2826
; 
32'd118531: dataIn1 = 32'd3121
; 
32'd118532: dataIn1 = 32'd3128
; 
32'd118533: dataIn1 = 32'd4125
; 
32'd118534: dataIn1 = 32'd4126
; 
32'd118535: dataIn1 = 32'd164
; 
32'd118536: dataIn1 = 32'd5348
; 
32'd118537: dataIn1 = 32'd5349
; 
32'd118538: dataIn1 = 32'd5470
; 
32'd118539: dataIn1 = 32'd5471
; 
32'd118540: dataIn1 = 32'd5556
; 
32'd118541: dataIn1 = 32'd5557
; 
32'd118542: dataIn1 = 32'd165
; 
32'd118543: dataIn1 = 32'd2850
; 
32'd118544: dataIn1 = 32'd2851
; 
32'd118545: dataIn1 = 32'd3138
; 
32'd118546: dataIn1 = 32'd3163
; 
32'd118547: dataIn1 = 32'd4152
; 
32'd118548: dataIn1 = 32'd4153
; 
32'd118549: dataIn1 = 32'd166
; 
32'd118550: dataIn1 = 32'd5356
; 
32'd118551: dataIn1 = 32'd5357
; 
32'd118552: dataIn1 = 32'd5474
; 
32'd118553: dataIn1 = 32'd5475
; 
32'd118554: dataIn1 = 32'd5564
; 
32'd118555: dataIn1 = 32'd5565
; 
32'd118556: dataIn1 = 32'd167
; 
32'd118557: dataIn1 = 32'd2845
; 
32'd118558: dataIn1 = 32'd2846
; 
32'd118559: dataIn1 = 32'd3150
; 
32'd118560: dataIn1 = 32'd3158
; 
32'd118561: dataIn1 = 32'd4174
; 
32'd118562: dataIn1 = 32'd4175
; 
32'd118563: dataIn1 = 32'd168
; 
32'd118564: dataIn1 = 32'd2860
; 
32'd118565: dataIn1 = 32'd2861
; 
32'd118566: dataIn1 = 32'd3145
; 
32'd118567: dataIn1 = 32'd3173
; 
32'd118568: dataIn1 = 32'd4200
; 
32'd118569: dataIn1 = 32'd4201
; 
32'd118570: dataIn1 = 32'd169
; 
32'd118571: dataIn1 = 32'd2865
; 
32'd118572: dataIn1 = 32'd2866
; 
32'd118573: dataIn1 = 32'd3177
; 
32'd118574: dataIn1 = 32'd3184
; 
32'd118575: dataIn1 = 32'd4221
; 
32'd118576: dataIn1 = 32'd4222
; 
32'd118577: dataIn1 = 32'd170
; 
32'd118578: dataIn1 = 32'd5364
; 
32'd118579: dataIn1 = 32'd5365
; 
32'd118580: dataIn1 = 32'd5478
; 
32'd118581: dataIn1 = 32'd5479
; 
32'd118582: dataIn1 = 32'd5572
; 
32'd118583: dataIn1 = 32'd5573
; 
32'd118584: dataIn1 = 32'd171
; 
32'd118585: dataIn1 = 32'd2890
; 
32'd118586: dataIn1 = 32'd2891
; 
32'd118587: dataIn1 = 32'd3194
; 
32'd118588: dataIn1 = 32'd3219
; 
32'd118589: dataIn1 = 32'd4248
; 
32'd118590: dataIn1 = 32'd4249
; 
32'd118591: dataIn1 = 32'd172
; 
32'd118592: dataIn1 = 32'd5372
; 
32'd118593: dataIn1 = 32'd5373
; 
32'd118594: dataIn1 = 32'd5482
; 
32'd118595: dataIn1 = 32'd5483
; 
32'd118596: dataIn1 = 32'd5580
; 
32'd118597: dataIn1 = 32'd5581
; 
32'd118598: dataIn1 = 32'd173
; 
32'd118599: dataIn1 = 32'd2885
; 
32'd118600: dataIn1 = 32'd2886
; 
32'd118601: dataIn1 = 32'd3206
; 
32'd118602: dataIn1 = 32'd3214
; 
32'd118603: dataIn1 = 32'd4270
; 
32'd118604: dataIn1 = 32'd4271
; 
32'd118605: dataIn1 = 32'd174
; 
32'd118606: dataIn1 = 32'd2900
; 
32'd118607: dataIn1 = 32'd2901
; 
32'd118608: dataIn1 = 32'd3201
; 
32'd118609: dataIn1 = 32'd3229
; 
32'd118610: dataIn1 = 32'd4296
; 
32'd118611: dataIn1 = 32'd4297
; 
32'd118612: dataIn1 = 32'd175
; 
32'd118613: dataIn1 = 32'd2905
; 
32'd118614: dataIn1 = 32'd2906
; 
32'd118615: dataIn1 = 32'd3233
; 
32'd118616: dataIn1 = 32'd3240
; 
32'd118617: dataIn1 = 32'd4317
; 
32'd118618: dataIn1 = 32'd4318
; 
32'd118619: dataIn1 = 32'd176
; 
32'd118620: dataIn1 = 32'd5380
; 
32'd118621: dataIn1 = 32'd5381
; 
32'd118622: dataIn1 = 32'd5486
; 
32'd118623: dataIn1 = 32'd5487
; 
32'd118624: dataIn1 = 32'd5588
; 
32'd118625: dataIn1 = 32'd5589
; 
32'd118626: dataIn1 = 32'd177
; 
32'd118627: dataIn1 = 32'd2930
; 
32'd118628: dataIn1 = 32'd2931
; 
32'd118629: dataIn1 = 32'd3250
; 
32'd118630: dataIn1 = 32'd3275
; 
32'd118631: dataIn1 = 32'd4344
; 
32'd118632: dataIn1 = 32'd4345
; 
32'd118633: dataIn1 = 32'd178
; 
32'd118634: dataIn1 = 32'd5388
; 
32'd118635: dataIn1 = 32'd5389
; 
32'd118636: dataIn1 = 32'd5490
; 
32'd118637: dataIn1 = 32'd5491
; 
32'd118638: dataIn1 = 32'd5596
; 
32'd118639: dataIn1 = 32'd5597
; 
32'd118640: dataIn1 = 32'd179
; 
32'd118641: dataIn1 = 32'd2925
; 
32'd118642: dataIn1 = 32'd2926
; 
32'd118643: dataIn1 = 32'd3262
; 
32'd118644: dataIn1 = 32'd3270
; 
32'd118645: dataIn1 = 32'd4366
; 
32'd118646: dataIn1 = 32'd4367
; 
32'd118647: dataIn1 = 32'd180
; 
32'd118648: dataIn1 = 32'd2940
; 
32'd118649: dataIn1 = 32'd2941
; 
32'd118650: dataIn1 = 32'd3257
; 
32'd118651: dataIn1 = 32'd3285
; 
32'd118652: dataIn1 = 32'd4392
; 
32'd118653: dataIn1 = 32'd4393
; 
32'd118654: dataIn1 = 32'd181
; 
32'd118655: dataIn1 = 32'd2945
; 
32'd118656: dataIn1 = 32'd2946
; 
32'd118657: dataIn1 = 32'd3289
; 
32'd118658: dataIn1 = 32'd3296
; 
32'd118659: dataIn1 = 32'd4413
; 
32'd118660: dataIn1 = 32'd4414
; 
32'd118661: dataIn1 = 32'd182
; 
32'd118662: dataIn1 = 32'd5396
; 
32'd118663: dataIn1 = 32'd5397
; 
32'd118664: dataIn1 = 32'd5494
; 
32'd118665: dataIn1 = 32'd5495
; 
32'd118666: dataIn1 = 32'd5604
; 
32'd118667: dataIn1 = 32'd5605
; 
32'd118668: dataIn1 = 32'd183
; 
32'd118669: dataIn1 = 32'd2970
; 
32'd118670: dataIn1 = 32'd2971
; 
32'd118671: dataIn1 = 32'd3306
; 
32'd118672: dataIn1 = 32'd3331
; 
32'd118673: dataIn1 = 32'd4440
; 
32'd118674: dataIn1 = 32'd4441
; 
32'd118675: dataIn1 = 32'd184
; 
32'd118676: dataIn1 = 32'd5404
; 
32'd118677: dataIn1 = 32'd5405
; 
32'd118678: dataIn1 = 32'd5498
; 
32'd118679: dataIn1 = 32'd5499
; 
32'd118680: dataIn1 = 32'd5612
; 
32'd118681: dataIn1 = 32'd5613
; 
32'd118682: dataIn1 = 32'd185
; 
32'd118683: dataIn1 = 32'd2965
; 
32'd118684: dataIn1 = 32'd2966
; 
32'd118685: dataIn1 = 32'd3318
; 
32'd118686: dataIn1 = 32'd3326
; 
32'd118687: dataIn1 = 32'd4462
; 
32'd118688: dataIn1 = 32'd4463
; 
32'd118689: dataIn1 = 32'd186
; 
32'd118690: dataIn1 = 32'd2980
; 
32'd118691: dataIn1 = 32'd2981
; 
32'd118692: dataIn1 = 32'd3313
; 
32'd118693: dataIn1 = 32'd3341
; 
32'd118694: dataIn1 = 32'd4488
; 
32'd118695: dataIn1 = 32'd4489
; 
32'd118696: dataIn1 = 32'd187
; 
32'd118697: dataIn1 = 32'd2985
; 
32'd118698: dataIn1 = 32'd2986
; 
32'd118699: dataIn1 = 32'd3345
; 
32'd118700: dataIn1 = 32'd3352
; 
32'd118701: dataIn1 = 32'd4509
; 
32'd118702: dataIn1 = 32'd4510
; 
32'd118703: dataIn1 = 32'd188
; 
32'd118704: dataIn1 = 32'd5412
; 
32'd118705: dataIn1 = 32'd5413
; 
32'd118706: dataIn1 = 32'd5502
; 
32'd118707: dataIn1 = 32'd5503
; 
32'd118708: dataIn1 = 32'd5620
; 
32'd118709: dataIn1 = 32'd5621
; 
32'd118710: dataIn1 = 32'd189
; 
32'd118711: dataIn1 = 32'd3010
; 
32'd118712: dataIn1 = 32'd3011
; 
32'd118713: dataIn1 = 32'd3362
; 
32'd118714: dataIn1 = 32'd3387
; 
32'd118715: dataIn1 = 32'd4536
; 
32'd118716: dataIn1 = 32'd4537
; 
32'd118717: dataIn1 = 32'd190
; 
32'd118718: dataIn1 = 32'd5420
; 
32'd118719: dataIn1 = 32'd5421
; 
32'd118720: dataIn1 = 32'd5506
; 
32'd118721: dataIn1 = 32'd5507
; 
32'd118722: dataIn1 = 32'd5628
; 
32'd118723: dataIn1 = 32'd5629
; 
32'd118724: dataIn1 = 32'd191
; 
32'd118725: dataIn1 = 32'd3005
; 
32'd118726: dataIn1 = 32'd3006
; 
32'd118727: dataIn1 = 32'd3374
; 
32'd118728: dataIn1 = 32'd3382
; 
32'd118729: dataIn1 = 32'd4558
; 
32'd118730: dataIn1 = 32'd4559
; 
32'd118731: dataIn1 = 32'd192
; 
32'd118732: dataIn1 = 32'd3020
; 
32'd118733: dataIn1 = 32'd3021
; 
32'd118734: dataIn1 = 32'd3369
; 
32'd118735: dataIn1 = 32'd3397
; 
32'd118736: dataIn1 = 32'd4584
; 
32'd118737: dataIn1 = 32'd4585
; 
32'd118738: dataIn1 = 32'd193
; 
32'd118739: dataIn1 = 32'd3025
; 
32'd118740: dataIn1 = 32'd3026
; 
32'd118741: dataIn1 = 32'd3401
; 
32'd118742: dataIn1 = 32'd5305
; 
32'd118743: dataIn1 = 32'd194
; 
32'd118744: dataIn1 = 32'd1397
; 
32'd118745: dataIn1 = 32'd1401
; 
32'd118746: dataIn1 = 32'd1830
; 
32'd118747: dataIn1 = 32'd10753
; 
32'd118748: dataIn1 = 32'd10754
; 
32'd118749: dataIn1 = 32'd195
; 
32'd118750: dataIn1 = 32'd962
; 
32'd118751: dataIn1 = 32'd1034
; 
32'd118752: dataIn1 = 32'd1035
; 
32'd118753: dataIn1 = 32'd2029
; 
32'd118754: dataIn1 = 32'd2030
; 
32'd118755: dataIn1 = 32'd3488
; 
32'd118756: dataIn1 = 32'd3492
; 
32'd118757: dataIn1 = 32'd196
; 
32'd118758: dataIn1 = 32'd1400
; 
32'd118759: dataIn1 = 32'd1408
; 
32'd118760: dataIn1 = 32'd1839
; 
32'd118761: dataIn1 = 32'd10744
; 
32'd118762: dataIn1 = 32'd10745
; 
32'd118763: dataIn1 = 32'd197
; 
32'd118764: dataIn1 = 32'd1403
; 
32'd118765: dataIn1 = 32'd1836
; 
32'd118766: dataIn1 = 32'd10760
; 
32'd118767: dataIn1 = 32'd10761
; 
32'd118768: dataIn1 = 32'd198
; 
32'd118769: dataIn1 = 32'd1406
; 
32'd118770: dataIn1 = 32'd1410
; 
32'd118771: dataIn1 = 32'd1837
; 
32'd118772: dataIn1 = 32'd1841
; 
32'd118773: dataIn1 = 32'd10736
; 
32'd118774: dataIn1 = 32'd10737
; 
32'd118775: dataIn1 = 32'd199
; 
32'd118776: dataIn1 = 32'd967
; 
32'd118777: dataIn1 = 32'd968
; 
32'd118778: dataIn1 = 32'd1036
; 
32'd118779: dataIn1 = 32'd1037
; 
32'd118780: dataIn1 = 32'd2035
; 
32'd118781: dataIn1 = 32'd3472
; 
32'd118782: dataIn1 = 32'd3476
; 
32'd118783: dataIn1 = 32'd200
; 
32'd118784: dataIn1 = 32'd1412
; 
32'd118785: dataIn1 = 32'd1419
; 
32'd118786: dataIn1 = 32'd1843
; 
32'd118787: dataIn1 = 32'd1852
; 
32'd118788: dataIn1 = 32'd10728
; 
32'd118789: dataIn1 = 32'd10729
; 
32'd118790: dataIn1 = 32'd201
; 
32'd118791: dataIn1 = 32'd1413
; 
32'd118792: dataIn1 = 32'd1417
; 
32'd118793: dataIn1 = 32'd1846
; 
32'd118794: dataIn1 = 32'd1850
; 
32'd118795: dataIn1 = 32'd10720
; 
32'd118796: dataIn1 = 32'd10721
; 
32'd118797: dataIn1 = 32'd202
; 
32'd118798: dataIn1 = 32'd969
; 
32'd118799: dataIn1 = 32'd970
; 
32'd118800: dataIn1 = 32'd1038
; 
32'd118801: dataIn1 = 32'd1039
; 
32'd118802: dataIn1 = 32'd2038
; 
32'd118803: dataIn1 = 32'd2534
; 
32'd118804: dataIn1 = 32'd2553
; 
32'd118805: dataIn1 = 32'd3430
; 
32'd118806: dataIn1 = 32'd203
; 
32'd118807: dataIn1 = 32'd1416
; 
32'd118808: dataIn1 = 32'd1426
; 
32'd118809: dataIn1 = 32'd3409
; 
32'd118810: dataIn1 = 32'd3410
; 
32'd118811: dataIn1 = 32'd10712
; 
32'd118812: dataIn1 = 32'd10713
; 
32'd118813: dataIn1 = 32'd204
; 
32'd118814: dataIn1 = 32'd1430
; 
32'd118815: dataIn1 = 32'd1440
; 
32'd118816: dataIn1 = 32'd3414
; 
32'd118817: dataIn1 = 32'd3416
; 
32'd118818: dataIn1 = 32'd10551
; 
32'd118819: dataIn1 = 32'd10552
; 
32'd118820: dataIn1 = 32'd10553
; 
32'd118821: dataIn1 = 32'd205
; 
32'd118822: dataIn1 = 32'd3874
; 
32'd118823: dataIn1 = 32'd3875
; 
32'd118824: dataIn1 = 32'd3890
; 
32'd118825: dataIn1 = 32'd3897
; 
32'd118826: dataIn1 = 32'd4602
; 
32'd118827: dataIn1 = 32'd5426
; 
32'd118828: dataIn1 = 32'd5656
; 
32'd118829: dataIn1 = 32'd206
; 
32'd118830: dataIn1 = 32'd2290
; 
32'd118831: dataIn1 = 32'd2291
; 
32'd118832: dataIn1 = 32'd2293
; 
32'd118833: dataIn1 = 32'd2527
; 
32'd118834: dataIn1 = 32'd3905
; 
32'd118835: dataIn1 = 32'd3906
; 
32'd118836: dataIn1 = 32'd5703
; 
32'd118837: dataIn1 = 32'd207
; 
32'd118838: dataIn1 = 32'd767
; 
32'd118839: dataIn1 = 32'd1463
; 
32'd118840: dataIn1 = 32'd1487
; 
32'd118841: dataIn1 = 32'd1862
; 
32'd118842: dataIn1 = 32'd10524
; 
32'd118843: dataIn1 = 32'd10525
; 
32'd118844: dataIn1 = 32'd208
; 
32'd118845: dataIn1 = 32'd1484
; 
32'd118846: dataIn1 = 32'd1495
; 
32'd118847: dataIn1 = 32'd1860
; 
32'd118848: dataIn1 = 32'd1864
; 
32'd118849: dataIn1 = 32'd10516
; 
32'd118850: dataIn1 = 32'd10517
; 
32'd118851: dataIn1 = 32'd209
; 
32'd118852: dataIn1 = 32'd2529
; 
32'd118853: dataIn1 = 32'd2530
; 
32'd118854: dataIn1 = 32'd5890
; 
32'd118855: dataIn1 = 32'd5891
; 
32'd118856: dataIn1 = 32'd5920
; 
32'd118857: dataIn1 = 32'd5930
; 
32'd118858: dataIn1 = 32'd210
; 
32'd118859: dataIn1 = 32'd1498
; 
32'd118860: dataIn1 = 32'd1511
; 
32'd118861: dataIn1 = 32'd1866
; 
32'd118862: dataIn1 = 32'd1876
; 
32'd118863: dataIn1 = 32'd10508
; 
32'd118864: dataIn1 = 32'd10509
; 
32'd118865: dataIn1 = 32'd211
; 
32'd118866: dataIn1 = 32'd1501
; 
32'd118867: dataIn1 = 32'd1508
; 
32'd118868: dataIn1 = 32'd3444
; 
32'd118869: dataIn1 = 32'd10262
; 
32'd118870: dataIn1 = 32'd10500
; 
32'd118871: dataIn1 = 32'd10501
; 
32'd118872: dataIn1 = 32'd212
; 
32'd118873: dataIn1 = 32'd1043
; 
32'd118874: dataIn1 = 32'd2565
; 
32'd118875: dataIn1 = 32'd5428
; 
32'd118876: dataIn1 = 32'd5429
; 
32'd118877: dataIn1 = 32'd5511
; 
32'd118878: dataIn1 = 32'd10275
; 
32'd118879: dataIn1 = 32'd213
; 
32'd118880: dataIn1 = 32'd1505
; 
32'd118881: dataIn1 = 32'd1525
; 
32'd118882: dataIn1 = 32'd1870
; 
32'd118883: dataIn1 = 32'd1879
; 
32'd118884: dataIn1 = 32'd10492
; 
32'd118885: dataIn1 = 32'd10493
; 
32'd118886: dataIn1 = 32'd214
; 
32'd118887: dataIn1 = 32'd1522
; 
32'd118888: dataIn1 = 32'd1531
; 
32'd118889: dataIn1 = 32'd1877
; 
32'd118890: dataIn1 = 32'd1881
; 
32'd118891: dataIn1 = 32'd10484
; 
32'd118892: dataIn1 = 32'd10485
; 
32'd118893: dataIn1 = 32'd215
; 
32'd118894: dataIn1 = 32'd986
; 
32'd118895: dataIn1 = 32'd987
; 
32'd118896: dataIn1 = 32'd1044
; 
32'd118897: dataIn1 = 32'd1045
; 
32'd118898: dataIn1 = 32'd2054
; 
32'd118899: dataIn1 = 32'd3456
; 
32'd118900: dataIn1 = 32'd3466
; 
32'd118901: dataIn1 = 32'd216
; 
32'd118902: dataIn1 = 32'd1534
; 
32'd118903: dataIn1 = 32'd1547
; 
32'd118904: dataIn1 = 32'd1883
; 
32'd118905: dataIn1 = 32'd1892
; 
32'd118906: dataIn1 = 32'd10476
; 
32'd118907: dataIn1 = 32'd10477
; 
32'd118908: dataIn1 = 32'd217
; 
32'd118909: dataIn1 = 32'd1537
; 
32'd118910: dataIn1 = 32'd1544
; 
32'd118911: dataIn1 = 32'd1886
; 
32'd118912: dataIn1 = 32'd1890
; 
32'd118913: dataIn1 = 32'd10468
; 
32'd118914: dataIn1 = 32'd10469
; 
32'd118915: dataIn1 = 32'd218
; 
32'd118916: dataIn1 = 32'd988
; 
32'd118917: dataIn1 = 32'd989
; 
32'd118918: dataIn1 = 32'd1046
; 
32'd118919: dataIn1 = 32'd1047
; 
32'd118920: dataIn1 = 32'd2057
; 
32'd118921: dataIn1 = 32'd3481
; 
32'd118922: dataIn1 = 32'd3485
; 
32'd118923: dataIn1 = 32'd219
; 
32'd118924: dataIn1 = 32'd1541
; 
32'd118925: dataIn1 = 32'd1557
; 
32'd118926: dataIn1 = 32'd1887
; 
32'd118927: dataIn1 = 32'd1895
; 
32'd118928: dataIn1 = 32'd10460
; 
32'd118929: dataIn1 = 32'd10461
; 
32'd118930: dataIn1 = 32'd220
; 
32'd118931: dataIn1 = 32'd1554
; 
32'd118932: dataIn1 = 32'd1563
; 
32'd118933: dataIn1 = 32'd1893
; 
32'd118934: dataIn1 = 32'd1897
; 
32'd118935: dataIn1 = 32'd10452
; 
32'd118936: dataIn1 = 32'd10453
; 
32'd118937: dataIn1 = 32'd221
; 
32'd118938: dataIn1 = 32'd994
; 
32'd118939: dataIn1 = 32'd995
; 
32'd118940: dataIn1 = 32'd1048
; 
32'd118941: dataIn1 = 32'd1049
; 
32'd118942: dataIn1 = 32'd2062
; 
32'd118943: dataIn1 = 32'd3497
; 
32'd118944: dataIn1 = 32'd3500
; 
32'd118945: dataIn1 = 32'd222
; 
32'd118946: dataIn1 = 32'd1566
; 
32'd118947: dataIn1 = 32'd1579
; 
32'd118948: dataIn1 = 32'd1899
; 
32'd118949: dataIn1 = 32'd1908
; 
32'd118950: dataIn1 = 32'd10444
; 
32'd118951: dataIn1 = 32'd10445
; 
32'd118952: dataIn1 = 32'd223
; 
32'd118953: dataIn1 = 32'd1569
; 
32'd118954: dataIn1 = 32'd1576
; 
32'd118955: dataIn1 = 32'd1902
; 
32'd118956: dataIn1 = 32'd1906
; 
32'd118957: dataIn1 = 32'd10436
; 
32'd118958: dataIn1 = 32'd10437
; 
32'd118959: dataIn1 = 32'd224
; 
32'd118960: dataIn1 = 32'd996
; 
32'd118961: dataIn1 = 32'd997
; 
32'd118962: dataIn1 = 32'd1050
; 
32'd118963: dataIn1 = 32'd1051
; 
32'd118964: dataIn1 = 32'd2065
; 
32'd118965: dataIn1 = 32'd3507
; 
32'd118966: dataIn1 = 32'd3509
; 
32'd118967: dataIn1 = 32'd225
; 
32'd118968: dataIn1 = 32'd1573
; 
32'd118969: dataIn1 = 32'd1589
; 
32'd118970: dataIn1 = 32'd1903
; 
32'd118971: dataIn1 = 32'd1911
; 
32'd118972: dataIn1 = 32'd10428
; 
32'd118973: dataIn1 = 32'd10429
; 
32'd118974: dataIn1 = 32'd226
; 
32'd118975: dataIn1 = 32'd1586
; 
32'd118976: dataIn1 = 32'd1595
; 
32'd118977: dataIn1 = 32'd1909
; 
32'd118978: dataIn1 = 32'd1913
; 
32'd118979: dataIn1 = 32'd10420
; 
32'd118980: dataIn1 = 32'd10421
; 
32'd118981: dataIn1 = 32'd227
; 
32'd118982: dataIn1 = 32'd1002
; 
32'd118983: dataIn1 = 32'd1003
; 
32'd118984: dataIn1 = 32'd1052
; 
32'd118985: dataIn1 = 32'd1053
; 
32'd118986: dataIn1 = 32'd2070
; 
32'd118987: dataIn1 = 32'd3515
; 
32'd118988: dataIn1 = 32'd3517
; 
32'd118989: dataIn1 = 32'd228
; 
32'd118990: dataIn1 = 32'd1598
; 
32'd118991: dataIn1 = 32'd1611
; 
32'd118992: dataIn1 = 32'd1915
; 
32'd118993: dataIn1 = 32'd1924
; 
32'd118994: dataIn1 = 32'd10412
; 
32'd118995: dataIn1 = 32'd10413
; 
32'd118996: dataIn1 = 32'd229
; 
32'd118997: dataIn1 = 32'd1601
; 
32'd118998: dataIn1 = 32'd1608
; 
32'd118999: dataIn1 = 32'd1918
; 
32'd119000: dataIn1 = 32'd1922
; 
32'd119001: dataIn1 = 32'd10404
; 
32'd119002: dataIn1 = 32'd10405
; 
32'd119003: dataIn1 = 32'd230
; 
32'd119004: dataIn1 = 32'd1004
; 
32'd119005: dataIn1 = 32'd1005
; 
32'd119006: dataIn1 = 32'd1054
; 
32'd119007: dataIn1 = 32'd1055
; 
32'd119008: dataIn1 = 32'd2073
; 
32'd119009: dataIn1 = 32'd3523
; 
32'd119010: dataIn1 = 32'd3525
; 
32'd119011: dataIn1 = 32'd231
; 
32'd119012: dataIn1 = 32'd1605
; 
32'd119013: dataIn1 = 32'd1621
; 
32'd119014: dataIn1 = 32'd1919
; 
32'd119015: dataIn1 = 32'd1927
; 
32'd119016: dataIn1 = 32'd10396
; 
32'd119017: dataIn1 = 32'd10397
; 
32'd119018: dataIn1 = 32'd232
; 
32'd119019: dataIn1 = 32'd1618
; 
32'd119020: dataIn1 = 32'd1627
; 
32'd119021: dataIn1 = 32'd1925
; 
32'd119022: dataIn1 = 32'd1929
; 
32'd119023: dataIn1 = 32'd10388
; 
32'd119024: dataIn1 = 32'd10389
; 
32'd119025: dataIn1 = 32'd233
; 
32'd119026: dataIn1 = 32'd1010
; 
32'd119027: dataIn1 = 32'd1011
; 
32'd119028: dataIn1 = 32'd1056
; 
32'd119029: dataIn1 = 32'd1057
; 
32'd119030: dataIn1 = 32'd2078
; 
32'd119031: dataIn1 = 32'd3531
; 
32'd119032: dataIn1 = 32'd3533
; 
32'd119033: dataIn1 = 32'd234
; 
32'd119034: dataIn1 = 32'd1630
; 
32'd119035: dataIn1 = 32'd1643
; 
32'd119036: dataIn1 = 32'd1931
; 
32'd119037: dataIn1 = 32'd1940
; 
32'd119038: dataIn1 = 32'd10380
; 
32'd119039: dataIn1 = 32'd10381
; 
32'd119040: dataIn1 = 32'd235
; 
32'd119041: dataIn1 = 32'd1633
; 
32'd119042: dataIn1 = 32'd1640
; 
32'd119043: dataIn1 = 32'd1934
; 
32'd119044: dataIn1 = 32'd1938
; 
32'd119045: dataIn1 = 32'd10372
; 
32'd119046: dataIn1 = 32'd10373
; 
32'd119047: dataIn1 = 32'd236
; 
32'd119048: dataIn1 = 32'd1012
; 
32'd119049: dataIn1 = 32'd1013
; 
32'd119050: dataIn1 = 32'd1058
; 
32'd119051: dataIn1 = 32'd1059
; 
32'd119052: dataIn1 = 32'd2081
; 
32'd119053: dataIn1 = 32'd3539
; 
32'd119054: dataIn1 = 32'd3541
; 
32'd119055: dataIn1 = 32'd237
; 
32'd119056: dataIn1 = 32'd1637
; 
32'd119057: dataIn1 = 32'd1653
; 
32'd119058: dataIn1 = 32'd1935
; 
32'd119059: dataIn1 = 32'd1943
; 
32'd119060: dataIn1 = 32'd10364
; 
32'd119061: dataIn1 = 32'd10365
; 
32'd119062: dataIn1 = 32'd238
; 
32'd119063: dataIn1 = 32'd1650
; 
32'd119064: dataIn1 = 32'd1659
; 
32'd119065: dataIn1 = 32'd1941
; 
32'd119066: dataIn1 = 32'd1945
; 
32'd119067: dataIn1 = 32'd10356
; 
32'd119068: dataIn1 = 32'd10357
; 
32'd119069: dataIn1 = 32'd239
; 
32'd119070: dataIn1 = 32'd1018
; 
32'd119071: dataIn1 = 32'd1019
; 
32'd119072: dataIn1 = 32'd1060
; 
32'd119073: dataIn1 = 32'd1061
; 
32'd119074: dataIn1 = 32'd2086
; 
32'd119075: dataIn1 = 32'd3547
; 
32'd119076: dataIn1 = 32'd3549
; 
32'd119077: dataIn1 = 32'd240
; 
32'd119078: dataIn1 = 32'd1662
; 
32'd119079: dataIn1 = 32'd1675
; 
32'd119080: dataIn1 = 32'd1947
; 
32'd119081: dataIn1 = 32'd1956
; 
32'd119082: dataIn1 = 32'd10348
; 
32'd119083: dataIn1 = 32'd10349
; 
32'd119084: dataIn1 = 32'd241
; 
32'd119085: dataIn1 = 32'd1665
; 
32'd119086: dataIn1 = 32'd1672
; 
32'd119087: dataIn1 = 32'd1950
; 
32'd119088: dataIn1 = 32'd1954
; 
32'd119089: dataIn1 = 32'd10340
; 
32'd119090: dataIn1 = 32'd10341
; 
32'd119091: dataIn1 = 32'd242
; 
32'd119092: dataIn1 = 32'd1020
; 
32'd119093: dataIn1 = 32'd1021
; 
32'd119094: dataIn1 = 32'd1062
; 
32'd119095: dataIn1 = 32'd1063
; 
32'd119096: dataIn1 = 32'd2089
; 
32'd119097: dataIn1 = 32'd3555
; 
32'd119098: dataIn1 = 32'd3557
; 
32'd119099: dataIn1 = 32'd243
; 
32'd119100: dataIn1 = 32'd1669
; 
32'd119101: dataIn1 = 32'd1685
; 
32'd119102: dataIn1 = 32'd1951
; 
32'd119103: dataIn1 = 32'd1959
; 
32'd119104: dataIn1 = 32'd10332
; 
32'd119105: dataIn1 = 32'd10333
; 
32'd119106: dataIn1 = 32'd244
; 
32'd119107: dataIn1 = 32'd1682
; 
32'd119108: dataIn1 = 32'd1691
; 
32'd119109: dataIn1 = 32'd1957
; 
32'd119110: dataIn1 = 32'd1961
; 
32'd119111: dataIn1 = 32'd10324
; 
32'd119112: dataIn1 = 32'd10325
; 
32'd119113: dataIn1 = 32'd245
; 
32'd119114: dataIn1 = 32'd1026
; 
32'd119115: dataIn1 = 32'd1027
; 
32'd119116: dataIn1 = 32'd1064
; 
32'd119117: dataIn1 = 32'd1065
; 
32'd119118: dataIn1 = 32'd2094
; 
32'd119119: dataIn1 = 32'd3563
; 
32'd119120: dataIn1 = 32'd3565
; 
32'd119121: dataIn1 = 32'd246
; 
32'd119122: dataIn1 = 32'd1694
; 
32'd119123: dataIn1 = 32'd1707
; 
32'd119124: dataIn1 = 32'd1963
; 
32'd119125: dataIn1 = 32'd1972
; 
32'd119126: dataIn1 = 32'd10315
; 
32'd119127: dataIn1 = 32'd10316
; 
32'd119128: dataIn1 = 32'd10317
; 
32'd119129: dataIn1 = 32'd247
; 
32'd119130: dataIn1 = 32'd1697
; 
32'd119131: dataIn1 = 32'd1704
; 
32'd119132: dataIn1 = 32'd1970
; 
32'd119133: dataIn1 = 32'd10307
; 
32'd119134: dataIn1 = 32'd10308
; 
32'd119135: dataIn1 = 32'd248
; 
32'd119136: dataIn1 = 32'd1028
; 
32'd119137: dataIn1 = 32'd1066
; 
32'd119138: dataIn1 = 32'd1067
; 
32'd119139: dataIn1 = 32'd2097
; 
32'd119140: dataIn1 = 32'd2098
; 
32'd119141: dataIn1 = 32'd3571
; 
32'd119142: dataIn1 = 32'd3573
; 
32'd119143: dataIn1 = 32'd249
; 
32'd119144: dataIn1 = 32'd1701
; 
32'd119145: dataIn1 = 32'd1717
; 
32'd119146: dataIn1 = 32'd1967
; 
32'd119147: dataIn1 = 32'd10300
; 
32'd119148: dataIn1 = 32'd10301
; 
32'd119149: dataIn1 = 32'd250
; 
32'd119150: dataIn1 = 32'd1714
; 
32'd119151: dataIn1 = 32'd1973
; 
32'd119152: dataIn1 = 32'd10292
; 
32'd119153: dataIn1 = 32'd10293
; 
32'd119154: dataIn1 = 32'd251
; 
32'd119155: dataIn1 = 32'd1145
; 
32'd119156: dataIn1 = 32'd1146
; 
32'd119157: dataIn1 = 32'd1151
; 
32'd119158: dataIn1 = 32'd1191
; 
32'd119159: dataIn1 = 32'd3554
; 
32'd119160: dataIn1 = 32'd3556
; 
32'd119161: dataIn1 = 32'd252
; 
32'd119162: dataIn1 = 32'd1147
; 
32'd119163: dataIn1 = 32'd1148
; 
32'd119164: dataIn1 = 32'd1150
; 
32'd119165: dataIn1 = 32'd1166
; 
32'd119166: dataIn1 = 32'd3562
; 
32'd119167: dataIn1 = 32'd3564
; 
32'd119168: dataIn1 = 32'd253
; 
32'd119169: dataIn1 = 32'd1154
; 
32'd119170: dataIn1 = 32'd1155
; 
32'd119171: dataIn1 = 32'd1159
; 
32'd119172: dataIn1 = 32'd1165
; 
32'd119173: dataIn1 = 32'd3570
; 
32'd119174: dataIn1 = 32'd3572
; 
32'd119175: dataIn1 = 32'd254
; 
32'd119176: dataIn1 = 32'd1156
; 
32'd119177: dataIn1 = 32'd1157
; 
32'd119178: dataIn1 = 32'd1158
; 
32'd119179: dataIn1 = 32'd1171
; 
32'd119180: dataIn1 = 32'd3577
; 
32'd119181: dataIn1 = 32'd3578
; 
32'd119182: dataIn1 = 32'd255
; 
32'd119183: dataIn1 = 32'd1172
; 
32'd119184: dataIn1 = 32'd1173
; 
32'd119185: dataIn1 = 32'd3581
; 
32'd119186: dataIn1 = 32'd3582
; 
32'd119187: dataIn1 = 32'd256
; 
32'd119188: dataIn1 = 32'd1178
; 
32'd119189: dataIn1 = 32'd1179
; 
32'd119190: dataIn1 = 32'd1184
; 
32'd119191: dataIn1 = 32'd1190
; 
32'd119192: dataIn1 = 32'd3546
; 
32'd119193: dataIn1 = 32'd3548
; 
32'd119194: dataIn1 = 32'd257
; 
32'd119195: dataIn1 = 32'd1180
; 
32'd119196: dataIn1 = 32'd1181
; 
32'd119197: dataIn1 = 32'd1182
; 
32'd119198: dataIn1 = 32'd1197
; 
32'd119199: dataIn1 = 32'd3538
; 
32'd119200: dataIn1 = 32'd3540
; 
32'd119201: dataIn1 = 32'd258
; 
32'd119202: dataIn1 = 32'd1195
; 
32'd119203: dataIn1 = 32'd1196
; 
32'd119204: dataIn1 = 32'd1204
; 
32'd119205: dataIn1 = 32'd1205
; 
32'd119206: dataIn1 = 32'd3530
; 
32'd119207: dataIn1 = 32'd3532
; 
32'd119208: dataIn1 = 32'd259
; 
32'd119209: dataIn1 = 32'd1202
; 
32'd119210: dataIn1 = 32'd1203
; 
32'd119211: dataIn1 = 32'd1207
; 
32'd119212: dataIn1 = 32'd1237
; 
32'd119213: dataIn1 = 32'd3522
; 
32'd119214: dataIn1 = 32'd3524
; 
32'd119215: dataIn1 = 32'd260
; 
32'd119216: dataIn1 = 32'd1210
; 
32'd119217: dataIn1 = 32'd1211
; 
32'd119218: dataIn1 = 32'd1216
; 
32'd119219: dataIn1 = 32'd1257
; 
32'd119220: dataIn1 = 32'd3478
; 
32'd119221: dataIn1 = 32'd3482
; 
32'd119222: dataIn1 = 32'd261
; 
32'd119223: dataIn1 = 32'd1212
; 
32'd119224: dataIn1 = 32'd1213
; 
32'd119225: dataIn1 = 32'd1215
; 
32'd119226: dataIn1 = 32'd1231
; 
32'd119227: dataIn1 = 32'd3494
; 
32'd119228: dataIn1 = 32'd3498
; 
32'd119229: dataIn1 = 32'd262
; 
32'd119230: dataIn1 = 32'd1219
; 
32'd119231: dataIn1 = 32'd1220
; 
32'd119232: dataIn1 = 32'd1224
; 
32'd119233: dataIn1 = 32'd1230
; 
32'd119234: dataIn1 = 32'd3506
; 
32'd119235: dataIn1 = 32'd3508
; 
32'd119236: dataIn1 = 32'd263
; 
32'd119237: dataIn1 = 32'd1221
; 
32'd119238: dataIn1 = 32'd1222
; 
32'd119239: dataIn1 = 32'd1223
; 
32'd119240: dataIn1 = 32'd1236
; 
32'd119241: dataIn1 = 32'd3514
; 
32'd119242: dataIn1 = 32'd3516
; 
32'd119243: dataIn1 = 32'd264
; 
32'd119244: dataIn1 = 32'd1242
; 
32'd119245: dataIn1 = 32'd1243
; 
32'd119246: dataIn1 = 32'd1250
; 
32'd119247: dataIn1 = 32'd1256
; 
32'd119248: dataIn1 = 32'd3438
; 
32'd119249: dataIn1 = 32'd3458
; 
32'd119250: dataIn1 = 32'd265
; 
32'd119251: dataIn1 = 32'd1244
; 
32'd119252: dataIn1 = 32'd1245
; 
32'd119253: dataIn1 = 32'd1246
; 
32'd119254: dataIn1 = 32'd1260
; 
32'd119255: dataIn1 = 32'd2480
; 
32'd119256: dataIn1 = 32'd2481
; 
32'd119257: dataIn1 = 32'd266
; 
32'd119258: dataIn1 = 32'd548
; 
32'd119259: dataIn1 = 32'd549
; 
32'd119260: dataIn1 = 32'd750
; 
32'd119261: dataIn1 = 32'd958
; 
32'd119262: dataIn1 = 32'd959
; 
32'd119263: dataIn1 = 32'd2042
; 
32'd119264: dataIn1 = 32'd2756
; 
32'd119265: dataIn1 = 32'd10269
; 
32'd119266: dataIn1 = 32'd267
; 
32'd119267: dataIn1 = 32'd1259
; 
32'd119268: dataIn1 = 32'd1266
; 
32'd119269: dataIn1 = 32'd10249
; 
32'd119270: dataIn1 = 32'd10654
; 
32'd119271: dataIn1 = 32'd10655
; 
32'd119272: dataIn1 = 32'd10656
; 
32'd119273: dataIn1 = 32'd268
; 
32'd119274: dataIn1 = 32'd552
; 
32'd119275: dataIn1 = 32'd553
; 
32'd119276: dataIn1 = 32'd555
; 
32'd119277: dataIn1 = 32'd558
; 
32'd119278: dataIn1 = 32'd960
; 
32'd119279: dataIn1 = 32'd1270
; 
32'd119280: dataIn1 = 32'd3463
; 
32'd119281: dataIn1 = 32'd10255
; 
32'd119282: dataIn1 = 32'd269
; 
32'd119283: dataIn1 = 32'd551
; 
32'd119284: dataIn1 = 32'd552
; 
32'd119285: dataIn1 = 32'd554
; 
32'd119286: dataIn1 = 32'd559
; 
32'd119287: dataIn1 = 32'd1269
; 
32'd119288: dataIn1 = 32'd3471
; 
32'd119289: dataIn1 = 32'd3475
; 
32'd119290: dataIn1 = 32'd270
; 
32'd119291: dataIn1 = 32'd556
; 
32'd119292: dataIn1 = 32'd782
; 
32'd119293: dataIn1 = 32'd960
; 
32'd119294: dataIn1 = 32'd976
; 
32'd119295: dataIn1 = 32'd1271
; 
32'd119296: dataIn1 = 32'd1488
; 
32'd119297: dataIn1 = 32'd3450
; 
32'd119298: dataIn1 = 32'd10564
; 
32'd119299: dataIn1 = 32'd271
; 
32'd119300: dataIn1 = 32'd3424
; 
32'd119301: dataIn1 = 32'd3425
; 
32'd119302: dataIn1 = 32'd3451
; 
32'd119303: dataIn1 = 32'd3452
; 
32'd119304: dataIn1 = 32'd3475
; 
32'd119305: dataIn1 = 32'd3479
; 
32'd119306: dataIn1 = 32'd272
; 
32'd119307: dataIn1 = 32'd559
; 
32'd119308: dataIn1 = 32'd560
; 
32'd119309: dataIn1 = 32'd568
; 
32'd119310: dataIn1 = 32'd569
; 
32'd119311: dataIn1 = 32'd1287
; 
32'd119312: dataIn1 = 32'd3479
; 
32'd119313: dataIn1 = 32'd3483
; 
32'd119314: dataIn1 = 32'd273
; 
32'd119315: dataIn1 = 32'd1277
; 
32'd119316: dataIn1 = 32'd1278
; 
32'd119317: dataIn1 = 32'd1291
; 
32'd119318: dataIn1 = 32'd1292
; 
32'd119319: dataIn1 = 32'd1721
; 
32'd119320: dataIn1 = 32'd11600
; 
32'd119321: dataIn1 = 32'd274
; 
32'd119322: dataIn1 = 32'd561
; 
32'd119323: dataIn1 = 32'd562
; 
32'd119324: dataIn1 = 32'd563
; 
32'd119325: dataIn1 = 32'd567
; 
32'd119326: dataIn1 = 32'd1276
; 
32'd119327: dataIn1 = 32'd1279
; 
32'd119328: dataIn1 = 32'd1720
; 
32'd119329: dataIn1 = 32'd5526
; 
32'd119330: dataIn1 = 32'd275
; 
32'd119331: dataIn1 = 32'd566
; 
32'd119332: dataIn1 = 32'd567
; 
32'd119333: dataIn1 = 32'd1280
; 
32'd119334: dataIn1 = 32'd1281
; 
32'd119335: dataIn1 = 32'd1282
; 
32'd119336: dataIn1 = 32'd5525
; 
32'd119337: dataIn1 = 32'd276
; 
32'd119338: dataIn1 = 32'd5319
; 
32'd119339: dataIn1 = 32'd5320
; 
32'd119340: dataIn1 = 32'd5457
; 
32'd119341: dataIn1 = 32'd5525
; 
32'd119342: dataIn1 = 32'd5526
; 
32'd119343: dataIn1 = 32'd5527
; 
32'd119344: dataIn1 = 32'd277
; 
32'd119345: dataIn1 = 32'd569
; 
32'd119346: dataIn1 = 32'd570
; 
32'd119347: dataIn1 = 32'd571
; 
32'd119348: dataIn1 = 32'd3487
; 
32'd119349: dataIn1 = 32'd3491
; 
32'd119350: dataIn1 = 32'd3495
; 
32'd119351: dataIn1 = 32'd278
; 
32'd119352: dataIn1 = 32'd572
; 
32'd119353: dataIn1 = 32'd573
; 
32'd119354: dataIn1 = 32'd574
; 
32'd119355: dataIn1 = 32'd582
; 
32'd119356: dataIn1 = 32'd1290
; 
32'd119357: dataIn1 = 32'd1293
; 
32'd119358: dataIn1 = 32'd1722
; 
32'd119359: dataIn1 = 32'd5530
; 
32'd119360: dataIn1 = 32'd279
; 
32'd119361: dataIn1 = 32'd2764
; 
32'd119362: dataIn1 = 32'd2765
; 
32'd119363: dataIn1 = 32'd3044
; 
32'd119364: dataIn1 = 32'd3051
; 
32'd119365: dataIn1 = 32'd3989
; 
32'd119366: dataIn1 = 32'd3990
; 
32'd119367: dataIn1 = 32'd280
; 
32'd119368: dataIn1 = 32'd575
; 
32'd119369: dataIn1 = 32'd577
; 
32'd119370: dataIn1 = 32'd579
; 
32'd119371: dataIn1 = 32'd581
; 
32'd119372: dataIn1 = 32'd1296
; 
32'd119373: dataIn1 = 32'd5533
; 
32'd119374: dataIn1 = 32'd5534
; 
32'd119375: dataIn1 = 32'd281
; 
32'd119376: dataIn1 = 32'd575
; 
32'd119377: dataIn1 = 32'd576
; 
32'd119378: dataIn1 = 32'd578
; 
32'd119379: dataIn1 = 32'd582
; 
32'd119380: dataIn1 = 32'd1295
; 
32'd119381: dataIn1 = 32'd5531
; 
32'd119382: dataIn1 = 32'd5532
; 
32'd119383: dataIn1 = 32'd282
; 
32'd119384: dataIn1 = 32'd580
; 
32'd119385: dataIn1 = 32'd581
; 
32'd119386: dataIn1 = 32'd597
; 
32'd119387: dataIn1 = 32'd598
; 
32'd119388: dataIn1 = 32'd1308
; 
32'd119389: dataIn1 = 32'd5535
; 
32'd119390: dataIn1 = 32'd5536
; 
32'd119391: dataIn1 = 32'd283
; 
32'd119392: dataIn1 = 32'd5326
; 
32'd119393: dataIn1 = 32'd5327
; 
32'd119394: dataIn1 = 32'd5459
; 
32'd119395: dataIn1 = 32'd5460
; 
32'd119396: dataIn1 = 32'd5534
; 
32'd119397: dataIn1 = 32'd5535
; 
32'd119398: dataIn1 = 32'd284
; 
32'd119399: dataIn1 = 32'd5321
; 
32'd119400: dataIn1 = 32'd5322
; 
32'd119401: dataIn1 = 32'd5458
; 
32'd119402: dataIn1 = 32'd5529
; 
32'd119403: dataIn1 = 32'd5530
; 
32'd119404: dataIn1 = 32'd5531
; 
32'd119405: dataIn1 = 32'd285
; 
32'd119406: dataIn1 = 32'd2484
; 
32'd119407: dataIn1 = 32'd2485
; 
32'd119408: dataIn1 = 32'd2757
; 
32'd119409: dataIn1 = 32'd2769
; 
32'd119410: dataIn1 = 32'd3421
; 
32'd119411: dataIn1 = 32'd5304
; 
32'd119412: dataIn1 = 32'd286
; 
32'd119413: dataIn1 = 32'd2775
; 
32'd119414: dataIn1 = 32'd2776
; 
32'd119415: dataIn1 = 32'd3060
; 
32'd119416: dataIn1 = 32'd3066
; 
32'd119417: dataIn1 = 32'd4015
; 
32'd119418: dataIn1 = 32'd4016
; 
32'd119419: dataIn1 = 32'd287
; 
32'd119420: dataIn1 = 32'd588
; 
32'd119421: dataIn1 = 32'd589
; 
32'd119422: dataIn1 = 32'd591
; 
32'd119423: dataIn1 = 32'd593
; 
32'd119424: dataIn1 = 32'd1303
; 
32'd119425: dataIn1 = 32'd5541
; 
32'd119426: dataIn1 = 32'd5542
; 
32'd119427: dataIn1 = 32'd288
; 
32'd119428: dataIn1 = 32'd587
; 
32'd119429: dataIn1 = 32'd588
; 
32'd119430: dataIn1 = 32'd590
; 
32'd119431: dataIn1 = 32'd594
; 
32'd119432: dataIn1 = 32'd1302
; 
32'd119433: dataIn1 = 32'd5539
; 
32'd119434: dataIn1 = 32'd5540
; 
32'd119435: dataIn1 = 32'd289
; 
32'd119436: dataIn1 = 32'd592
; 
32'd119437: dataIn1 = 32'd593
; 
32'd119438: dataIn1 = 32'd599
; 
32'd119439: dataIn1 = 32'd601
; 
32'd119440: dataIn1 = 32'd1311
; 
32'd119441: dataIn1 = 32'd5543
; 
32'd119442: dataIn1 = 32'd5544
; 
32'd119443: dataIn1 = 32'd290
; 
32'd119444: dataIn1 = 32'd5334
; 
32'd119445: dataIn1 = 32'd5335
; 
32'd119446: dataIn1 = 32'd5463
; 
32'd119447: dataIn1 = 32'd5464
; 
32'd119448: dataIn1 = 32'd5542
; 
32'd119449: dataIn1 = 32'd5543
; 
32'd119450: dataIn1 = 32'd291
; 
32'd119451: dataIn1 = 32'd5330
; 
32'd119452: dataIn1 = 32'd5331
; 
32'd119453: dataIn1 = 32'd5461
; 
32'd119454: dataIn1 = 32'd5462
; 
32'd119455: dataIn1 = 32'd5538
; 
32'd119456: dataIn1 = 32'd5539
; 
32'd119457: dataIn1 = 32'd292
; 
32'd119458: dataIn1 = 32'd594
; 
32'd119459: dataIn1 = 32'd595
; 
32'd119460: dataIn1 = 32'd596
; 
32'd119461: dataIn1 = 32'd598
; 
32'd119462: dataIn1 = 32'd1307
; 
32'd119463: dataIn1 = 32'd5537
; 
32'd119464: dataIn1 = 32'd5538
; 
32'd119465: dataIn1 = 32'd293
; 
32'd119466: dataIn1 = 32'd2790
; 
32'd119467: dataIn1 = 32'd2791
; 
32'd119468: dataIn1 = 32'd3073
; 
32'd119469: dataIn1 = 32'd3081
; 
32'd119470: dataIn1 = 32'd4039
; 
32'd119471: dataIn1 = 32'd4040
; 
32'd119472: dataIn1 = 32'd294
; 
32'd119473: dataIn1 = 32'd599
; 
32'd119474: dataIn1 = 32'd600
; 
32'd119475: dataIn1 = 32'd602
; 
32'd119476: dataIn1 = 32'd610
; 
32'd119477: dataIn1 = 32'd1310
; 
32'd119478: dataIn1 = 32'd5545
; 
32'd119479: dataIn1 = 32'd5546
; 
32'd119480: dataIn1 = 32'd295
; 
32'd119481: dataIn1 = 32'd2795
; 
32'd119482: dataIn1 = 32'd2796
; 
32'd119483: dataIn1 = 32'd3086
; 
32'd119484: dataIn1 = 32'd3093
; 
32'd119485: dataIn1 = 32'd4085
; 
32'd119486: dataIn1 = 32'd4086
; 
32'd119487: dataIn1 = 32'd296
; 
32'd119488: dataIn1 = 32'd603
; 
32'd119489: dataIn1 = 32'd605
; 
32'd119490: dataIn1 = 32'd607
; 
32'd119491: dataIn1 = 32'd609
; 
32'd119492: dataIn1 = 32'd1314
; 
32'd119493: dataIn1 = 32'd5549
; 
32'd119494: dataIn1 = 32'd5550
; 
32'd119495: dataIn1 = 32'd297
; 
32'd119496: dataIn1 = 32'd603
; 
32'd119497: dataIn1 = 32'd604
; 
32'd119498: dataIn1 = 32'd606
; 
32'd119499: dataIn1 = 32'd610
; 
32'd119500: dataIn1 = 32'd1313
; 
32'd119501: dataIn1 = 32'd5547
; 
32'd119502: dataIn1 = 32'd5548
; 
32'd119503: dataIn1 = 32'd298
; 
32'd119504: dataIn1 = 32'd608
; 
32'd119505: dataIn1 = 32'd609
; 
32'd119506: dataIn1 = 32'd621
; 
32'd119507: dataIn1 = 32'd622
; 
32'd119508: dataIn1 = 32'd1324
; 
32'd119509: dataIn1 = 32'd5551
; 
32'd119510: dataIn1 = 32'd5552
; 
32'd119511: dataIn1 = 32'd299
; 
32'd119512: dataIn1 = 32'd5342
; 
32'd119513: dataIn1 = 32'd5343
; 
32'd119514: dataIn1 = 32'd5467
; 
32'd119515: dataIn1 = 32'd5468
; 
32'd119516: dataIn1 = 32'd5550
; 
32'd119517: dataIn1 = 32'd5551
; 
32'd119518: dataIn1 = 32'd300
; 
32'd119519: dataIn1 = 32'd5338
; 
32'd119520: dataIn1 = 32'd5339
; 
32'd119521: dataIn1 = 32'd5465
; 
32'd119522: dataIn1 = 32'd5466
; 
32'd119523: dataIn1 = 32'd5546
; 
32'd119524: dataIn1 = 32'd5547
; 
32'd119525: dataIn1 = 32'd301
; 
32'd119526: dataIn1 = 32'd2800
; 
32'd119527: dataIn1 = 32'd2801
; 
32'd119528: dataIn1 = 32'd3103
; 
32'd119529: dataIn1 = 32'd3110
; 
32'd119530: dataIn1 = 32'd4065
; 
32'd119531: dataIn1 = 32'd4066
; 
32'd119532: dataIn1 = 32'd302
; 
32'd119533: dataIn1 = 32'd2815
; 
32'd119534: dataIn1 = 32'd2816
; 
32'd119535: dataIn1 = 32'd3116
; 
32'd119536: dataIn1 = 32'd3122
; 
32'd119537: dataIn1 = 32'd4111
; 
32'd119538: dataIn1 = 32'd4112
; 
32'd119539: dataIn1 = 32'd303
; 
32'd119540: dataIn1 = 32'd612
; 
32'd119541: dataIn1 = 32'd613
; 
32'd119542: dataIn1 = 32'd615
; 
32'd119543: dataIn1 = 32'd617
; 
32'd119544: dataIn1 = 32'd1319
; 
32'd119545: dataIn1 = 32'd5557
; 
32'd119546: dataIn1 = 32'd5558
; 
32'd119547: dataIn1 = 32'd304
; 
32'd119548: dataIn1 = 32'd611
; 
32'd119549: dataIn1 = 32'd612
; 
32'd119550: dataIn1 = 32'd614
; 
32'd119551: dataIn1 = 32'd618
; 
32'd119552: dataIn1 = 32'd1318
; 
32'd119553: dataIn1 = 32'd5555
; 
32'd119554: dataIn1 = 32'd5556
; 
32'd119555: dataIn1 = 32'd305
; 
32'd119556: dataIn1 = 32'd616
; 
32'd119557: dataIn1 = 32'd617
; 
32'd119558: dataIn1 = 32'd623
; 
32'd119559: dataIn1 = 32'd625
; 
32'd119560: dataIn1 = 32'd1327
; 
32'd119561: dataIn1 = 32'd5559
; 
32'd119562: dataIn1 = 32'd5560
; 
32'd119563: dataIn1 = 32'd306
; 
32'd119564: dataIn1 = 32'd5350
; 
32'd119565: dataIn1 = 32'd5351
; 
32'd119566: dataIn1 = 32'd5471
; 
32'd119567: dataIn1 = 32'd5472
; 
32'd119568: dataIn1 = 32'd5558
; 
32'd119569: dataIn1 = 32'd5559
; 
32'd119570: dataIn1 = 32'd307
; 
32'd119571: dataIn1 = 32'd5346
; 
32'd119572: dataIn1 = 32'd5347
; 
32'd119573: dataIn1 = 32'd5469
; 
32'd119574: dataIn1 = 32'd5470
; 
32'd119575: dataIn1 = 32'd5554
; 
32'd119576: dataIn1 = 32'd5555
; 
32'd119577: dataIn1 = 32'd308
; 
32'd119578: dataIn1 = 32'd618
; 
32'd119579: dataIn1 = 32'd619
; 
32'd119580: dataIn1 = 32'd620
; 
32'd119581: dataIn1 = 32'd622
; 
32'd119582: dataIn1 = 32'd1323
; 
32'd119583: dataIn1 = 32'd5553
; 
32'd119584: dataIn1 = 32'd5554
; 
32'd119585: dataIn1 = 32'd309
; 
32'd119586: dataIn1 = 32'd2830
; 
32'd119587: dataIn1 = 32'd2831
; 
32'd119588: dataIn1 = 32'd3129
; 
32'd119589: dataIn1 = 32'd3137
; 
32'd119590: dataIn1 = 32'd4135
; 
32'd119591: dataIn1 = 32'd4136
; 
32'd119592: dataIn1 = 32'd310
; 
32'd119593: dataIn1 = 32'd623
; 
32'd119594: dataIn1 = 32'd624
; 
32'd119595: dataIn1 = 32'd626
; 
32'd119596: dataIn1 = 32'd634
; 
32'd119597: dataIn1 = 32'd1326
; 
32'd119598: dataIn1 = 32'd5561
; 
32'd119599: dataIn1 = 32'd5562
; 
32'd119600: dataIn1 = 32'd311
; 
32'd119601: dataIn1 = 32'd2835
; 
32'd119602: dataIn1 = 32'd2836
; 
32'd119603: dataIn1 = 32'd3142
; 
32'd119604: dataIn1 = 32'd3149
; 
32'd119605: dataIn1 = 32'd4181
; 
32'd119606: dataIn1 = 32'd4182
; 
32'd119607: dataIn1 = 32'd312
; 
32'd119608: dataIn1 = 32'd627
; 
32'd119609: dataIn1 = 32'd629
; 
32'd119610: dataIn1 = 32'd631
; 
32'd119611: dataIn1 = 32'd633
; 
32'd119612: dataIn1 = 32'd1330
; 
32'd119613: dataIn1 = 32'd5565
; 
32'd119614: dataIn1 = 32'd5566
; 
32'd119615: dataIn1 = 32'd313
; 
32'd119616: dataIn1 = 32'd627
; 
32'd119617: dataIn1 = 32'd628
; 
32'd119618: dataIn1 = 32'd630
; 
32'd119619: dataIn1 = 32'd634
; 
32'd119620: dataIn1 = 32'd1329
; 
32'd119621: dataIn1 = 32'd5563
; 
32'd119622: dataIn1 = 32'd5564
; 
32'd119623: dataIn1 = 32'd314
; 
32'd119624: dataIn1 = 32'd632
; 
32'd119625: dataIn1 = 32'd633
; 
32'd119626: dataIn1 = 32'd645
; 
32'd119627: dataIn1 = 32'd646
; 
32'd119628: dataIn1 = 32'd1340
; 
32'd119629: dataIn1 = 32'd5567
; 
32'd119630: dataIn1 = 32'd5568
; 
32'd119631: dataIn1 = 32'd315
; 
32'd119632: dataIn1 = 32'd5358
; 
32'd119633: dataIn1 = 32'd5359
; 
32'd119634: dataIn1 = 32'd5475
; 
32'd119635: dataIn1 = 32'd5476
; 
32'd119636: dataIn1 = 32'd5566
; 
32'd119637: dataIn1 = 32'd5567
; 
32'd119638: dataIn1 = 32'd316
; 
32'd119639: dataIn1 = 32'd5354
; 
32'd119640: dataIn1 = 32'd5355
; 
32'd119641: dataIn1 = 32'd5473
; 
32'd119642: dataIn1 = 32'd5474
; 
32'd119643: dataIn1 = 32'd5562
; 
32'd119644: dataIn1 = 32'd5563
; 
32'd119645: dataIn1 = 32'd317
; 
32'd119646: dataIn1 = 32'd2840
; 
32'd119647: dataIn1 = 32'd2841
; 
32'd119648: dataIn1 = 32'd3159
; 
32'd119649: dataIn1 = 32'd3166
; 
32'd119650: dataIn1 = 32'd4161
; 
32'd119651: dataIn1 = 32'd4162
; 
32'd119652: dataIn1 = 32'd318
; 
32'd119653: dataIn1 = 32'd2855
; 
32'd119654: dataIn1 = 32'd2856
; 
32'd119655: dataIn1 = 32'd3172
; 
32'd119656: dataIn1 = 32'd3178
; 
32'd119657: dataIn1 = 32'd4207
; 
32'd119658: dataIn1 = 32'd4208
; 
32'd119659: dataIn1 = 32'd319
; 
32'd119660: dataIn1 = 32'd636
; 
32'd119661: dataIn1 = 32'd637
; 
32'd119662: dataIn1 = 32'd639
; 
32'd119663: dataIn1 = 32'd641
; 
32'd119664: dataIn1 = 32'd1335
; 
32'd119665: dataIn1 = 32'd5573
; 
32'd119666: dataIn1 = 32'd5574
; 
32'd119667: dataIn1 = 32'd320
; 
32'd119668: dataIn1 = 32'd635
; 
32'd119669: dataIn1 = 32'd636
; 
32'd119670: dataIn1 = 32'd638
; 
32'd119671: dataIn1 = 32'd642
; 
32'd119672: dataIn1 = 32'd1334
; 
32'd119673: dataIn1 = 32'd5571
; 
32'd119674: dataIn1 = 32'd5572
; 
32'd119675: dataIn1 = 32'd321
; 
32'd119676: dataIn1 = 32'd640
; 
32'd119677: dataIn1 = 32'd641
; 
32'd119678: dataIn1 = 32'd647
; 
32'd119679: dataIn1 = 32'd649
; 
32'd119680: dataIn1 = 32'd1343
; 
32'd119681: dataIn1 = 32'd5575
; 
32'd119682: dataIn1 = 32'd5576
; 
32'd119683: dataIn1 = 32'd322
; 
32'd119684: dataIn1 = 32'd5366
; 
32'd119685: dataIn1 = 32'd5367
; 
32'd119686: dataIn1 = 32'd5479
; 
32'd119687: dataIn1 = 32'd5480
; 
32'd119688: dataIn1 = 32'd5574
; 
32'd119689: dataIn1 = 32'd5575
; 
32'd119690: dataIn1 = 32'd323
; 
32'd119691: dataIn1 = 32'd5362
; 
32'd119692: dataIn1 = 32'd5363
; 
32'd119693: dataIn1 = 32'd5477
; 
32'd119694: dataIn1 = 32'd5478
; 
32'd119695: dataIn1 = 32'd5570
; 
32'd119696: dataIn1 = 32'd5571
; 
32'd119697: dataIn1 = 32'd324
; 
32'd119698: dataIn1 = 32'd642
; 
32'd119699: dataIn1 = 32'd643
; 
32'd119700: dataIn1 = 32'd644
; 
32'd119701: dataIn1 = 32'd646
; 
32'd119702: dataIn1 = 32'd1339
; 
32'd119703: dataIn1 = 32'd5569
; 
32'd119704: dataIn1 = 32'd5570
; 
32'd119705: dataIn1 = 32'd325
; 
32'd119706: dataIn1 = 32'd2870
; 
32'd119707: dataIn1 = 32'd2871
; 
32'd119708: dataIn1 = 32'd3185
; 
32'd119709: dataIn1 = 32'd3193
; 
32'd119710: dataIn1 = 32'd4231
; 
32'd119711: dataIn1 = 32'd4232
; 
32'd119712: dataIn1 = 32'd326
; 
32'd119713: dataIn1 = 32'd647
; 
32'd119714: dataIn1 = 32'd648
; 
32'd119715: dataIn1 = 32'd650
; 
32'd119716: dataIn1 = 32'd658
; 
32'd119717: dataIn1 = 32'd1342
; 
32'd119718: dataIn1 = 32'd5577
; 
32'd119719: dataIn1 = 32'd5578
; 
32'd119720: dataIn1 = 32'd327
; 
32'd119721: dataIn1 = 32'd2875
; 
32'd119722: dataIn1 = 32'd2876
; 
32'd119723: dataIn1 = 32'd3198
; 
32'd119724: dataIn1 = 32'd3205
; 
32'd119725: dataIn1 = 32'd4277
; 
32'd119726: dataIn1 = 32'd4278
; 
32'd119727: dataIn1 = 32'd328
; 
32'd119728: dataIn1 = 32'd651
; 
32'd119729: dataIn1 = 32'd653
; 
32'd119730: dataIn1 = 32'd655
; 
32'd119731: dataIn1 = 32'd657
; 
32'd119732: dataIn1 = 32'd1346
; 
32'd119733: dataIn1 = 32'd5581
; 
32'd119734: dataIn1 = 32'd5582
; 
32'd119735: dataIn1 = 32'd329
; 
32'd119736: dataIn1 = 32'd651
; 
32'd119737: dataIn1 = 32'd652
; 
32'd119738: dataIn1 = 32'd654
; 
32'd119739: dataIn1 = 32'd658
; 
32'd119740: dataIn1 = 32'd1345
; 
32'd119741: dataIn1 = 32'd5579
; 
32'd119742: dataIn1 = 32'd5580
; 
32'd119743: dataIn1 = 32'd330
; 
32'd119744: dataIn1 = 32'd656
; 
32'd119745: dataIn1 = 32'd657
; 
32'd119746: dataIn1 = 32'd669
; 
32'd119747: dataIn1 = 32'd670
; 
32'd119748: dataIn1 = 32'd1356
; 
32'd119749: dataIn1 = 32'd5583
; 
32'd119750: dataIn1 = 32'd5584
; 
32'd119751: dataIn1 = 32'd331
; 
32'd119752: dataIn1 = 32'd5374
; 
32'd119753: dataIn1 = 32'd5375
; 
32'd119754: dataIn1 = 32'd5483
; 
32'd119755: dataIn1 = 32'd5484
; 
32'd119756: dataIn1 = 32'd5582
; 
32'd119757: dataIn1 = 32'd5583
; 
32'd119758: dataIn1 = 32'd332
; 
32'd119759: dataIn1 = 32'd5370
; 
32'd119760: dataIn1 = 32'd5371
; 
32'd119761: dataIn1 = 32'd5481
; 
32'd119762: dataIn1 = 32'd5482
; 
32'd119763: dataIn1 = 32'd5578
; 
32'd119764: dataIn1 = 32'd5579
; 
32'd119765: dataIn1 = 32'd333
; 
32'd119766: dataIn1 = 32'd2880
; 
32'd119767: dataIn1 = 32'd2881
; 
32'd119768: dataIn1 = 32'd3215
; 
32'd119769: dataIn1 = 32'd3222
; 
32'd119770: dataIn1 = 32'd4257
; 
32'd119771: dataIn1 = 32'd4258
; 
32'd119772: dataIn1 = 32'd334
; 
32'd119773: dataIn1 = 32'd2895
; 
32'd119774: dataIn1 = 32'd2896
; 
32'd119775: dataIn1 = 32'd3228
; 
32'd119776: dataIn1 = 32'd3234
; 
32'd119777: dataIn1 = 32'd4303
; 
32'd119778: dataIn1 = 32'd4304
; 
32'd119779: dataIn1 = 32'd335
; 
32'd119780: dataIn1 = 32'd660
; 
32'd119781: dataIn1 = 32'd661
; 
32'd119782: dataIn1 = 32'd663
; 
32'd119783: dataIn1 = 32'd665
; 
32'd119784: dataIn1 = 32'd1351
; 
32'd119785: dataIn1 = 32'd5589
; 
32'd119786: dataIn1 = 32'd5590
; 
32'd119787: dataIn1 = 32'd336
; 
32'd119788: dataIn1 = 32'd659
; 
32'd119789: dataIn1 = 32'd660
; 
32'd119790: dataIn1 = 32'd662
; 
32'd119791: dataIn1 = 32'd666
; 
32'd119792: dataIn1 = 32'd1350
; 
32'd119793: dataIn1 = 32'd5587
; 
32'd119794: dataIn1 = 32'd5588
; 
32'd119795: dataIn1 = 32'd337
; 
32'd119796: dataIn1 = 32'd664
; 
32'd119797: dataIn1 = 32'd665
; 
32'd119798: dataIn1 = 32'd671
; 
32'd119799: dataIn1 = 32'd673
; 
32'd119800: dataIn1 = 32'd1359
; 
32'd119801: dataIn1 = 32'd5591
; 
32'd119802: dataIn1 = 32'd5592
; 
32'd119803: dataIn1 = 32'd338
; 
32'd119804: dataIn1 = 32'd5382
; 
32'd119805: dataIn1 = 32'd5383
; 
32'd119806: dataIn1 = 32'd5487
; 
32'd119807: dataIn1 = 32'd5488
; 
32'd119808: dataIn1 = 32'd5590
; 
32'd119809: dataIn1 = 32'd5591
; 
32'd119810: dataIn1 = 32'd339
; 
32'd119811: dataIn1 = 32'd5378
; 
32'd119812: dataIn1 = 32'd5379
; 
32'd119813: dataIn1 = 32'd5485
; 
32'd119814: dataIn1 = 32'd5486
; 
32'd119815: dataIn1 = 32'd5586
; 
32'd119816: dataIn1 = 32'd5587
; 
32'd119817: dataIn1 = 32'd340
; 
32'd119818: dataIn1 = 32'd666
; 
32'd119819: dataIn1 = 32'd667
; 
32'd119820: dataIn1 = 32'd668
; 
32'd119821: dataIn1 = 32'd670
; 
32'd119822: dataIn1 = 32'd1355
; 
32'd119823: dataIn1 = 32'd5585
; 
32'd119824: dataIn1 = 32'd5586
; 
32'd119825: dataIn1 = 32'd341
; 
32'd119826: dataIn1 = 32'd2910
; 
32'd119827: dataIn1 = 32'd2911
; 
32'd119828: dataIn1 = 32'd3241
; 
32'd119829: dataIn1 = 32'd3249
; 
32'd119830: dataIn1 = 32'd4327
; 
32'd119831: dataIn1 = 32'd4328
; 
32'd119832: dataIn1 = 32'd342
; 
32'd119833: dataIn1 = 32'd671
; 
32'd119834: dataIn1 = 32'd672
; 
32'd119835: dataIn1 = 32'd674
; 
32'd119836: dataIn1 = 32'd682
; 
32'd119837: dataIn1 = 32'd1358
; 
32'd119838: dataIn1 = 32'd5593
; 
32'd119839: dataIn1 = 32'd5594
; 
32'd119840: dataIn1 = 32'd343
; 
32'd119841: dataIn1 = 32'd2915
; 
32'd119842: dataIn1 = 32'd2916
; 
32'd119843: dataIn1 = 32'd3254
; 
32'd119844: dataIn1 = 32'd3261
; 
32'd119845: dataIn1 = 32'd4373
; 
32'd119846: dataIn1 = 32'd4374
; 
32'd119847: dataIn1 = 32'd344
; 
32'd119848: dataIn1 = 32'd675
; 
32'd119849: dataIn1 = 32'd677
; 
32'd119850: dataIn1 = 32'd679
; 
32'd119851: dataIn1 = 32'd681
; 
32'd119852: dataIn1 = 32'd1362
; 
32'd119853: dataIn1 = 32'd5597
; 
32'd119854: dataIn1 = 32'd5598
; 
32'd119855: dataIn1 = 32'd345
; 
32'd119856: dataIn1 = 32'd675
; 
32'd119857: dataIn1 = 32'd676
; 
32'd119858: dataIn1 = 32'd678
; 
32'd119859: dataIn1 = 32'd682
; 
32'd119860: dataIn1 = 32'd1361
; 
32'd119861: dataIn1 = 32'd5595
; 
32'd119862: dataIn1 = 32'd5596
; 
32'd119863: dataIn1 = 32'd346
; 
32'd119864: dataIn1 = 32'd680
; 
32'd119865: dataIn1 = 32'd681
; 
32'd119866: dataIn1 = 32'd693
; 
32'd119867: dataIn1 = 32'd694
; 
32'd119868: dataIn1 = 32'd1372
; 
32'd119869: dataIn1 = 32'd5599
; 
32'd119870: dataIn1 = 32'd5600
; 
32'd119871: dataIn1 = 32'd347
; 
32'd119872: dataIn1 = 32'd5390
; 
32'd119873: dataIn1 = 32'd5391
; 
32'd119874: dataIn1 = 32'd5491
; 
32'd119875: dataIn1 = 32'd5492
; 
32'd119876: dataIn1 = 32'd5598
; 
32'd119877: dataIn1 = 32'd5599
; 
32'd119878: dataIn1 = 32'd348
; 
32'd119879: dataIn1 = 32'd5386
; 
32'd119880: dataIn1 = 32'd5387
; 
32'd119881: dataIn1 = 32'd5489
; 
32'd119882: dataIn1 = 32'd5490
; 
32'd119883: dataIn1 = 32'd5594
; 
32'd119884: dataIn1 = 32'd5595
; 
32'd119885: dataIn1 = 32'd349
; 
32'd119886: dataIn1 = 32'd2920
; 
32'd119887: dataIn1 = 32'd2921
; 
32'd119888: dataIn1 = 32'd3271
; 
32'd119889: dataIn1 = 32'd3278
; 
32'd119890: dataIn1 = 32'd4353
; 
32'd119891: dataIn1 = 32'd4354
; 
32'd119892: dataIn1 = 32'd350
; 
32'd119893: dataIn1 = 32'd2935
; 
32'd119894: dataIn1 = 32'd2936
; 
32'd119895: dataIn1 = 32'd3284
; 
32'd119896: dataIn1 = 32'd3290
; 
32'd119897: dataIn1 = 32'd4399
; 
32'd119898: dataIn1 = 32'd4400
; 
32'd119899: dataIn1 = 32'd351
; 
32'd119900: dataIn1 = 32'd684
; 
32'd119901: dataIn1 = 32'd685
; 
32'd119902: dataIn1 = 32'd687
; 
32'd119903: dataIn1 = 32'd689
; 
32'd119904: dataIn1 = 32'd1367
; 
32'd119905: dataIn1 = 32'd5605
; 
32'd119906: dataIn1 = 32'd5606
; 
32'd119907: dataIn1 = 32'd352
; 
32'd119908: dataIn1 = 32'd683
; 
32'd119909: dataIn1 = 32'd684
; 
32'd119910: dataIn1 = 32'd686
; 
32'd119911: dataIn1 = 32'd690
; 
32'd119912: dataIn1 = 32'd1366
; 
32'd119913: dataIn1 = 32'd5603
; 
32'd119914: dataIn1 = 32'd5604
; 
32'd119915: dataIn1 = 32'd353
; 
32'd119916: dataIn1 = 32'd688
; 
32'd119917: dataIn1 = 32'd689
; 
32'd119918: dataIn1 = 32'd695
; 
32'd119919: dataIn1 = 32'd697
; 
32'd119920: dataIn1 = 32'd1375
; 
32'd119921: dataIn1 = 32'd5607
; 
32'd119922: dataIn1 = 32'd5608
; 
32'd119923: dataIn1 = 32'd354
; 
32'd119924: dataIn1 = 32'd5398
; 
32'd119925: dataIn1 = 32'd5399
; 
32'd119926: dataIn1 = 32'd5495
; 
32'd119927: dataIn1 = 32'd5496
; 
32'd119928: dataIn1 = 32'd5606
; 
32'd119929: dataIn1 = 32'd5607
; 
32'd119930: dataIn1 = 32'd355
; 
32'd119931: dataIn1 = 32'd5394
; 
32'd119932: dataIn1 = 32'd5395
; 
32'd119933: dataIn1 = 32'd5493
; 
32'd119934: dataIn1 = 32'd5494
; 
32'd119935: dataIn1 = 32'd5602
; 
32'd119936: dataIn1 = 32'd5603
; 
32'd119937: dataIn1 = 32'd356
; 
32'd119938: dataIn1 = 32'd690
; 
32'd119939: dataIn1 = 32'd691
; 
32'd119940: dataIn1 = 32'd692
; 
32'd119941: dataIn1 = 32'd694
; 
32'd119942: dataIn1 = 32'd1371
; 
32'd119943: dataIn1 = 32'd5601
; 
32'd119944: dataIn1 = 32'd5602
; 
32'd119945: dataIn1 = 32'd357
; 
32'd119946: dataIn1 = 32'd2950
; 
32'd119947: dataIn1 = 32'd2951
; 
32'd119948: dataIn1 = 32'd3297
; 
32'd119949: dataIn1 = 32'd3305
; 
32'd119950: dataIn1 = 32'd4423
; 
32'd119951: dataIn1 = 32'd4424
; 
32'd119952: dataIn1 = 32'd358
; 
32'd119953: dataIn1 = 32'd695
; 
32'd119954: dataIn1 = 32'd696
; 
32'd119955: dataIn1 = 32'd698
; 
32'd119956: dataIn1 = 32'd706
; 
32'd119957: dataIn1 = 32'd1374
; 
32'd119958: dataIn1 = 32'd5609
; 
32'd119959: dataIn1 = 32'd5610
; 
32'd119960: dataIn1 = 32'd359
; 
32'd119961: dataIn1 = 32'd2955
; 
32'd119962: dataIn1 = 32'd2956
; 
32'd119963: dataIn1 = 32'd3310
; 
32'd119964: dataIn1 = 32'd3317
; 
32'd119965: dataIn1 = 32'd4469
; 
32'd119966: dataIn1 = 32'd4470
; 
32'd119967: dataIn1 = 32'd360
; 
32'd119968: dataIn1 = 32'd699
; 
32'd119969: dataIn1 = 32'd701
; 
32'd119970: dataIn1 = 32'd703
; 
32'd119971: dataIn1 = 32'd705
; 
32'd119972: dataIn1 = 32'd1378
; 
32'd119973: dataIn1 = 32'd5613
; 
32'd119974: dataIn1 = 32'd5614
; 
32'd119975: dataIn1 = 32'd361
; 
32'd119976: dataIn1 = 32'd699
; 
32'd119977: dataIn1 = 32'd700
; 
32'd119978: dataIn1 = 32'd702
; 
32'd119979: dataIn1 = 32'd706
; 
32'd119980: dataIn1 = 32'd1377
; 
32'd119981: dataIn1 = 32'd5611
; 
32'd119982: dataIn1 = 32'd5612
; 
32'd119983: dataIn1 = 32'd362
; 
32'd119984: dataIn1 = 32'd704
; 
32'd119985: dataIn1 = 32'd705
; 
32'd119986: dataIn1 = 32'd717
; 
32'd119987: dataIn1 = 32'd718
; 
32'd119988: dataIn1 = 32'd1388
; 
32'd119989: dataIn1 = 32'd5615
; 
32'd119990: dataIn1 = 32'd5616
; 
32'd119991: dataIn1 = 32'd363
; 
32'd119992: dataIn1 = 32'd5406
; 
32'd119993: dataIn1 = 32'd5407
; 
32'd119994: dataIn1 = 32'd5499
; 
32'd119995: dataIn1 = 32'd5500
; 
32'd119996: dataIn1 = 32'd5614
; 
32'd119997: dataIn1 = 32'd5615
; 
32'd119998: dataIn1 = 32'd364
; 
32'd119999: dataIn1 = 32'd5402
; 
32'd120000: dataIn1 = 32'd5403
; 
32'd120001: dataIn1 = 32'd5497
; 
32'd120002: dataIn1 = 32'd5498
; 
32'd120003: dataIn1 = 32'd5610
; 
32'd120004: dataIn1 = 32'd5611
; 
32'd120005: dataIn1 = 32'd365
; 
32'd120006: dataIn1 = 32'd2960
; 
32'd120007: dataIn1 = 32'd2961
; 
32'd120008: dataIn1 = 32'd3327
; 
32'd120009: dataIn1 = 32'd3334
; 
32'd120010: dataIn1 = 32'd4449
; 
32'd120011: dataIn1 = 32'd4450
; 
32'd120012: dataIn1 = 32'd366
; 
32'd120013: dataIn1 = 32'd2975
; 
32'd120014: dataIn1 = 32'd2976
; 
32'd120015: dataIn1 = 32'd3340
; 
32'd120016: dataIn1 = 32'd3346
; 
32'd120017: dataIn1 = 32'd4495
; 
32'd120018: dataIn1 = 32'd4496
; 
32'd120019: dataIn1 = 32'd367
; 
32'd120020: dataIn1 = 32'd708
; 
32'd120021: dataIn1 = 32'd709
; 
32'd120022: dataIn1 = 32'd711
; 
32'd120023: dataIn1 = 32'd713
; 
32'd120024: dataIn1 = 32'd1383
; 
32'd120025: dataIn1 = 32'd5621
; 
32'd120026: dataIn1 = 32'd5622
; 
32'd120027: dataIn1 = 32'd368
; 
32'd120028: dataIn1 = 32'd707
; 
32'd120029: dataIn1 = 32'd708
; 
32'd120030: dataIn1 = 32'd710
; 
32'd120031: dataIn1 = 32'd714
; 
32'd120032: dataIn1 = 32'd1382
; 
32'd120033: dataIn1 = 32'd5619
; 
32'd120034: dataIn1 = 32'd5620
; 
32'd120035: dataIn1 = 32'd369
; 
32'd120036: dataIn1 = 32'd712
; 
32'd120037: dataIn1 = 32'd713
; 
32'd120038: dataIn1 = 32'd719
; 
32'd120039: dataIn1 = 32'd721
; 
32'd120040: dataIn1 = 32'd1391
; 
32'd120041: dataIn1 = 32'd5623
; 
32'd120042: dataIn1 = 32'd5624
; 
32'd120043: dataIn1 = 32'd370
; 
32'd120044: dataIn1 = 32'd5414
; 
32'd120045: dataIn1 = 32'd5415
; 
32'd120046: dataIn1 = 32'd5503
; 
32'd120047: dataIn1 = 32'd5504
; 
32'd120048: dataIn1 = 32'd5622
; 
32'd120049: dataIn1 = 32'd5623
; 
32'd120050: dataIn1 = 32'd371
; 
32'd120051: dataIn1 = 32'd5410
; 
32'd120052: dataIn1 = 32'd5411
; 
32'd120053: dataIn1 = 32'd5501
; 
32'd120054: dataIn1 = 32'd5502
; 
32'd120055: dataIn1 = 32'd5618
; 
32'd120056: dataIn1 = 32'd5619
; 
32'd120057: dataIn1 = 32'd372
; 
32'd120058: dataIn1 = 32'd714
; 
32'd120059: dataIn1 = 32'd715
; 
32'd120060: dataIn1 = 32'd716
; 
32'd120061: dataIn1 = 32'd718
; 
32'd120062: dataIn1 = 32'd1387
; 
32'd120063: dataIn1 = 32'd5617
; 
32'd120064: dataIn1 = 32'd5618
; 
32'd120065: dataIn1 = 32'd373
; 
32'd120066: dataIn1 = 32'd2990
; 
32'd120067: dataIn1 = 32'd2991
; 
32'd120068: dataIn1 = 32'd3353
; 
32'd120069: dataIn1 = 32'd3361
; 
32'd120070: dataIn1 = 32'd4519
; 
32'd120071: dataIn1 = 32'd4520
; 
32'd120072: dataIn1 = 32'd374
; 
32'd120073: dataIn1 = 32'd719
; 
32'd120074: dataIn1 = 32'd720
; 
32'd120075: dataIn1 = 32'd722
; 
32'd120076: dataIn1 = 32'd730
; 
32'd120077: dataIn1 = 32'd1390
; 
32'd120078: dataIn1 = 32'd5625
; 
32'd120079: dataIn1 = 32'd5626
; 
32'd120080: dataIn1 = 32'd375
; 
32'd120081: dataIn1 = 32'd2995
; 
32'd120082: dataIn1 = 32'd2996
; 
32'd120083: dataIn1 = 32'd3366
; 
32'd120084: dataIn1 = 32'd3373
; 
32'd120085: dataIn1 = 32'd4565
; 
32'd120086: dataIn1 = 32'd4566
; 
32'd120087: dataIn1 = 32'd376
; 
32'd120088: dataIn1 = 32'd723
; 
32'd120089: dataIn1 = 32'd725
; 
32'd120090: dataIn1 = 32'd729
; 
32'd120091: dataIn1 = 32'd1392
; 
32'd120092: dataIn1 = 32'd1394
; 
32'd120093: dataIn1 = 32'd5629
; 
32'd120094: dataIn1 = 32'd5630
; 
32'd120095: dataIn1 = 32'd377
; 
32'd120096: dataIn1 = 32'd723
; 
32'd120097: dataIn1 = 32'd726
; 
32'd120098: dataIn1 = 32'd730
; 
32'd120099: dataIn1 = 32'd1393
; 
32'd120100: dataIn1 = 32'd1396
; 
32'd120101: dataIn1 = 32'd5627
; 
32'd120102: dataIn1 = 32'd5628
; 
32'd120103: dataIn1 = 32'd378
; 
32'd120104: dataIn1 = 32'd728
; 
32'd120105: dataIn1 = 32'd729
; 
32'd120106: dataIn1 = 32'd1395
; 
32'd120107: dataIn1 = 32'd5631
; 
32'd120108: dataIn1 = 32'd5632
; 
32'd120109: dataIn1 = 32'd379
; 
32'd120110: dataIn1 = 32'd5422
; 
32'd120111: dataIn1 = 32'd5423
; 
32'd120112: dataIn1 = 32'd5507
; 
32'd120113: dataIn1 = 32'd5508
; 
32'd120114: dataIn1 = 32'd5630
; 
32'd120115: dataIn1 = 32'd5631
; 
32'd120116: dataIn1 = 32'd380
; 
32'd120117: dataIn1 = 32'd5418
; 
32'd120118: dataIn1 = 32'd5419
; 
32'd120119: dataIn1 = 32'd5505
; 
32'd120120: dataIn1 = 32'd5506
; 
32'd120121: dataIn1 = 32'd5626
; 
32'd120122: dataIn1 = 32'd5627
; 
32'd120123: dataIn1 = 32'd381
; 
32'd120124: dataIn1 = 32'd3000
; 
32'd120125: dataIn1 = 32'd3001
; 
32'd120126: dataIn1 = 32'd3383
; 
32'd120127: dataIn1 = 32'd3390
; 
32'd120128: dataIn1 = 32'd4545
; 
32'd120129: dataIn1 = 32'd4546
; 
32'd120130: dataIn1 = 32'd382
; 
32'd120131: dataIn1 = 32'd3015
; 
32'd120132: dataIn1 = 32'd3016
; 
32'd120133: dataIn1 = 32'd3396
; 
32'd120134: dataIn1 = 32'd3402
; 
32'd120135: dataIn1 = 32'd4591
; 
32'd120136: dataIn1 = 32'd4592
; 
32'd120137: dataIn1 = 32'd383
; 
32'd120138: dataIn1 = 32'd1398
; 
32'd120139: dataIn1 = 32'd1399
; 
32'd120140: dataIn1 = 32'd1832
; 
32'd120141: dataIn1 = 32'd10748
; 
32'd120142: dataIn1 = 32'd10749
; 
32'd120143: dataIn1 = 32'd384
; 
32'd120144: dataIn1 = 32'd1402
; 
32'd120145: dataIn1 = 32'd1404
; 
32'd120146: dataIn1 = 32'd1833
; 
32'd120147: dataIn1 = 32'd10757
; 
32'd120148: dataIn1 = 32'd10758
; 
32'd120149: dataIn1 = 32'd385
; 
32'd120150: dataIn1 = 32'd1405
; 
32'd120151: dataIn1 = 32'd1407
; 
32'd120152: dataIn1 = 32'd1838
; 
32'd120153: dataIn1 = 32'd10740
; 
32'd120154: dataIn1 = 32'd10741
; 
32'd120155: dataIn1 = 32'd386
; 
32'd120156: dataIn1 = 32'd1409
; 
32'd120157: dataIn1 = 32'd1411
; 
32'd120158: dataIn1 = 32'd1842
; 
32'd120159: dataIn1 = 32'd1844
; 
32'd120160: dataIn1 = 32'd10732
; 
32'd120161: dataIn1 = 32'd10733
; 
32'd120162: dataIn1 = 32'd387
; 
32'd120163: dataIn1 = 32'd1414
; 
32'd120164: dataIn1 = 32'd1415
; 
32'd120165: dataIn1 = 32'd1845
; 
32'd120166: dataIn1 = 32'd1848
; 
32'd120167: dataIn1 = 32'd10716
; 
32'd120168: dataIn1 = 32'd10717
; 
32'd120169: dataIn1 = 32'd388
; 
32'd120170: dataIn1 = 32'd1418
; 
32'd120171: dataIn1 = 32'd1420
; 
32'd120172: dataIn1 = 32'd1849
; 
32'd120173: dataIn1 = 32'd1851
; 
32'd120174: dataIn1 = 32'd10724
; 
32'd120175: dataIn1 = 32'd10725
; 
32'd120176: dataIn1 = 32'd389
; 
32'd120177: dataIn1 = 32'd1425
; 
32'd120178: dataIn1 = 32'd1429
; 
32'd120179: dataIn1 = 32'd3442
; 
32'd120180: dataIn1 = 32'd10559
; 
32'd120181: dataIn1 = 32'd10560
; 
32'd120182: dataIn1 = 32'd10561
; 
32'd120183: dataIn1 = 32'd10708
; 
32'd120184: dataIn1 = 32'd10709
; 
32'd120185: dataIn1 = 32'd390
; 
32'd120186: dataIn1 = 32'd750
; 
32'd120187: dataIn1 = 32'd1421
; 
32'd120188: dataIn1 = 32'd1422
; 
32'd120189: dataIn1 = 32'd1423
; 
32'd120190: dataIn1 = 32'd2041
; 
32'd120191: dataIn1 = 32'd3470
; 
32'd120192: dataIn1 = 32'd391
; 
32'd120193: dataIn1 = 32'd3030
; 
32'd120194: dataIn1 = 32'd3031
; 
32'd120195: dataIn1 = 32'd3408
; 
32'd120196: dataIn1 = 32'd4611
; 
32'd120197: dataIn1 = 32'd4612
; 
32'd120198: dataIn1 = 32'd10257
; 
32'd120199: dataIn1 = 32'd392
; 
32'd120200: dataIn1 = 32'd748
; 
32'd120201: dataIn1 = 32'd749
; 
32'd120202: dataIn1 = 32'd761
; 
32'd120203: dataIn1 = 32'd1428
; 
32'd120204: dataIn1 = 32'd1855
; 
32'd120205: dataIn1 = 32'd2286
; 
32'd120206: dataIn1 = 32'd2289
; 
32'd120207: dataIn1 = 32'd10271
; 
32'd120208: dataIn1 = 32'd10272
; 
32'd120209: dataIn1 = 32'd393
; 
32'd120210: dataIn1 = 32'd1856
; 
32'd120211: dataIn1 = 32'd1857
; 
32'd120212: dataIn1 = 32'd1858
; 
32'd120213: dataIn1 = 32'd1859
; 
32'd120214: dataIn1 = 32'd2041
; 
32'd120215: dataIn1 = 32'd2042
; 
32'd120216: dataIn1 = 32'd3034
; 
32'd120217: dataIn1 = 32'd10270
; 
32'd120218: dataIn1 = 32'd394
; 
32'd120219: dataIn1 = 32'd1439
; 
32'd120220: dataIn1 = 32'd1445
; 
32'd120221: dataIn1 = 32'd3412
; 
32'd120222: dataIn1 = 32'd3413
; 
32'd120223: dataIn1 = 32'd10544
; 
32'd120224: dataIn1 = 32'd10545
; 
32'd120225: dataIn1 = 32'd10546
; 
32'd120226: dataIn1 = 32'd395
; 
32'd120227: dataIn1 = 32'd751
; 
32'd120228: dataIn1 = 32'd753
; 
32'd120229: dataIn1 = 32'd756
; 
32'd120230: dataIn1 = 32'd760
; 
32'd120231: dataIn1 = 32'd1443
; 
32'd120232: dataIn1 = 32'd5426
; 
32'd120233: dataIn1 = 32'd5509
; 
32'd120234: dataIn1 = 32'd396
; 
32'd120235: dataIn1 = 32'd751
; 
32'd120236: dataIn1 = 32'd752
; 
32'd120237: dataIn1 = 32'd754
; 
32'd120238: dataIn1 = 32'd761
; 
32'd120239: dataIn1 = 32'd1438
; 
32'd120240: dataIn1 = 32'd2489
; 
32'd120241: dataIn1 = 32'd4602
; 
32'd120242: dataIn1 = 32'd397
; 
32'd120243: dataIn1 = 32'd1466
; 
32'd120244: dataIn1 = 32'd1470
; 
32'd120245: dataIn1 = 32'd1471
; 
32'd120246: dataIn1 = 32'd3469
; 
32'd120247: dataIn1 = 32'd10259
; 
32'd120248: dataIn1 = 32'd10671
; 
32'd120249: dataIn1 = 32'd398
; 
32'd120250: dataIn1 = 32'd759
; 
32'd120251: dataIn1 = 32'd760
; 
32'd120252: dataIn1 = 32'd773
; 
32'd120253: dataIn1 = 32'd774
; 
32'd120254: dataIn1 = 32'd1478
; 
32'd120255: dataIn1 = 32'd5427
; 
32'd120256: dataIn1 = 32'd5510
; 
32'd120257: dataIn1 = 32'd399
; 
32'd120258: dataIn1 = 32'd3887
; 
32'd120259: dataIn1 = 32'd3888
; 
32'd120260: dataIn1 = 32'd3890
; 
32'd120261: dataIn1 = 32'd3891
; 
32'd120262: dataIn1 = 32'd5509
; 
32'd120263: dataIn1 = 32'd5510
; 
32'd120264: dataIn1 = 32'd400
; 
32'd120265: dataIn1 = 32'd2289
; 
32'd120266: dataIn1 = 32'd2489
; 
32'd120267: dataIn1 = 32'd3897
; 
32'd120268: dataIn1 = 32'd5682
; 
32'd120269: dataIn1 = 32'd5683
; 
32'd120270: dataIn1 = 32'd5692
; 
32'd120271: dataIn1 = 32'd401
; 
32'd120272: dataIn1 = 32'd763
; 
32'd120273: dataIn1 = 32'd764
; 
32'd120274: dataIn1 = 32'd767
; 
32'd120275: dataIn1 = 32'd2045
; 
32'd120276: dataIn1 = 32'd2291
; 
32'd120277: dataIn1 = 32'd2524
; 
32'd120278: dataIn1 = 32'd402
; 
32'd120279: dataIn1 = 32'd1458
; 
32'd120280: dataIn1 = 32'd1460
; 
32'd120281: dataIn1 = 32'd10530
; 
32'd120282: dataIn1 = 32'd10531
; 
32'd120283: dataIn1 = 32'd10532
; 
32'd120284: dataIn1 = 32'd10679
; 
32'd120285: dataIn1 = 32'd10680
; 
32'd120286: dataIn1 = 32'd10681
; 
32'd120287: dataIn1 = 32'd403
; 
32'd120288: dataIn1 = 32'd762
; 
32'd120289: dataIn1 = 32'd763
; 
32'd120290: dataIn1 = 32'd765
; 
32'd120291: dataIn1 = 32'd769
; 
32'd120292: dataIn1 = 32'd1456
; 
32'd120293: dataIn1 = 32'd2290
; 
32'd120294: dataIn1 = 32'd2292
; 
32'd120295: dataIn1 = 32'd404
; 
32'd120296: dataIn1 = 32'd2292
; 
32'd120297: dataIn1 = 32'd2293
; 
32'd120298: dataIn1 = 32'd2490
; 
32'd120299: dataIn1 = 32'd3922
; 
32'd120300: dataIn1 = 32'd3923
; 
32'd120301: dataIn1 = 32'd3926
; 
32'd120302: dataIn1 = 32'd5745
; 
32'd120303: dataIn1 = 32'd405
; 
32'd120304: dataIn1 = 32'd769
; 
32'd120305: dataIn1 = 32'd770
; 
32'd120306: dataIn1 = 32'd772
; 
32'd120307: dataIn1 = 32'd774
; 
32'd120308: dataIn1 = 32'd1476
; 
32'd120309: dataIn1 = 32'd2490
; 
32'd120310: dataIn1 = 32'd4603
; 
32'd120311: dataIn1 = 32'd406
; 
32'd120312: dataIn1 = 32'd1483
; 
32'd120313: dataIn1 = 32'd1486
; 
32'd120314: dataIn1 = 32'd1861
; 
32'd120315: dataIn1 = 32'd1863
; 
32'd120316: dataIn1 = 32'd10520
; 
32'd120317: dataIn1 = 32'd10521
; 
32'd120318: dataIn1 = 32'd407
; 
32'd120319: dataIn1 = 32'd976
; 
32'd120320: dataIn1 = 32'd2491
; 
32'd120321: dataIn1 = 32'd2493
; 
32'd120322: dataIn1 = 32'd2497
; 
32'd120323: dataIn1 = 32'd2499
; 
32'd120324: dataIn1 = 32'd3423
; 
32'd120325: dataIn1 = 32'd408
; 
32'd120326: dataIn1 = 32'd2494
; 
32'd120327: dataIn1 = 32'd2495
; 
32'd120328: dataIn1 = 32'd2503
; 
32'd120329: dataIn1 = 32'd2504
; 
32'd120330: dataIn1 = 32'd3422
; 
32'd120331: dataIn1 = 32'd3424
; 
32'd120332: dataIn1 = 32'd409
; 
32'd120333: dataIn1 = 32'd2501
; 
32'd120334: dataIn1 = 32'd2502
; 
32'd120335: dataIn1 = 32'd2509
; 
32'd120336: dataIn1 = 32'd2510
; 
32'd120337: dataIn1 = 32'd3425
; 
32'd120338: dataIn1 = 32'd3426
; 
32'd120339: dataIn1 = 32'd410
; 
32'd120340: dataIn1 = 32'd1494
; 
32'd120341: dataIn1 = 32'd1497
; 
32'd120342: dataIn1 = 32'd1865
; 
32'd120343: dataIn1 = 32'd1867
; 
32'd120344: dataIn1 = 32'd10512
; 
32'd120345: dataIn1 = 32'd10513
; 
32'd120346: dataIn1 = 32'd411
; 
32'd120347: dataIn1 = 32'd2506
; 
32'd120348: dataIn1 = 32'd2508
; 
32'd120349: dataIn1 = 32'd2518
; 
32'd120350: dataIn1 = 32'd2519
; 
32'd120351: dataIn1 = 32'd3427
; 
32'd120352: dataIn1 = 32'd3428
; 
32'd120353: dataIn1 = 32'd412
; 
32'd120354: dataIn1 = 32'd1502
; 
32'd120355: dataIn1 = 32'd1504
; 
32'd120356: dataIn1 = 32'd1871
; 
32'd120357: dataIn1 = 32'd3443
; 
32'd120358: dataIn1 = 32'd10496
; 
32'd120359: dataIn1 = 32'd10497
; 
32'd120360: dataIn1 = 32'd413
; 
32'd120361: dataIn1 = 32'd2513
; 
32'd120362: dataIn1 = 32'd2514
; 
32'd120363: dataIn1 = 32'd2516
; 
32'd120364: dataIn1 = 32'd2517
; 
32'd120365: dataIn1 = 32'd3429
; 
32'd120366: dataIn1 = 32'd10264
; 
32'd120367: dataIn1 = 32'd414
; 
32'd120368: dataIn1 = 32'd1514
; 
32'd120369: dataIn1 = 32'd1517
; 
32'd120370: dataIn1 = 32'd1872
; 
32'd120371: dataIn1 = 32'd3040
; 
32'd120372: dataIn1 = 32'd3440
; 
32'd120373: dataIn1 = 32'd10973
; 
32'd120374: dataIn1 = 32'd10974
; 
32'd120375: dataIn1 = 32'd415
; 
32'd120376: dataIn1 = 32'd1509
; 
32'd120377: dataIn1 = 32'd1512
; 
32'd120378: dataIn1 = 32'd1873
; 
32'd120379: dataIn1 = 32'd1875
; 
32'd120380: dataIn1 = 32'd10504
; 
32'd120381: dataIn1 = 32'd10505
; 
32'd120382: dataIn1 = 32'd416
; 
32'd120383: dataIn1 = 32'd3428
; 
32'd120384: dataIn1 = 32'd3429
; 
32'd120385: dataIn1 = 32'd3453
; 
32'd120386: dataIn1 = 32'd3454
; 
32'd120387: dataIn1 = 32'd3464
; 
32'd120388: dataIn1 = 32'd3491
; 
32'd120389: dataIn1 = 32'd417
; 
32'd120390: dataIn1 = 32'd1521
; 
32'd120391: dataIn1 = 32'd1524
; 
32'd120392: dataIn1 = 32'd1878
; 
32'd120393: dataIn1 = 32'd1880
; 
32'd120394: dataIn1 = 32'd10488
; 
32'd120395: dataIn1 = 32'd10489
; 
32'd120396: dataIn1 = 32'd418
; 
32'd120397: dataIn1 = 32'd1530
; 
32'd120398: dataIn1 = 32'd1533
; 
32'd120399: dataIn1 = 32'd1882
; 
32'd120400: dataIn1 = 32'd1884
; 
32'd120401: dataIn1 = 32'd10480
; 
32'd120402: dataIn1 = 32'd10481
; 
32'd120403: dataIn1 = 32'd419
; 
32'd120404: dataIn1 = 32'd1538
; 
32'd120405: dataIn1 = 32'd1540
; 
32'd120406: dataIn1 = 32'd1885
; 
32'd120407: dataIn1 = 32'd1888
; 
32'd120408: dataIn1 = 32'd10464
; 
32'd120409: dataIn1 = 32'd10465
; 
32'd120410: dataIn1 = 32'd420
; 
32'd120411: dataIn1 = 32'd1545
; 
32'd120412: dataIn1 = 32'd1548
; 
32'd120413: dataIn1 = 32'd1889
; 
32'd120414: dataIn1 = 32'd1891
; 
32'd120415: dataIn1 = 32'd10472
; 
32'd120416: dataIn1 = 32'd10473
; 
32'd120417: dataIn1 = 32'd421
; 
32'd120418: dataIn1 = 32'd1553
; 
32'd120419: dataIn1 = 32'd1556
; 
32'd120420: dataIn1 = 32'd1894
; 
32'd120421: dataIn1 = 32'd1896
; 
32'd120422: dataIn1 = 32'd10456
; 
32'd120423: dataIn1 = 32'd10457
; 
32'd120424: dataIn1 = 32'd422
; 
32'd120425: dataIn1 = 32'd1562
; 
32'd120426: dataIn1 = 32'd1565
; 
32'd120427: dataIn1 = 32'd1898
; 
32'd120428: dataIn1 = 32'd1900
; 
32'd120429: dataIn1 = 32'd10448
; 
32'd120430: dataIn1 = 32'd10449
; 
32'd120431: dataIn1 = 32'd423
; 
32'd120432: dataIn1 = 32'd1570
; 
32'd120433: dataIn1 = 32'd1572
; 
32'd120434: dataIn1 = 32'd1901
; 
32'd120435: dataIn1 = 32'd1904
; 
32'd120436: dataIn1 = 32'd10432
; 
32'd120437: dataIn1 = 32'd10433
; 
32'd120438: dataIn1 = 32'd424
; 
32'd120439: dataIn1 = 32'd1577
; 
32'd120440: dataIn1 = 32'd1580
; 
32'd120441: dataIn1 = 32'd1905
; 
32'd120442: dataIn1 = 32'd1907
; 
32'd120443: dataIn1 = 32'd10440
; 
32'd120444: dataIn1 = 32'd10441
; 
32'd120445: dataIn1 = 32'd425
; 
32'd120446: dataIn1 = 32'd1585
; 
32'd120447: dataIn1 = 32'd1588
; 
32'd120448: dataIn1 = 32'd1910
; 
32'd120449: dataIn1 = 32'd1912
; 
32'd120450: dataIn1 = 32'd10424
; 
32'd120451: dataIn1 = 32'd10425
; 
32'd120452: dataIn1 = 32'd426
; 
32'd120453: dataIn1 = 32'd1594
; 
32'd120454: dataIn1 = 32'd1597
; 
32'd120455: dataIn1 = 32'd1914
; 
32'd120456: dataIn1 = 32'd1916
; 
32'd120457: dataIn1 = 32'd10416
; 
32'd120458: dataIn1 = 32'd10417
; 
32'd120459: dataIn1 = 32'd427
; 
32'd120460: dataIn1 = 32'd1602
; 
32'd120461: dataIn1 = 32'd1604
; 
32'd120462: dataIn1 = 32'd1917
; 
32'd120463: dataIn1 = 32'd1920
; 
32'd120464: dataIn1 = 32'd10400
; 
32'd120465: dataIn1 = 32'd10401
; 
32'd120466: dataIn1 = 32'd428
; 
32'd120467: dataIn1 = 32'd1609
; 
32'd120468: dataIn1 = 32'd1612
; 
32'd120469: dataIn1 = 32'd1921
; 
32'd120470: dataIn1 = 32'd1923
; 
32'd120471: dataIn1 = 32'd10408
; 
32'd120472: dataIn1 = 32'd10409
; 
32'd120473: dataIn1 = 32'd429
; 
32'd120474: dataIn1 = 32'd1617
; 
32'd120475: dataIn1 = 32'd1620
; 
32'd120476: dataIn1 = 32'd1926
; 
32'd120477: dataIn1 = 32'd1928
; 
32'd120478: dataIn1 = 32'd10392
; 
32'd120479: dataIn1 = 32'd10393
; 
32'd120480: dataIn1 = 32'd430
; 
32'd120481: dataIn1 = 32'd1626
; 
32'd120482: dataIn1 = 32'd1629
; 
32'd120483: dataIn1 = 32'd1930
; 
32'd120484: dataIn1 = 32'd1932
; 
32'd120485: dataIn1 = 32'd10384
; 
32'd120486: dataIn1 = 32'd10385
; 
32'd120487: dataIn1 = 32'd431
; 
32'd120488: dataIn1 = 32'd1634
; 
32'd120489: dataIn1 = 32'd1636
; 
32'd120490: dataIn1 = 32'd1933
; 
32'd120491: dataIn1 = 32'd1936
; 
32'd120492: dataIn1 = 32'd10368
; 
32'd120493: dataIn1 = 32'd10369
; 
32'd120494: dataIn1 = 32'd432
; 
32'd120495: dataIn1 = 32'd1641
; 
32'd120496: dataIn1 = 32'd1644
; 
32'd120497: dataIn1 = 32'd1937
; 
32'd120498: dataIn1 = 32'd1939
; 
32'd120499: dataIn1 = 32'd10376
; 
32'd120500: dataIn1 = 32'd10377
; 
32'd120501: dataIn1 = 32'd433
; 
32'd120502: dataIn1 = 32'd1649
; 
32'd120503: dataIn1 = 32'd1652
; 
32'd120504: dataIn1 = 32'd1942
; 
32'd120505: dataIn1 = 32'd1944
; 
32'd120506: dataIn1 = 32'd10360
; 
32'd120507: dataIn1 = 32'd10361
; 
32'd120508: dataIn1 = 32'd434
; 
32'd120509: dataIn1 = 32'd1658
; 
32'd120510: dataIn1 = 32'd1661
; 
32'd120511: dataIn1 = 32'd1946
; 
32'd120512: dataIn1 = 32'd1948
; 
32'd120513: dataIn1 = 32'd10352
; 
32'd120514: dataIn1 = 32'd10353
; 
32'd120515: dataIn1 = 32'd435
; 
32'd120516: dataIn1 = 32'd1666
; 
32'd120517: dataIn1 = 32'd1668
; 
32'd120518: dataIn1 = 32'd1949
; 
32'd120519: dataIn1 = 32'd1952
; 
32'd120520: dataIn1 = 32'd10336
; 
32'd120521: dataIn1 = 32'd10337
; 
32'd120522: dataIn1 = 32'd436
; 
32'd120523: dataIn1 = 32'd1673
; 
32'd120524: dataIn1 = 32'd1676
; 
32'd120525: dataIn1 = 32'd1953
; 
32'd120526: dataIn1 = 32'd1955
; 
32'd120527: dataIn1 = 32'd10344
; 
32'd120528: dataIn1 = 32'd10345
; 
32'd120529: dataIn1 = 32'd437
; 
32'd120530: dataIn1 = 32'd1681
; 
32'd120531: dataIn1 = 32'd1684
; 
32'd120532: dataIn1 = 32'd1958
; 
32'd120533: dataIn1 = 32'd1960
; 
32'd120534: dataIn1 = 32'd10328
; 
32'd120535: dataIn1 = 32'd10329
; 
32'd120536: dataIn1 = 32'd438
; 
32'd120537: dataIn1 = 32'd1690
; 
32'd120538: dataIn1 = 32'd1693
; 
32'd120539: dataIn1 = 32'd1962
; 
32'd120540: dataIn1 = 32'd1964
; 
32'd120541: dataIn1 = 32'd10320
; 
32'd120542: dataIn1 = 32'd10321
; 
32'd120543: dataIn1 = 32'd439
; 
32'd120544: dataIn1 = 32'd1698
; 
32'd120545: dataIn1 = 32'd1700
; 
32'd120546: dataIn1 = 32'd1965
; 
32'd120547: dataIn1 = 32'd10304
; 
32'd120548: dataIn1 = 32'd10305
; 
32'd120549: dataIn1 = 32'd440
; 
32'd120550: dataIn1 = 32'd1705
; 
32'd120551: dataIn1 = 32'd1708
; 
32'd120552: dataIn1 = 32'd1971
; 
32'd120553: dataIn1 = 32'd10312
; 
32'd120554: dataIn1 = 32'd441
; 
32'd120555: dataIn1 = 32'd1713
; 
32'd120556: dataIn1 = 32'd1716
; 
32'd120557: dataIn1 = 32'd1976
; 
32'd120558: dataIn1 = 32'd10296
; 
32'd120559: dataIn1 = 32'd10297
; 
32'd120560: dataIn1 = 32'd442
; 
32'd120561: dataIn1 = 32'd3420
; 
32'd120562: dataIn1 = 32'd3421
; 
32'd120563: dataIn1 = 32'd3449
; 
32'd120564: dataIn1 = 32'd3464
; 
32'd120565: dataIn1 = 32'd3495
; 
32'd120566: dataIn1 = 32'd3499
; 
32'd120567: dataIn1 = 32'd443
; 
32'd120568: dataIn1 = 32'd2294
; 
32'd120569: dataIn1 = 32'd2295
; 
32'd120570: dataIn1 = 32'd2310
; 
32'd120571: dataIn1 = 32'd3449
; 
32'd120572: dataIn1 = 32'd3502
; 
32'd120573: dataIn1 = 32'd3870
; 
32'd120574: dataIn1 = 32'd3929
; 
32'd120575: dataIn1 = 32'd5319
; 
32'd120576: dataIn1 = 32'd444
; 
32'd120577: dataIn1 = 32'd3876
; 
32'd120578: dataIn1 = 32'd3877
; 
32'd120579: dataIn1 = 32'd3885
; 
32'd120580: dataIn1 = 32'd3898
; 
32'd120581: dataIn1 = 32'd4823
; 
32'd120582: dataIn1 = 32'd4824
; 
32'd120583: dataIn1 = 32'd445
; 
32'd120584: dataIn1 = 32'd3878
; 
32'd120585: dataIn1 = 32'd3879
; 
32'd120586: dataIn1 = 32'd3886
; 
32'd120587: dataIn1 = 32'd3893
; 
32'd120588: dataIn1 = 32'd3941
; 
32'd120589: dataIn1 = 32'd3942
; 
32'd120590: dataIn1 = 32'd5674
; 
32'd120591: dataIn1 = 32'd446
; 
32'd120592: dataIn1 = 32'd3903
; 
32'd120593: dataIn1 = 32'd3904
; 
32'd120594: dataIn1 = 32'd3917
; 
32'd120595: dataIn1 = 32'd3924
; 
32'd120596: dataIn1 = 32'd3937
; 
32'd120597: dataIn1 = 32'd3938
; 
32'd120598: dataIn1 = 32'd5752
; 
32'd120599: dataIn1 = 32'd5814
; 
32'd120600: dataIn1 = 32'd447
; 
32'd120601: dataIn1 = 32'd3907
; 
32'd120602: dataIn1 = 32'd3908
; 
32'd120603: dataIn1 = 32'd3913
; 
32'd120604: dataIn1 = 32'd3920
; 
32'd120605: dataIn1 = 32'd4865
; 
32'd120606: dataIn1 = 32'd4866
; 
32'd120607: dataIn1 = 32'd6700
; 
32'd120608: dataIn1 = 32'd6732
; 
32'd120609: dataIn1 = 32'd448
; 
32'd120610: dataIn1 = 32'd3930
; 
32'd120611: dataIn1 = 32'd3931
; 
32'd120612: dataIn1 = 32'd3959
; 
32'd120613: dataIn1 = 32'd5320
; 
32'd120614: dataIn1 = 32'd5322
; 
32'd120615: dataIn1 = 32'd5528
; 
32'd120616: dataIn1 = 32'd449
; 
32'd120617: dataIn1 = 32'd5770
; 
32'd120618: dataIn1 = 32'd5771
; 
32'd120619: dataIn1 = 32'd5793
; 
32'd120620: dataIn1 = 32'd5821
; 
32'd120621: dataIn1 = 32'd7001
; 
32'd120622: dataIn1 = 32'd7002
; 
32'd120623: dataIn1 = 32'd450
; 
32'd120624: dataIn1 = 32'd3961
; 
32'd120625: dataIn1 = 32'd3962
; 
32'd120626: dataIn1 = 32'd3993
; 
32'd120627: dataIn1 = 32'd3994
; 
32'd120628: dataIn1 = 32'd5321
; 
32'd120629: dataIn1 = 32'd5324
; 
32'd120630: dataIn1 = 32'd451
; 
32'd120631: dataIn1 = 32'd3966
; 
32'd120632: dataIn1 = 32'd3967
; 
32'd120633: dataIn1 = 32'd3984
; 
32'd120634: dataIn1 = 32'd5273
; 
32'd120635: dataIn1 = 32'd5323
; 
32'd120636: dataIn1 = 32'd5633
; 
32'd120637: dataIn1 = 32'd9320
; 
32'd120638: dataIn1 = 32'd452
; 
32'd120639: dataIn1 = 32'd3980
; 
32'd120640: dataIn1 = 32'd5847
; 
32'd120641: dataIn1 = 32'd5848
; 
32'd120642: dataIn1 = 32'd5870
; 
32'd120643: dataIn1 = 32'd6589
; 
32'd120644: dataIn1 = 32'd6717
; 
32'd120645: dataIn1 = 32'd453
; 
32'd120646: dataIn1 = 32'd3991
; 
32'd120647: dataIn1 = 32'd3992
; 
32'd120648: dataIn1 = 32'd4001
; 
32'd120649: dataIn1 = 32'd4007
; 
32'd120650: dataIn1 = 32'd5325
; 
32'd120651: dataIn1 = 32'd5326
; 
32'd120652: dataIn1 = 32'd454
; 
32'd120653: dataIn1 = 32'd4005
; 
32'd120654: dataIn1 = 32'd4006
; 
32'd120655: dataIn1 = 32'd4013
; 
32'd120656: dataIn1 = 32'd4014
; 
32'd120657: dataIn1 = 32'd5327
; 
32'd120658: dataIn1 = 32'd5329
; 
32'd120659: dataIn1 = 32'd455
; 
32'd120660: dataIn1 = 32'd4017
; 
32'd120661: dataIn1 = 32'd4018
; 
32'd120662: dataIn1 = 32'd4022
; 
32'd120663: dataIn1 = 32'd4031
; 
32'd120664: dataIn1 = 32'd5328
; 
32'd120665: dataIn1 = 32'd5331
; 
32'd120666: dataIn1 = 32'd456
; 
32'd120667: dataIn1 = 32'd4032
; 
32'd120668: dataIn1 = 32'd4033
; 
32'd120669: dataIn1 = 32'd4041
; 
32'd120670: dataIn1 = 32'd4042
; 
32'd120671: dataIn1 = 32'd5330
; 
32'd120672: dataIn1 = 32'd5332
; 
32'd120673: dataIn1 = 32'd457
; 
32'd120674: dataIn1 = 32'd4037
; 
32'd120675: dataIn1 = 32'd4038
; 
32'd120676: dataIn1 = 32'd4049
; 
32'd120677: dataIn1 = 32'd4053
; 
32'd120678: dataIn1 = 32'd5333
; 
32'd120679: dataIn1 = 32'd5335
; 
32'd120680: dataIn1 = 32'd458
; 
32'd120681: dataIn1 = 32'd4054
; 
32'd120682: dataIn1 = 32'd4055
; 
32'd120683: dataIn1 = 32'd4063
; 
32'd120684: dataIn1 = 32'd4064
; 
32'd120685: dataIn1 = 32'd5334
; 
32'd120686: dataIn1 = 32'd5336
; 
32'd120687: dataIn1 = 32'd459
; 
32'd120688: dataIn1 = 32'd4061
; 
32'd120689: dataIn1 = 32'd4062
; 
32'd120690: dataIn1 = 32'd4073
; 
32'd120691: dataIn1 = 32'd4077
; 
32'd120692: dataIn1 = 32'd5337
; 
32'd120693: dataIn1 = 32'd5339
; 
32'd120694: dataIn1 = 32'd460
; 
32'd120695: dataIn1 = 32'd4080
; 
32'd120696: dataIn1 = 32'd4081
; 
32'd120697: dataIn1 = 32'd4089
; 
32'd120698: dataIn1 = 32'd4090
; 
32'd120699: dataIn1 = 32'd5338
; 
32'd120700: dataIn1 = 32'd5340
; 
32'd120701: dataIn1 = 32'd461
; 
32'd120702: dataIn1 = 32'd4087
; 
32'd120703: dataIn1 = 32'd4088
; 
32'd120704: dataIn1 = 32'd4097
; 
32'd120705: dataIn1 = 32'd4103
; 
32'd120706: dataIn1 = 32'd5341
; 
32'd120707: dataIn1 = 32'd5342
; 
32'd120708: dataIn1 = 32'd462
; 
32'd120709: dataIn1 = 32'd4101
; 
32'd120710: dataIn1 = 32'd4102
; 
32'd120711: dataIn1 = 32'd4109
; 
32'd120712: dataIn1 = 32'd4110
; 
32'd120713: dataIn1 = 32'd5343
; 
32'd120714: dataIn1 = 32'd5345
; 
32'd120715: dataIn1 = 32'd463
; 
32'd120716: dataIn1 = 32'd4113
; 
32'd120717: dataIn1 = 32'd4114
; 
32'd120718: dataIn1 = 32'd4118
; 
32'd120719: dataIn1 = 32'd4127
; 
32'd120720: dataIn1 = 32'd5344
; 
32'd120721: dataIn1 = 32'd5347
; 
32'd120722: dataIn1 = 32'd464
; 
32'd120723: dataIn1 = 32'd4128
; 
32'd120724: dataIn1 = 32'd4129
; 
32'd120725: dataIn1 = 32'd4137
; 
32'd120726: dataIn1 = 32'd4138
; 
32'd120727: dataIn1 = 32'd5346
; 
32'd120728: dataIn1 = 32'd5348
; 
32'd120729: dataIn1 = 32'd465
; 
32'd120730: dataIn1 = 32'd4133
; 
32'd120731: dataIn1 = 32'd4134
; 
32'd120732: dataIn1 = 32'd4145
; 
32'd120733: dataIn1 = 32'd4149
; 
32'd120734: dataIn1 = 32'd5349
; 
32'd120735: dataIn1 = 32'd5351
; 
32'd120736: dataIn1 = 32'd466
; 
32'd120737: dataIn1 = 32'd4150
; 
32'd120738: dataIn1 = 32'd4151
; 
32'd120739: dataIn1 = 32'd4159
; 
32'd120740: dataIn1 = 32'd4160
; 
32'd120741: dataIn1 = 32'd5350
; 
32'd120742: dataIn1 = 32'd5352
; 
32'd120743: dataIn1 = 32'd467
; 
32'd120744: dataIn1 = 32'd4157
; 
32'd120745: dataIn1 = 32'd4158
; 
32'd120746: dataIn1 = 32'd4169
; 
32'd120747: dataIn1 = 32'd4173
; 
32'd120748: dataIn1 = 32'd5353
; 
32'd120749: dataIn1 = 32'd5355
; 
32'd120750: dataIn1 = 32'd468
; 
32'd120751: dataIn1 = 32'd4176
; 
32'd120752: dataIn1 = 32'd4177
; 
32'd120753: dataIn1 = 32'd4185
; 
32'd120754: dataIn1 = 32'd4186
; 
32'd120755: dataIn1 = 32'd5354
; 
32'd120756: dataIn1 = 32'd5356
; 
32'd120757: dataIn1 = 32'd469
; 
32'd120758: dataIn1 = 32'd4183
; 
32'd120759: dataIn1 = 32'd4184
; 
32'd120760: dataIn1 = 32'd4193
; 
32'd120761: dataIn1 = 32'd4199
; 
32'd120762: dataIn1 = 32'd5357
; 
32'd120763: dataIn1 = 32'd5358
; 
32'd120764: dataIn1 = 32'd470
; 
32'd120765: dataIn1 = 32'd4197
; 
32'd120766: dataIn1 = 32'd4198
; 
32'd120767: dataIn1 = 32'd4205
; 
32'd120768: dataIn1 = 32'd4206
; 
32'd120769: dataIn1 = 32'd5359
; 
32'd120770: dataIn1 = 32'd5361
; 
32'd120771: dataIn1 = 32'd471
; 
32'd120772: dataIn1 = 32'd4209
; 
32'd120773: dataIn1 = 32'd4210
; 
32'd120774: dataIn1 = 32'd4214
; 
32'd120775: dataIn1 = 32'd4223
; 
32'd120776: dataIn1 = 32'd5360
; 
32'd120777: dataIn1 = 32'd5363
; 
32'd120778: dataIn1 = 32'd472
; 
32'd120779: dataIn1 = 32'd4224
; 
32'd120780: dataIn1 = 32'd4225
; 
32'd120781: dataIn1 = 32'd4233
; 
32'd120782: dataIn1 = 32'd4234
; 
32'd120783: dataIn1 = 32'd5362
; 
32'd120784: dataIn1 = 32'd5364
; 
32'd120785: dataIn1 = 32'd473
; 
32'd120786: dataIn1 = 32'd4229
; 
32'd120787: dataIn1 = 32'd4230
; 
32'd120788: dataIn1 = 32'd4241
; 
32'd120789: dataIn1 = 32'd4245
; 
32'd120790: dataIn1 = 32'd5365
; 
32'd120791: dataIn1 = 32'd5367
; 
32'd120792: dataIn1 = 32'd474
; 
32'd120793: dataIn1 = 32'd4246
; 
32'd120794: dataIn1 = 32'd4247
; 
32'd120795: dataIn1 = 32'd4255
; 
32'd120796: dataIn1 = 32'd4256
; 
32'd120797: dataIn1 = 32'd5366
; 
32'd120798: dataIn1 = 32'd5368
; 
32'd120799: dataIn1 = 32'd475
; 
32'd120800: dataIn1 = 32'd4253
; 
32'd120801: dataIn1 = 32'd4254
; 
32'd120802: dataIn1 = 32'd4265
; 
32'd120803: dataIn1 = 32'd4269
; 
32'd120804: dataIn1 = 32'd5369
; 
32'd120805: dataIn1 = 32'd5371
; 
32'd120806: dataIn1 = 32'd476
; 
32'd120807: dataIn1 = 32'd4272
; 
32'd120808: dataIn1 = 32'd4273
; 
32'd120809: dataIn1 = 32'd4281
; 
32'd120810: dataIn1 = 32'd4282
; 
32'd120811: dataIn1 = 32'd5370
; 
32'd120812: dataIn1 = 32'd5372
; 
32'd120813: dataIn1 = 32'd477
; 
32'd120814: dataIn1 = 32'd4279
; 
32'd120815: dataIn1 = 32'd4280
; 
32'd120816: dataIn1 = 32'd4289
; 
32'd120817: dataIn1 = 32'd4295
; 
32'd120818: dataIn1 = 32'd5373
; 
32'd120819: dataIn1 = 32'd5374
; 
32'd120820: dataIn1 = 32'd478
; 
32'd120821: dataIn1 = 32'd4293
; 
32'd120822: dataIn1 = 32'd4294
; 
32'd120823: dataIn1 = 32'd4301
; 
32'd120824: dataIn1 = 32'd4302
; 
32'd120825: dataIn1 = 32'd5375
; 
32'd120826: dataIn1 = 32'd5377
; 
32'd120827: dataIn1 = 32'd479
; 
32'd120828: dataIn1 = 32'd4305
; 
32'd120829: dataIn1 = 32'd4306
; 
32'd120830: dataIn1 = 32'd4310
; 
32'd120831: dataIn1 = 32'd4319
; 
32'd120832: dataIn1 = 32'd5376
; 
32'd120833: dataIn1 = 32'd5379
; 
32'd120834: dataIn1 = 32'd480
; 
32'd120835: dataIn1 = 32'd4320
; 
32'd120836: dataIn1 = 32'd4321
; 
32'd120837: dataIn1 = 32'd4329
; 
32'd120838: dataIn1 = 32'd4330
; 
32'd120839: dataIn1 = 32'd5378
; 
32'd120840: dataIn1 = 32'd5380
; 
32'd120841: dataIn1 = 32'd481
; 
32'd120842: dataIn1 = 32'd4325
; 
32'd120843: dataIn1 = 32'd4326
; 
32'd120844: dataIn1 = 32'd4337
; 
32'd120845: dataIn1 = 32'd4341
; 
32'd120846: dataIn1 = 32'd5381
; 
32'd120847: dataIn1 = 32'd5383
; 
32'd120848: dataIn1 = 32'd482
; 
32'd120849: dataIn1 = 32'd4342
; 
32'd120850: dataIn1 = 32'd4343
; 
32'd120851: dataIn1 = 32'd4351
; 
32'd120852: dataIn1 = 32'd4352
; 
32'd120853: dataIn1 = 32'd5382
; 
32'd120854: dataIn1 = 32'd5384
; 
32'd120855: dataIn1 = 32'd483
; 
32'd120856: dataIn1 = 32'd4349
; 
32'd120857: dataIn1 = 32'd4350
; 
32'd120858: dataIn1 = 32'd4361
; 
32'd120859: dataIn1 = 32'd4365
; 
32'd120860: dataIn1 = 32'd5385
; 
32'd120861: dataIn1 = 32'd5387
; 
32'd120862: dataIn1 = 32'd484
; 
32'd120863: dataIn1 = 32'd4368
; 
32'd120864: dataIn1 = 32'd4369
; 
32'd120865: dataIn1 = 32'd4377
; 
32'd120866: dataIn1 = 32'd4378
; 
32'd120867: dataIn1 = 32'd5386
; 
32'd120868: dataIn1 = 32'd5388
; 
32'd120869: dataIn1 = 32'd485
; 
32'd120870: dataIn1 = 32'd4375
; 
32'd120871: dataIn1 = 32'd4376
; 
32'd120872: dataIn1 = 32'd4385
; 
32'd120873: dataIn1 = 32'd4391
; 
32'd120874: dataIn1 = 32'd5389
; 
32'd120875: dataIn1 = 32'd5390
; 
32'd120876: dataIn1 = 32'd486
; 
32'd120877: dataIn1 = 32'd4389
; 
32'd120878: dataIn1 = 32'd4390
; 
32'd120879: dataIn1 = 32'd4397
; 
32'd120880: dataIn1 = 32'd4398
; 
32'd120881: dataIn1 = 32'd5391
; 
32'd120882: dataIn1 = 32'd5393
; 
32'd120883: dataIn1 = 32'd487
; 
32'd120884: dataIn1 = 32'd4401
; 
32'd120885: dataIn1 = 32'd4402
; 
32'd120886: dataIn1 = 32'd4406
; 
32'd120887: dataIn1 = 32'd4415
; 
32'd120888: dataIn1 = 32'd5392
; 
32'd120889: dataIn1 = 32'd5395
; 
32'd120890: dataIn1 = 32'd488
; 
32'd120891: dataIn1 = 32'd4416
; 
32'd120892: dataIn1 = 32'd4417
; 
32'd120893: dataIn1 = 32'd4425
; 
32'd120894: dataIn1 = 32'd4426
; 
32'd120895: dataIn1 = 32'd5394
; 
32'd120896: dataIn1 = 32'd5396
; 
32'd120897: dataIn1 = 32'd489
; 
32'd120898: dataIn1 = 32'd4421
; 
32'd120899: dataIn1 = 32'd4422
; 
32'd120900: dataIn1 = 32'd4433
; 
32'd120901: dataIn1 = 32'd4437
; 
32'd120902: dataIn1 = 32'd5397
; 
32'd120903: dataIn1 = 32'd5399
; 
32'd120904: dataIn1 = 32'd490
; 
32'd120905: dataIn1 = 32'd4438
; 
32'd120906: dataIn1 = 32'd4439
; 
32'd120907: dataIn1 = 32'd4447
; 
32'd120908: dataIn1 = 32'd4448
; 
32'd120909: dataIn1 = 32'd5398
; 
32'd120910: dataIn1 = 32'd5400
; 
32'd120911: dataIn1 = 32'd491
; 
32'd120912: dataIn1 = 32'd4445
; 
32'd120913: dataIn1 = 32'd4446
; 
32'd120914: dataIn1 = 32'd4457
; 
32'd120915: dataIn1 = 32'd4461
; 
32'd120916: dataIn1 = 32'd5401
; 
32'd120917: dataIn1 = 32'd5403
; 
32'd120918: dataIn1 = 32'd492
; 
32'd120919: dataIn1 = 32'd4464
; 
32'd120920: dataIn1 = 32'd4465
; 
32'd120921: dataIn1 = 32'd4473
; 
32'd120922: dataIn1 = 32'd4474
; 
32'd120923: dataIn1 = 32'd5402
; 
32'd120924: dataIn1 = 32'd5404
; 
32'd120925: dataIn1 = 32'd493
; 
32'd120926: dataIn1 = 32'd4471
; 
32'd120927: dataIn1 = 32'd4472
; 
32'd120928: dataIn1 = 32'd4481
; 
32'd120929: dataIn1 = 32'd4487
; 
32'd120930: dataIn1 = 32'd5405
; 
32'd120931: dataIn1 = 32'd5406
; 
32'd120932: dataIn1 = 32'd494
; 
32'd120933: dataIn1 = 32'd4485
; 
32'd120934: dataIn1 = 32'd4486
; 
32'd120935: dataIn1 = 32'd4493
; 
32'd120936: dataIn1 = 32'd4494
; 
32'd120937: dataIn1 = 32'd5407
; 
32'd120938: dataIn1 = 32'd5409
; 
32'd120939: dataIn1 = 32'd495
; 
32'd120940: dataIn1 = 32'd4497
; 
32'd120941: dataIn1 = 32'd4498
; 
32'd120942: dataIn1 = 32'd4502
; 
32'd120943: dataIn1 = 32'd4511
; 
32'd120944: dataIn1 = 32'd5408
; 
32'd120945: dataIn1 = 32'd5411
; 
32'd120946: dataIn1 = 32'd496
; 
32'd120947: dataIn1 = 32'd4512
; 
32'd120948: dataIn1 = 32'd4513
; 
32'd120949: dataIn1 = 32'd4521
; 
32'd120950: dataIn1 = 32'd4522
; 
32'd120951: dataIn1 = 32'd5410
; 
32'd120952: dataIn1 = 32'd5412
; 
32'd120953: dataIn1 = 32'd497
; 
32'd120954: dataIn1 = 32'd4517
; 
32'd120955: dataIn1 = 32'd4518
; 
32'd120956: dataIn1 = 32'd4529
; 
32'd120957: dataIn1 = 32'd4533
; 
32'd120958: dataIn1 = 32'd5413
; 
32'd120959: dataIn1 = 32'd5415
; 
32'd120960: dataIn1 = 32'd498
; 
32'd120961: dataIn1 = 32'd4534
; 
32'd120962: dataIn1 = 32'd4535
; 
32'd120963: dataIn1 = 32'd4543
; 
32'd120964: dataIn1 = 32'd4544
; 
32'd120965: dataIn1 = 32'd5414
; 
32'd120966: dataIn1 = 32'd5416
; 
32'd120967: dataIn1 = 32'd499
; 
32'd120968: dataIn1 = 32'd4541
; 
32'd120969: dataIn1 = 32'd4542
; 
32'd120970: dataIn1 = 32'd4553
; 
32'd120971: dataIn1 = 32'd4557
; 
32'd120972: dataIn1 = 32'd5417
; 
32'd120973: dataIn1 = 32'd500
; 
32'd120974: dataIn1 = 32'd4560
; 
32'd120975: dataIn1 = 32'd4561
; 
32'd120976: dataIn1 = 32'd4569
; 
32'd120977: dataIn1 = 32'd4570
; 
32'd120978: dataIn1 = 32'd5418
; 
32'd120979: dataIn1 = 32'd501
; 
32'd120980: dataIn1 = 32'd4567
; 
32'd120981: dataIn1 = 32'd4568
; 
32'd120982: dataIn1 = 32'd4577
; 
32'd120983: dataIn1 = 32'd4583
; 
32'd120984: dataIn1 = 32'd5421
; 
32'd120985: dataIn1 = 32'd502
; 
32'd120986: dataIn1 = 32'd4581
; 
32'd120987: dataIn1 = 32'd4582
; 
32'd120988: dataIn1 = 32'd4589
; 
32'd120989: dataIn1 = 32'd4590
; 
32'd120990: dataIn1 = 32'd5423
; 
32'd120991: dataIn1 = 32'd503
; 
32'd120992: dataIn1 = 32'd4593
; 
32'd120993: dataIn1 = 32'd4594
; 
32'd120994: dataIn1 = 32'd4598
; 
32'd120995: dataIn1 = 32'd5424
; 
32'd120996: dataIn1 = 32'd504
; 
32'd120997: dataIn1 = 32'd1143
; 
32'd120998: dataIn1 = 32'd1144
; 
32'd120999: dataIn1 = 32'd1146
; 
32'd121000: dataIn1 = 32'd1148
; 
32'd121001: dataIn1 = 32'd3558
; 
32'd121002: dataIn1 = 32'd3560
; 
32'd121003: dataIn1 = 32'd505
; 
32'd121004: dataIn1 = 32'd1149
; 
32'd121005: dataIn1 = 32'd1162
; 
32'd121006: dataIn1 = 32'd3560
; 
32'd121007: dataIn1 = 32'd3562
; 
32'd121008: dataIn1 = 32'd11686
; 
32'd121009: dataIn1 = 32'd11687
; 
32'd121010: dataIn1 = 32'd506
; 
32'd121011: dataIn1 = 32'd1149
; 
32'd121012: dataIn1 = 32'd1186
; 
32'd121013: dataIn1 = 32'd3556
; 
32'd121014: dataIn1 = 32'd3558
; 
32'd121015: dataIn1 = 32'd11688
; 
32'd121016: dataIn1 = 32'd11689
; 
32'd121017: dataIn1 = 32'd507
; 
32'd121018: dataIn1 = 32'd1152
; 
32'd121019: dataIn1 = 32'd1153
; 
32'd121020: dataIn1 = 32'd1154
; 
32'd121021: dataIn1 = 32'd1156
; 
32'd121022: dataIn1 = 32'd3574
; 
32'd121023: dataIn1 = 32'd3576
; 
32'd121024: dataIn1 = 32'd508
; 
32'd121025: dataIn1 = 32'd1160
; 
32'd121026: dataIn1 = 32'd1175
; 
32'd121027: dataIn1 = 32'd3576
; 
32'd121028: dataIn1 = 32'd3577
; 
32'd121029: dataIn1 = 32'd11678
; 
32'd121030: dataIn1 = 32'd11679
; 
32'd121031: dataIn1 = 32'd509
; 
32'd121032: dataIn1 = 32'd1160
; 
32'd121033: dataIn1 = 32'd1167
; 
32'd121034: dataIn1 = 32'd3572
; 
32'd121035: dataIn1 = 32'd3574
; 
32'd121036: dataIn1 = 32'd11680
; 
32'd121037: dataIn1 = 32'd11681
; 
32'd121038: dataIn1 = 32'd510
; 
32'd121039: dataIn1 = 32'd1161
; 
32'd121040: dataIn1 = 32'd1162
; 
32'd121041: dataIn1 = 32'd3564
; 
32'd121042: dataIn1 = 32'd3566
; 
32'd121043: dataIn1 = 32'd11684
; 
32'd121044: dataIn1 = 32'd11685
; 
32'd121045: dataIn1 = 32'd511
; 
32'd121046: dataIn1 = 32'd1163
; 
32'd121047: dataIn1 = 32'd1164
; 
32'd121048: dataIn1 = 32'd1165
; 
32'd121049: dataIn1 = 32'd1166
; 
32'd121050: dataIn1 = 32'd3566
; 
32'd121051: dataIn1 = 32'd3568
; 
32'd121052: dataIn1 = 32'd512
; 
32'd121053: dataIn1 = 32'd1161
; 
32'd121054: dataIn1 = 32'd1167
; 
32'd121055: dataIn1 = 32'd3568
; 
32'd121056: dataIn1 = 32'd3570
; 
32'd121057: dataIn1 = 32'd11682
; 
32'd121058: dataIn1 = 32'd11683
; 
32'd121059: dataIn1 = 32'd513
; 
32'd121060: dataIn1 = 32'd1169
; 
32'd121061: dataIn1 = 32'd1170
; 
32'd121062: dataIn1 = 32'd1171
; 
32'd121063: dataIn1 = 32'd1173
; 
32'd121064: dataIn1 = 32'd3579
; 
32'd121065: dataIn1 = 32'd3580
; 
32'd121066: dataIn1 = 32'd514
; 
32'd121067: dataIn1 = 32'd1168
; 
32'd121068: dataIn1 = 32'd1174
; 
32'd121069: dataIn1 = 32'd3580
; 
32'd121070: dataIn1 = 32'd3581
; 
32'd121071: dataIn1 = 32'd11675
; 
32'd121072: dataIn1 = 32'd11676
; 
32'd121073: dataIn1 = 32'd515
; 
32'd121074: dataIn1 = 32'd1168
; 
32'd121075: dataIn1 = 32'd1175
; 
32'd121076: dataIn1 = 32'd3578
; 
32'd121077: dataIn1 = 32'd3579
; 
32'd121078: dataIn1 = 32'd11677
; 
32'd121079: dataIn1 = 32'd516
; 
32'd121080: dataIn1 = 32'd1174
; 
32'd121081: dataIn1 = 32'd3582
; 
32'd121082: dataIn1 = 32'd10683
; 
32'd121083: dataIn1 = 32'd11674
; 
32'd121084: dataIn1 = 32'd517
; 
32'd121085: dataIn1 = 32'd1176
; 
32'd121086: dataIn1 = 32'd1177
; 
32'd121087: dataIn1 = 32'd1179
; 
32'd121088: dataIn1 = 32'd1180
; 
32'd121089: dataIn1 = 32'd3542
; 
32'd121090: dataIn1 = 32'd3544
; 
32'd121091: dataIn1 = 32'd518
; 
32'd121092: dataIn1 = 32'd1183
; 
32'd121093: dataIn1 = 32'd1198
; 
32'd121094: dataIn1 = 32'd3540
; 
32'd121095: dataIn1 = 32'd3542
; 
32'd121096: dataIn1 = 32'd11697
; 
32'd121097: dataIn1 = 32'd11698
; 
32'd121098: dataIn1 = 32'd519
; 
32'd121099: dataIn1 = 32'd1183
; 
32'd121100: dataIn1 = 32'd1187
; 
32'd121101: dataIn1 = 32'd3544
; 
32'd121102: dataIn1 = 32'd3546
; 
32'd121103: dataIn1 = 32'd11694
; 
32'd121104: dataIn1 = 32'd11695
; 
32'd121105: dataIn1 = 32'd11696
; 
32'd121106: dataIn1 = 32'd520
; 
32'd121107: dataIn1 = 32'd1185
; 
32'd121108: dataIn1 = 32'd1186
; 
32'd121109: dataIn1 = 32'd3552
; 
32'd121110: dataIn1 = 32'd3554
; 
32'd121111: dataIn1 = 32'd11690
; 
32'd121112: dataIn1 = 32'd11691
; 
32'd121113: dataIn1 = 32'd521
; 
32'd121114: dataIn1 = 32'd1185
; 
32'd121115: dataIn1 = 32'd1187
; 
32'd121116: dataIn1 = 32'd3548
; 
32'd121117: dataIn1 = 32'd3550
; 
32'd121118: dataIn1 = 32'd11692
; 
32'd121119: dataIn1 = 32'd11693
; 
32'd121120: dataIn1 = 32'd522
; 
32'd121121: dataIn1 = 32'd1188
; 
32'd121122: dataIn1 = 32'd1189
; 
32'd121123: dataIn1 = 32'd1190
; 
32'd121124: dataIn1 = 32'd1191
; 
32'd121125: dataIn1 = 32'd3550
; 
32'd121126: dataIn1 = 32'd3552
; 
32'd121127: dataIn1 = 32'd523
; 
32'd121128: dataIn1 = 32'd1193
; 
32'd121129: dataIn1 = 32'd1194
; 
32'd121130: dataIn1 = 32'd1196
; 
32'd121131: dataIn1 = 32'd1197
; 
32'd121132: dataIn1 = 32'd3534
; 
32'd121133: dataIn1 = 32'd3536
; 
32'd121134: dataIn1 = 32'd524
; 
32'd121135: dataIn1 = 32'd1192
; 
32'd121136: dataIn1 = 32'd1198
; 
32'd121137: dataIn1 = 32'd3536
; 
32'd121138: dataIn1 = 32'd3538
; 
32'd121139: dataIn1 = 32'd11699
; 
32'd121140: dataIn1 = 32'd11700
; 
32'd121141: dataIn1 = 32'd525
; 
32'd121142: dataIn1 = 32'd1192
; 
32'd121143: dataIn1 = 32'd1199
; 
32'd121144: dataIn1 = 32'd3532
; 
32'd121145: dataIn1 = 32'd3534
; 
32'd121146: dataIn1 = 32'd11701
; 
32'd121147: dataIn1 = 32'd11702
; 
32'd121148: dataIn1 = 32'd526
; 
32'd121149: dataIn1 = 32'd1199
; 
32'd121150: dataIn1 = 32'd1206
; 
32'd121151: dataIn1 = 32'd3528
; 
32'd121152: dataIn1 = 32'd3530
; 
32'd121153: dataIn1 = 32'd11703
; 
32'd121154: dataIn1 = 32'd11704
; 
32'd121155: dataIn1 = 32'd527
; 
32'd121156: dataIn1 = 32'd1200
; 
32'd121157: dataIn1 = 32'd1201
; 
32'd121158: dataIn1 = 32'd1203
; 
32'd121159: dataIn1 = 32'd1204
; 
32'd121160: dataIn1 = 32'd3526
; 
32'd121161: dataIn1 = 32'd3528
; 
32'd121162: dataIn1 = 32'd528
; 
32'd121163: dataIn1 = 32'd1206
; 
32'd121164: dataIn1 = 32'd1238
; 
32'd121165: dataIn1 = 32'd3524
; 
32'd121166: dataIn1 = 32'd3526
; 
32'd121167: dataIn1 = 32'd11705
; 
32'd121168: dataIn1 = 32'd11706
; 
32'd121169: dataIn1 = 32'd529
; 
32'd121170: dataIn1 = 32'd1208
; 
32'd121171: dataIn1 = 32'd1209
; 
32'd121172: dataIn1 = 32'd1211
; 
32'd121173: dataIn1 = 32'd1213
; 
32'd121174: dataIn1 = 32'd3486
; 
32'd121175: dataIn1 = 32'd3490
; 
32'd121176: dataIn1 = 32'd530
; 
32'd121177: dataIn1 = 32'd1214
; 
32'd121178: dataIn1 = 32'd1227
; 
32'd121179: dataIn1 = 32'd3490
; 
32'd121180: dataIn1 = 32'd3494
; 
32'd121181: dataIn1 = 32'd11719
; 
32'd121182: dataIn1 = 32'd11720
; 
32'd121183: dataIn1 = 32'd531
; 
32'd121184: dataIn1 = 32'd1214
; 
32'd121185: dataIn1 = 32'd1252
; 
32'd121186: dataIn1 = 32'd3482
; 
32'd121187: dataIn1 = 32'd3486
; 
32'd121188: dataIn1 = 32'd11721
; 
32'd121189: dataIn1 = 32'd11722
; 
32'd121190: dataIn1 = 32'd532
; 
32'd121191: dataIn1 = 32'd1217
; 
32'd121192: dataIn1 = 32'd1218
; 
32'd121193: dataIn1 = 32'd1219
; 
32'd121194: dataIn1 = 32'd1221
; 
32'd121195: dataIn1 = 32'd3510
; 
32'd121196: dataIn1 = 32'd3512
; 
32'd121197: dataIn1 = 32'd533
; 
32'd121198: dataIn1 = 32'd1225
; 
32'd121199: dataIn1 = 32'd1239
; 
32'd121200: dataIn1 = 32'd3512
; 
32'd121201: dataIn1 = 32'd3514
; 
32'd121202: dataIn1 = 32'd11711
; 
32'd121203: dataIn1 = 32'd11712
; 
32'd121204: dataIn1 = 32'd534
; 
32'd121205: dataIn1 = 32'd1225
; 
32'd121206: dataIn1 = 32'd1232
; 
32'd121207: dataIn1 = 32'd3508
; 
32'd121208: dataIn1 = 32'd3510
; 
32'd121209: dataIn1 = 32'd11713
; 
32'd121210: dataIn1 = 32'd11714
; 
32'd121211: dataIn1 = 32'd535
; 
32'd121212: dataIn1 = 32'd1226
; 
32'd121213: dataIn1 = 32'd1227
; 
32'd121214: dataIn1 = 32'd3498
; 
32'd121215: dataIn1 = 32'd3501
; 
32'd121216: dataIn1 = 32'd11717
; 
32'd121217: dataIn1 = 32'd11718
; 
32'd121218: dataIn1 = 32'd536
; 
32'd121219: dataIn1 = 32'd1228
; 
32'd121220: dataIn1 = 32'd1229
; 
32'd121221: dataIn1 = 32'd1230
; 
32'd121222: dataIn1 = 32'd1231
; 
32'd121223: dataIn1 = 32'd3501
; 
32'd121224: dataIn1 = 32'd3504
; 
32'd121225: dataIn1 = 32'd537
; 
32'd121226: dataIn1 = 32'd1226
; 
32'd121227: dataIn1 = 32'd1232
; 
32'd121228: dataIn1 = 32'd3504
; 
32'd121229: dataIn1 = 32'd3506
; 
32'd121230: dataIn1 = 32'd11715
; 
32'd121231: dataIn1 = 32'd11716
; 
32'd121232: dataIn1 = 32'd538
; 
32'd121233: dataIn1 = 32'd1234
; 
32'd121234: dataIn1 = 32'd1235
; 
32'd121235: dataIn1 = 32'd1236
; 
32'd121236: dataIn1 = 32'd1237
; 
32'd121237: dataIn1 = 32'd3518
; 
32'd121238: dataIn1 = 32'd3520
; 
32'd121239: dataIn1 = 32'd539
; 
32'd121240: dataIn1 = 32'd1233
; 
32'd121241: dataIn1 = 32'd1238
; 
32'd121242: dataIn1 = 32'd3520
; 
32'd121243: dataIn1 = 32'd3522
; 
32'd121244: dataIn1 = 32'd11707
; 
32'd121245: dataIn1 = 32'd11708
; 
32'd121246: dataIn1 = 32'd540
; 
32'd121247: dataIn1 = 32'd1233
; 
32'd121248: dataIn1 = 32'd1239
; 
32'd121249: dataIn1 = 32'd3516
; 
32'd121250: dataIn1 = 32'd3518
; 
32'd121251: dataIn1 = 32'd11709
; 
32'd121252: dataIn1 = 32'd11710
; 
32'd121253: dataIn1 = 32'd541
; 
32'd121254: dataIn1 = 32'd1240
; 
32'd121255: dataIn1 = 32'd1241
; 
32'd121256: dataIn1 = 32'd1243
; 
32'd121257: dataIn1 = 32'd1244
; 
32'd121258: dataIn1 = 32'd2753
; 
32'd121259: dataIn1 = 32'd2754
; 
32'd121260: dataIn1 = 32'd542
; 
32'd121261: dataIn1 = 32'd1248
; 
32'd121262: dataIn1 = 32'd1249
; 
32'd121263: dataIn1 = 32'd1262
; 
32'd121264: dataIn1 = 32'd2481
; 
32'd121265: dataIn1 = 32'd2482
; 
32'd121266: dataIn1 = 32'd2753
; 
32'd121267: dataIn1 = 32'd543
; 
32'd121268: dataIn1 = 32'd1247
; 
32'd121269: dataIn1 = 32'd1248
; 
32'd121270: dataIn1 = 32'd1253
; 
32'd121271: dataIn1 = 32'd2754
; 
32'd121272: dataIn1 = 32'd3438
; 
32'd121273: dataIn1 = 32'd11727
; 
32'd121274: dataIn1 = 32'd544
; 
32'd121275: dataIn1 = 32'd1251
; 
32'd121276: dataIn1 = 32'd1252
; 
32'd121277: dataIn1 = 32'd3474
; 
32'd121278: dataIn1 = 32'd3478
; 
32'd121279: dataIn1 = 32'd11723
; 
32'd121280: dataIn1 = 32'd11724
; 
32'd121281: dataIn1 = 32'd545
; 
32'd121282: dataIn1 = 32'd1251
; 
32'd121283: dataIn1 = 32'd1253
; 
32'd121284: dataIn1 = 32'd3458
; 
32'd121285: dataIn1 = 32'd3468
; 
32'd121286: dataIn1 = 32'd11725
; 
32'd121287: dataIn1 = 32'd11726
; 
32'd121288: dataIn1 = 32'd546
; 
32'd121289: dataIn1 = 32'd1254
; 
32'd121290: dataIn1 = 32'd1255
; 
32'd121291: dataIn1 = 32'd1256
; 
32'd121292: dataIn1 = 32'd1257
; 
32'd121293: dataIn1 = 32'd3468
; 
32'd121294: dataIn1 = 32'd3474
; 
32'd121295: dataIn1 = 32'd547
; 
32'd121296: dataIn1 = 32'd1258
; 
32'd121297: dataIn1 = 32'd1259
; 
32'd121298: dataIn1 = 32'd1260
; 
32'd121299: dataIn1 = 32'd2755
; 
32'd121300: dataIn1 = 32'd10250
; 
32'd121301: dataIn1 = 32'd10652
; 
32'd121302: dataIn1 = 32'd266
; 
32'd121303: dataIn1 = 32'd548
; 
32'd121304: dataIn1 = 32'd2480
; 
32'd121305: dataIn1 = 32'd2482
; 
32'd121306: dataIn1 = 32'd2755
; 
32'd121307: dataIn1 = 32'd2756
; 
32'd121308: dataIn1 = 32'd10269
; 
32'd121309: dataIn1 = 32'd266
; 
32'd121310: dataIn1 = 32'd549
; 
32'd121311: dataIn1 = 32'd750
; 
32'd121312: dataIn1 = 32'd1261
; 
32'd121313: dataIn1 = 32'd1262
; 
32'd121314: dataIn1 = 32'd1432
; 
32'd121315: dataIn1 = 32'd2756
; 
32'd121316: dataIn1 = 32'd550
; 
32'd121317: dataIn1 = 32'd959
; 
32'd121318: dataIn1 = 32'd1263
; 
32'd121319: dataIn1 = 32'd1265
; 
32'd121320: dataIn1 = 32'd1266
; 
32'd121321: dataIn1 = 32'd10253
; 
32'd121322: dataIn1 = 32'd10658
; 
32'd121323: dataIn1 = 32'd269
; 
32'd121324: dataIn1 = 32'd551
; 
32'd121325: dataIn1 = 32'd552
; 
32'd121326: dataIn1 = 32'd1268
; 
32'd121327: dataIn1 = 32'd1269
; 
32'd121328: dataIn1 = 32'd11638
; 
32'd121329: dataIn1 = 32'd11639
; 
32'd121330: dataIn1 = 32'd11640
; 
32'd121331: dataIn1 = 32'd268
; 
32'd121332: dataIn1 = 32'd269
; 
32'd121333: dataIn1 = 32'd551
; 
32'd121334: dataIn1 = 32'd552
; 
32'd121335: dataIn1 = 32'd553
; 
32'd121336: dataIn1 = 32'd1268
; 
32'd121337: dataIn1 = 32'd3463
; 
32'd121338: dataIn1 = 32'd3471
; 
32'd121339: dataIn1 = 32'd268
; 
32'd121340: dataIn1 = 32'd552
; 
32'd121341: dataIn1 = 32'd553
; 
32'd121342: dataIn1 = 32'd1268
; 
32'd121343: dataIn1 = 32'd1270
; 
32'd121344: dataIn1 = 32'd11642
; 
32'd121345: dataIn1 = 32'd11643
; 
32'd121346: dataIn1 = 32'd11644
; 
32'd121347: dataIn1 = 32'd269
; 
32'd121348: dataIn1 = 32'd554
; 
32'd121349: dataIn1 = 32'd559
; 
32'd121350: dataIn1 = 32'd1269
; 
32'd121351: dataIn1 = 32'd1274
; 
32'd121352: dataIn1 = 32'd11633
; 
32'd121353: dataIn1 = 32'd11634
; 
32'd121354: dataIn1 = 32'd11635
; 
32'd121355: dataIn1 = 32'd268
; 
32'd121356: dataIn1 = 32'd555
; 
32'd121357: dataIn1 = 32'd1270
; 
32'd121358: dataIn1 = 32'd1273
; 
32'd121359: dataIn1 = 32'd10255
; 
32'd121360: dataIn1 = 32'd11645
; 
32'd121361: dataIn1 = 32'd11646
; 
32'd121362: dataIn1 = 32'd11647
; 
32'd121363: dataIn1 = 32'd270
; 
32'd121364: dataIn1 = 32'd556
; 
32'd121365: dataIn1 = 32'd960
; 
32'd121366: dataIn1 = 32'd1271
; 
32'd121367: dataIn1 = 32'd1272
; 
32'd121368: dataIn1 = 32'd10254
; 
32'd121369: dataIn1 = 32'd11659
; 
32'd121370: dataIn1 = 32'd11660
; 
32'd121371: dataIn1 = 32'd557
; 
32'd121372: dataIn1 = 32'd1273
; 
32'd121373: dataIn1 = 32'd2101
; 
32'd121374: dataIn1 = 32'd10248
; 
32'd121375: dataIn1 = 32'd11650
; 
32'd121376: dataIn1 = 32'd11651
; 
32'd121377: dataIn1 = 32'd11652
; 
32'd121378: dataIn1 = 32'd11654
; 
32'd121379: dataIn1 = 32'd268
; 
32'd121380: dataIn1 = 32'd558
; 
32'd121381: dataIn1 = 32'd960
; 
32'd121382: dataIn1 = 32'd10247
; 
32'd121383: dataIn1 = 32'd10248
; 
32'd121384: dataIn1 = 32'd10254
; 
32'd121385: dataIn1 = 32'd10255
; 
32'd121386: dataIn1 = 32'd269
; 
32'd121387: dataIn1 = 32'd272
; 
32'd121388: dataIn1 = 32'd554
; 
32'd121389: dataIn1 = 32'd559
; 
32'd121390: dataIn1 = 32'd560
; 
32'd121391: dataIn1 = 32'd1274
; 
32'd121392: dataIn1 = 32'd3475
; 
32'd121393: dataIn1 = 32'd3479
; 
32'd121394: dataIn1 = 32'd272
; 
32'd121395: dataIn1 = 32'd559
; 
32'd121396: dataIn1 = 32'd560
; 
32'd121397: dataIn1 = 32'd1274
; 
32'd121398: dataIn1 = 32'd1287
; 
32'd121399: dataIn1 = 32'd11629
; 
32'd121400: dataIn1 = 32'd11630
; 
32'd121401: dataIn1 = 32'd11631
; 
32'd121402: dataIn1 = 32'd274
; 
32'd121403: dataIn1 = 32'd561
; 
32'd121404: dataIn1 = 32'd1275
; 
32'd121405: dataIn1 = 32'd1276
; 
32'd121406: dataIn1 = 32'd1278
; 
32'd121407: dataIn1 = 32'd1720
; 
32'd121408: dataIn1 = 32'd1721
; 
32'd121409: dataIn1 = 32'd274
; 
32'd121410: dataIn1 = 32'd562
; 
32'd121411: dataIn1 = 32'd1276
; 
32'd121412: dataIn1 = 32'd1279
; 
32'd121413: dataIn1 = 32'd11605
; 
32'd121414: dataIn1 = 32'd11606
; 
32'd121415: dataIn1 = 32'd11607
; 
32'd121416: dataIn1 = 32'd274
; 
32'd121417: dataIn1 = 32'd563
; 
32'd121418: dataIn1 = 32'd567
; 
32'd121419: dataIn1 = 32'd1279
; 
32'd121420: dataIn1 = 32'd1285
; 
32'd121421: dataIn1 = 32'd11610
; 
32'd121422: dataIn1 = 32'd11611
; 
32'd121423: dataIn1 = 32'd11612
; 
32'd121424: dataIn1 = 32'd564
; 
32'd121425: dataIn1 = 32'd566
; 
32'd121426: dataIn1 = 32'd1280
; 
32'd121427: dataIn1 = 32'd1283
; 
32'd121428: dataIn1 = 32'd11619
; 
32'd121429: dataIn1 = 32'd11620
; 
32'd121430: dataIn1 = 32'd11621
; 
32'd121431: dataIn1 = 32'd152
; 
32'd121432: dataIn1 = 32'd565
; 
32'd121433: dataIn1 = 32'd566
; 
32'd121434: dataIn1 = 32'd571
; 
32'd121435: dataIn1 = 32'd1283
; 
32'd121436: dataIn1 = 32'd1284
; 
32'd121437: dataIn1 = 32'd1288
; 
32'd121438: dataIn1 = 32'd152
; 
32'd121439: dataIn1 = 32'd275
; 
32'd121440: dataIn1 = 32'd564
; 
32'd121441: dataIn1 = 32'd565
; 
32'd121442: dataIn1 = 32'd566
; 
32'd121443: dataIn1 = 32'd1280
; 
32'd121444: dataIn1 = 32'd1283
; 
32'd121445: dataIn1 = 32'd5457
; 
32'd121446: dataIn1 = 32'd5525
; 
32'd121447: dataIn1 = 32'd274
; 
32'd121448: dataIn1 = 32'd275
; 
32'd121449: dataIn1 = 32'd563
; 
32'd121450: dataIn1 = 32'd567
; 
32'd121451: dataIn1 = 32'd1282
; 
32'd121452: dataIn1 = 32'd1285
; 
32'd121453: dataIn1 = 32'd5525
; 
32'd121454: dataIn1 = 32'd5526
; 
32'd121455: dataIn1 = 32'd272
; 
32'd121456: dataIn1 = 32'd568
; 
32'd121457: dataIn1 = 32'd569
; 
32'd121458: dataIn1 = 32'd1286
; 
32'd121459: dataIn1 = 32'd1287
; 
32'd121460: dataIn1 = 32'd11625
; 
32'd121461: dataIn1 = 32'd11626
; 
32'd121462: dataIn1 = 32'd11627
; 
32'd121463: dataIn1 = 32'd272
; 
32'd121464: dataIn1 = 32'd277
; 
32'd121465: dataIn1 = 32'd568
; 
32'd121466: dataIn1 = 32'd569
; 
32'd121467: dataIn1 = 32'd570
; 
32'd121468: dataIn1 = 32'd1286
; 
32'd121469: dataIn1 = 32'd3483
; 
32'd121470: dataIn1 = 32'd3487
; 
32'd121471: dataIn1 = 32'd277
; 
32'd121472: dataIn1 = 32'd569
; 
32'd121473: dataIn1 = 32'd570
; 
32'd121474: dataIn1 = 32'd571
; 
32'd121475: dataIn1 = 32'd1286
; 
32'd121476: dataIn1 = 32'd1288
; 
32'd121477: dataIn1 = 32'd11624
; 
32'd121478: dataIn1 = 32'd152
; 
32'd121479: dataIn1 = 32'd277
; 
32'd121480: dataIn1 = 32'd565
; 
32'd121481: dataIn1 = 32'd570
; 
32'd121482: dataIn1 = 32'd571
; 
32'd121483: dataIn1 = 32'd1288
; 
32'd121484: dataIn1 = 32'd3495
; 
32'd121485: dataIn1 = 32'd3499
; 
32'd121486: dataIn1 = 32'd278
; 
32'd121487: dataIn1 = 32'd572
; 
32'd121488: dataIn1 = 32'd1289
; 
32'd121489: dataIn1 = 32'd1290
; 
32'd121490: dataIn1 = 32'd1292
; 
32'd121491: dataIn1 = 32'd1721
; 
32'd121492: dataIn1 = 32'd1722
; 
32'd121493: dataIn1 = 32'd278
; 
32'd121494: dataIn1 = 32'd573
; 
32'd121495: dataIn1 = 32'd1290
; 
32'd121496: dataIn1 = 32'd1293
; 
32'd121497: dataIn1 = 32'd11594
; 
32'd121498: dataIn1 = 32'd11595
; 
32'd121499: dataIn1 = 32'd11596
; 
32'd121500: dataIn1 = 32'd278
; 
32'd121501: dataIn1 = 32'd574
; 
32'd121502: dataIn1 = 32'd582
; 
32'd121503: dataIn1 = 32'd1293
; 
32'd121504: dataIn1 = 32'd1298
; 
32'd121505: dataIn1 = 32'd11589
; 
32'd121506: dataIn1 = 32'd11590
; 
32'd121507: dataIn1 = 32'd11591
; 
32'd121508: dataIn1 = 32'd280
; 
32'd121509: dataIn1 = 32'd281
; 
32'd121510: dataIn1 = 32'd575
; 
32'd121511: dataIn1 = 32'd576
; 
32'd121512: dataIn1 = 32'd577
; 
32'd121513: dataIn1 = 32'd1294
; 
32'd121514: dataIn1 = 32'd5532
; 
32'd121515: dataIn1 = 32'd5533
; 
32'd121516: dataIn1 = 32'd281
; 
32'd121517: dataIn1 = 32'd575
; 
32'd121518: dataIn1 = 32'd576
; 
32'd121519: dataIn1 = 32'd1294
; 
32'd121520: dataIn1 = 32'd1295
; 
32'd121521: dataIn1 = 32'd11581
; 
32'd121522: dataIn1 = 32'd11582
; 
32'd121523: dataIn1 = 32'd11583
; 
32'd121524: dataIn1 = 32'd280
; 
32'd121525: dataIn1 = 32'd575
; 
32'd121526: dataIn1 = 32'd577
; 
32'd121527: dataIn1 = 32'd1294
; 
32'd121528: dataIn1 = 32'd1296
; 
32'd121529: dataIn1 = 32'd11577
; 
32'd121530: dataIn1 = 32'd11578
; 
32'd121531: dataIn1 = 32'd11579
; 
32'd121532: dataIn1 = 32'd281
; 
32'd121533: dataIn1 = 32'd578
; 
32'd121534: dataIn1 = 32'd582
; 
32'd121535: dataIn1 = 32'd1295
; 
32'd121536: dataIn1 = 32'd1298
; 
32'd121537: dataIn1 = 32'd11585
; 
32'd121538: dataIn1 = 32'd11586
; 
32'd121539: dataIn1 = 32'd11587
; 
32'd121540: dataIn1 = 32'd280
; 
32'd121541: dataIn1 = 32'd579
; 
32'd121542: dataIn1 = 32'd581
; 
32'd121543: dataIn1 = 32'd1296
; 
32'd121544: dataIn1 = 32'd1297
; 
32'd121545: dataIn1 = 32'd11573
; 
32'd121546: dataIn1 = 32'd11574
; 
32'd121547: dataIn1 = 32'd11575
; 
32'd121548: dataIn1 = 32'd282
; 
32'd121549: dataIn1 = 32'd580
; 
32'd121550: dataIn1 = 32'd581
; 
32'd121551: dataIn1 = 32'd1297
; 
32'd121552: dataIn1 = 32'd1308
; 
32'd121553: dataIn1 = 32'd11569
; 
32'd121554: dataIn1 = 32'd11570
; 
32'd121555: dataIn1 = 32'd11571
; 
32'd121556: dataIn1 = 32'd280
; 
32'd121557: dataIn1 = 32'd282
; 
32'd121558: dataIn1 = 32'd579
; 
32'd121559: dataIn1 = 32'd580
; 
32'd121560: dataIn1 = 32'd581
; 
32'd121561: dataIn1 = 32'd1297
; 
32'd121562: dataIn1 = 32'd5534
; 
32'd121563: dataIn1 = 32'd5535
; 
32'd121564: dataIn1 = 32'd278
; 
32'd121565: dataIn1 = 32'd281
; 
32'd121566: dataIn1 = 32'd574
; 
32'd121567: dataIn1 = 32'd578
; 
32'd121568: dataIn1 = 32'd582
; 
32'd121569: dataIn1 = 32'd1298
; 
32'd121570: dataIn1 = 32'd5530
; 
32'd121571: dataIn1 = 32'd5531
; 
32'd121572: dataIn1 = 32'd583
; 
32'd121573: dataIn1 = 32'd1299
; 
32'd121574: dataIn1 = 32'd2757
; 
32'd121575: dataIn1 = 32'd2766
; 
32'd121576: dataIn1 = 32'd2768
; 
32'd121577: dataIn1 = 32'd10985
; 
32'd121578: dataIn1 = 32'd10986
; 
32'd121579: dataIn1 = 32'd10987
; 
32'd121580: dataIn1 = 32'd584
; 
32'd121581: dataIn1 = 32'd1300
; 
32'd121582: dataIn1 = 32'd2483
; 
32'd121583: dataIn1 = 32'd2484
; 
32'd121584: dataIn1 = 32'd10981
; 
32'd121585: dataIn1 = 32'd10982
; 
32'd121586: dataIn1 = 32'd10983
; 
32'd121587: dataIn1 = 32'd585
; 
32'd121588: dataIn1 = 32'd1300
; 
32'd121589: dataIn1 = 32'd1518
; 
32'd121590: dataIn1 = 32'd2487
; 
32'd121591: dataIn1 = 32'd2488
; 
32'd121592: dataIn1 = 32'd2522
; 
32'd121593: dataIn1 = 32'd10978
; 
32'd121594: dataIn1 = 32'd10979
; 
32'd121595: dataIn1 = 32'd586
; 
32'd121596: dataIn1 = 32'd2483
; 
32'd121597: dataIn1 = 32'd2485
; 
32'd121598: dataIn1 = 32'd2486
; 
32'd121599: dataIn1 = 32'd2488
; 
32'd121600: dataIn1 = 32'd3420
; 
32'd121601: dataIn1 = 32'd3421
; 
32'd121602: dataIn1 = 32'd288
; 
32'd121603: dataIn1 = 32'd587
; 
32'd121604: dataIn1 = 32'd588
; 
32'd121605: dataIn1 = 32'd1301
; 
32'd121606: dataIn1 = 32'd1302
; 
32'd121607: dataIn1 = 32'd11549
; 
32'd121608: dataIn1 = 32'd11550
; 
32'd121609: dataIn1 = 32'd11551
; 
32'd121610: dataIn1 = 32'd287
; 
32'd121611: dataIn1 = 32'd288
; 
32'd121612: dataIn1 = 32'd587
; 
32'd121613: dataIn1 = 32'd588
; 
32'd121614: dataIn1 = 32'd589
; 
32'd121615: dataIn1 = 32'd1301
; 
32'd121616: dataIn1 = 32'd5540
; 
32'd121617: dataIn1 = 32'd5541
; 
32'd121618: dataIn1 = 32'd287
; 
32'd121619: dataIn1 = 32'd588
; 
32'd121620: dataIn1 = 32'd589
; 
32'd121621: dataIn1 = 32'd1301
; 
32'd121622: dataIn1 = 32'd1303
; 
32'd121623: dataIn1 = 32'd11546
; 
32'd121624: dataIn1 = 32'd11547
; 
32'd121625: dataIn1 = 32'd11548
; 
32'd121626: dataIn1 = 32'd288
; 
32'd121627: dataIn1 = 32'd590
; 
32'd121628: dataIn1 = 32'd594
; 
32'd121629: dataIn1 = 32'd1302
; 
32'd121630: dataIn1 = 32'd1305
; 
32'd121631: dataIn1 = 32'd11553
; 
32'd121632: dataIn1 = 32'd11554
; 
32'd121633: dataIn1 = 32'd11555
; 
32'd121634: dataIn1 = 32'd11556
; 
32'd121635: dataIn1 = 32'd287
; 
32'd121636: dataIn1 = 32'd591
; 
32'd121637: dataIn1 = 32'd593
; 
32'd121638: dataIn1 = 32'd1303
; 
32'd121639: dataIn1 = 32'd1304
; 
32'd121640: dataIn1 = 32'd11542
; 
32'd121641: dataIn1 = 32'd11543
; 
32'd121642: dataIn1 = 32'd11544
; 
32'd121643: dataIn1 = 32'd289
; 
32'd121644: dataIn1 = 32'd592
; 
32'd121645: dataIn1 = 32'd593
; 
32'd121646: dataIn1 = 32'd1304
; 
32'd121647: dataIn1 = 32'd1311
; 
32'd121648: dataIn1 = 32'd11537
; 
32'd121649: dataIn1 = 32'd11538
; 
32'd121650: dataIn1 = 32'd11539
; 
32'd121651: dataIn1 = 32'd287
; 
32'd121652: dataIn1 = 32'd289
; 
32'd121653: dataIn1 = 32'd591
; 
32'd121654: dataIn1 = 32'd592
; 
32'd121655: dataIn1 = 32'd593
; 
32'd121656: dataIn1 = 32'd1304
; 
32'd121657: dataIn1 = 32'd5542
; 
32'd121658: dataIn1 = 32'd5543
; 
32'd121659: dataIn1 = 32'd288
; 
32'd121660: dataIn1 = 32'd292
; 
32'd121661: dataIn1 = 32'd590
; 
32'd121662: dataIn1 = 32'd594
; 
32'd121663: dataIn1 = 32'd595
; 
32'd121664: dataIn1 = 32'd1305
; 
32'd121665: dataIn1 = 32'd5538
; 
32'd121666: dataIn1 = 32'd5539
; 
32'd121667: dataIn1 = 32'd292
; 
32'd121668: dataIn1 = 32'd594
; 
32'd121669: dataIn1 = 32'd595
; 
32'd121670: dataIn1 = 32'd1305
; 
32'd121671: dataIn1 = 32'd1307
; 
32'd121672: dataIn1 = 32'd11558
; 
32'd121673: dataIn1 = 32'd11559
; 
32'd121674: dataIn1 = 32'd11560
; 
32'd121675: dataIn1 = 32'd292
; 
32'd121676: dataIn1 = 32'd596
; 
32'd121677: dataIn1 = 32'd598
; 
32'd121678: dataIn1 = 32'd1306
; 
32'd121679: dataIn1 = 32'd1307
; 
32'd121680: dataIn1 = 32'd11562
; 
32'd121681: dataIn1 = 32'd11563
; 
32'd121682: dataIn1 = 32'd11564
; 
32'd121683: dataIn1 = 32'd282
; 
32'd121684: dataIn1 = 32'd597
; 
32'd121685: dataIn1 = 32'd598
; 
32'd121686: dataIn1 = 32'd1306
; 
32'd121687: dataIn1 = 32'd1308
; 
32'd121688: dataIn1 = 32'd11566
; 
32'd121689: dataIn1 = 32'd11567
; 
32'd121690: dataIn1 = 32'd282
; 
32'd121691: dataIn1 = 32'd292
; 
32'd121692: dataIn1 = 32'd596
; 
32'd121693: dataIn1 = 32'd597
; 
32'd121694: dataIn1 = 32'd598
; 
32'd121695: dataIn1 = 32'd1306
; 
32'd121696: dataIn1 = 32'd5536
; 
32'd121697: dataIn1 = 32'd5537
; 
32'd121698: dataIn1 = 32'd289
; 
32'd121699: dataIn1 = 32'd294
; 
32'd121700: dataIn1 = 32'd599
; 
32'd121701: dataIn1 = 32'd600
; 
32'd121702: dataIn1 = 32'd601
; 
32'd121703: dataIn1 = 32'd1309
; 
32'd121704: dataIn1 = 32'd5544
; 
32'd121705: dataIn1 = 32'd5545
; 
32'd121706: dataIn1 = 32'd294
; 
32'd121707: dataIn1 = 32'd599
; 
32'd121708: dataIn1 = 32'd600
; 
32'd121709: dataIn1 = 32'd1309
; 
32'd121710: dataIn1 = 32'd1310
; 
32'd121711: dataIn1 = 32'd11530
; 
32'd121712: dataIn1 = 32'd11531
; 
32'd121713: dataIn1 = 32'd11532
; 
32'd121714: dataIn1 = 32'd289
; 
32'd121715: dataIn1 = 32'd599
; 
32'd121716: dataIn1 = 32'd601
; 
32'd121717: dataIn1 = 32'd1309
; 
32'd121718: dataIn1 = 32'd1311
; 
32'd121719: dataIn1 = 32'd11534
; 
32'd121720: dataIn1 = 32'd11535
; 
32'd121721: dataIn1 = 32'd11536
; 
32'd121722: dataIn1 = 32'd294
; 
32'd121723: dataIn1 = 32'd602
; 
32'd121724: dataIn1 = 32'd610
; 
32'd121725: dataIn1 = 32'd1310
; 
32'd121726: dataIn1 = 32'd1316
; 
32'd121727: dataIn1 = 32'd11526
; 
32'd121728: dataIn1 = 32'd11527
; 
32'd121729: dataIn1 = 32'd11528
; 
32'd121730: dataIn1 = 32'd296
; 
32'd121731: dataIn1 = 32'd297
; 
32'd121732: dataIn1 = 32'd603
; 
32'd121733: dataIn1 = 32'd604
; 
32'd121734: dataIn1 = 32'd605
; 
32'd121735: dataIn1 = 32'd1312
; 
32'd121736: dataIn1 = 32'd5548
; 
32'd121737: dataIn1 = 32'd5549
; 
32'd121738: dataIn1 = 32'd297
; 
32'd121739: dataIn1 = 32'd603
; 
32'd121740: dataIn1 = 32'd604
; 
32'd121741: dataIn1 = 32'd1312
; 
32'd121742: dataIn1 = 32'd1313
; 
32'd121743: dataIn1 = 32'd11517
; 
32'd121744: dataIn1 = 32'd11518
; 
32'd121745: dataIn1 = 32'd11519
; 
32'd121746: dataIn1 = 32'd296
; 
32'd121747: dataIn1 = 32'd603
; 
32'd121748: dataIn1 = 32'd605
; 
32'd121749: dataIn1 = 32'd1312
; 
32'd121750: dataIn1 = 32'd1314
; 
32'd121751: dataIn1 = 32'd11513
; 
32'd121752: dataIn1 = 32'd11514
; 
32'd121753: dataIn1 = 32'd11515
; 
32'd121754: dataIn1 = 32'd297
; 
32'd121755: dataIn1 = 32'd606
; 
32'd121756: dataIn1 = 32'd610
; 
32'd121757: dataIn1 = 32'd1313
; 
32'd121758: dataIn1 = 32'd1316
; 
32'd121759: dataIn1 = 32'd11521
; 
32'd121760: dataIn1 = 32'd11522
; 
32'd121761: dataIn1 = 32'd11523
; 
32'd121762: dataIn1 = 32'd11524
; 
32'd121763: dataIn1 = 32'd296
; 
32'd121764: dataIn1 = 32'd607
; 
32'd121765: dataIn1 = 32'd609
; 
32'd121766: dataIn1 = 32'd1314
; 
32'd121767: dataIn1 = 32'd1315
; 
32'd121768: dataIn1 = 32'd11509
; 
32'd121769: dataIn1 = 32'd11510
; 
32'd121770: dataIn1 = 32'd11511
; 
32'd121771: dataIn1 = 32'd298
; 
32'd121772: dataIn1 = 32'd608
; 
32'd121773: dataIn1 = 32'd609
; 
32'd121774: dataIn1 = 32'd1315
; 
32'd121775: dataIn1 = 32'd1324
; 
32'd121776: dataIn1 = 32'd11505
; 
32'd121777: dataIn1 = 32'd11506
; 
32'd121778: dataIn1 = 32'd11507
; 
32'd121779: dataIn1 = 32'd296
; 
32'd121780: dataIn1 = 32'd298
; 
32'd121781: dataIn1 = 32'd607
; 
32'd121782: dataIn1 = 32'd608
; 
32'd121783: dataIn1 = 32'd609
; 
32'd121784: dataIn1 = 32'd1315
; 
32'd121785: dataIn1 = 32'd5550
; 
32'd121786: dataIn1 = 32'd5551
; 
32'd121787: dataIn1 = 32'd294
; 
32'd121788: dataIn1 = 32'd297
; 
32'd121789: dataIn1 = 32'd602
; 
32'd121790: dataIn1 = 32'd606
; 
32'd121791: dataIn1 = 32'd610
; 
32'd121792: dataIn1 = 32'd1316
; 
32'd121793: dataIn1 = 32'd5546
; 
32'd121794: dataIn1 = 32'd5547
; 
32'd121795: dataIn1 = 32'd304
; 
32'd121796: dataIn1 = 32'd611
; 
32'd121797: dataIn1 = 32'd612
; 
32'd121798: dataIn1 = 32'd1317
; 
32'd121799: dataIn1 = 32'd1318
; 
32'd121800: dataIn1 = 32'd11486
; 
32'd121801: dataIn1 = 32'd11487
; 
32'd121802: dataIn1 = 32'd11488
; 
32'd121803: dataIn1 = 32'd303
; 
32'd121804: dataIn1 = 32'd304
; 
32'd121805: dataIn1 = 32'd611
; 
32'd121806: dataIn1 = 32'd612
; 
32'd121807: dataIn1 = 32'd613
; 
32'd121808: dataIn1 = 32'd1317
; 
32'd121809: dataIn1 = 32'd5556
; 
32'd121810: dataIn1 = 32'd5557
; 
32'd121811: dataIn1 = 32'd303
; 
32'd121812: dataIn1 = 32'd612
; 
32'd121813: dataIn1 = 32'd613
; 
32'd121814: dataIn1 = 32'd1317
; 
32'd121815: dataIn1 = 32'd1319
; 
32'd121816: dataIn1 = 32'd11482
; 
32'd121817: dataIn1 = 32'd11483
; 
32'd121818: dataIn1 = 32'd11484
; 
32'd121819: dataIn1 = 32'd304
; 
32'd121820: dataIn1 = 32'd614
; 
32'd121821: dataIn1 = 32'd618
; 
32'd121822: dataIn1 = 32'd1318
; 
32'd121823: dataIn1 = 32'd1321
; 
32'd121824: dataIn1 = 32'd11490
; 
32'd121825: dataIn1 = 32'd11491
; 
32'd121826: dataIn1 = 32'd11492
; 
32'd121827: dataIn1 = 32'd303
; 
32'd121828: dataIn1 = 32'd615
; 
32'd121829: dataIn1 = 32'd617
; 
32'd121830: dataIn1 = 32'd1319
; 
32'd121831: dataIn1 = 32'd1320
; 
32'd121832: dataIn1 = 32'd11478
; 
32'd121833: dataIn1 = 32'd11479
; 
32'd121834: dataIn1 = 32'd11480
; 
32'd121835: dataIn1 = 32'd305
; 
32'd121836: dataIn1 = 32'd616
; 
32'd121837: dataIn1 = 32'd617
; 
32'd121838: dataIn1 = 32'd1320
; 
32'd121839: dataIn1 = 32'd1327
; 
32'd121840: dataIn1 = 32'd11474
; 
32'd121841: dataIn1 = 32'd11475
; 
32'd121842: dataIn1 = 32'd11476
; 
32'd121843: dataIn1 = 32'd303
; 
32'd121844: dataIn1 = 32'd305
; 
32'd121845: dataIn1 = 32'd615
; 
32'd121846: dataIn1 = 32'd616
; 
32'd121847: dataIn1 = 32'd617
; 
32'd121848: dataIn1 = 32'd1320
; 
32'd121849: dataIn1 = 32'd5558
; 
32'd121850: dataIn1 = 32'd5559
; 
32'd121851: dataIn1 = 32'd304
; 
32'd121852: dataIn1 = 32'd308
; 
32'd121853: dataIn1 = 32'd614
; 
32'd121854: dataIn1 = 32'd618
; 
32'd121855: dataIn1 = 32'd619
; 
32'd121856: dataIn1 = 32'd1321
; 
32'd121857: dataIn1 = 32'd5554
; 
32'd121858: dataIn1 = 32'd5555
; 
32'd121859: dataIn1 = 32'd308
; 
32'd121860: dataIn1 = 32'd618
; 
32'd121861: dataIn1 = 32'd619
; 
32'd121862: dataIn1 = 32'd1321
; 
32'd121863: dataIn1 = 32'd1323
; 
32'd121864: dataIn1 = 32'd11494
; 
32'd121865: dataIn1 = 32'd11495
; 
32'd121866: dataIn1 = 32'd11496
; 
32'd121867: dataIn1 = 32'd308
; 
32'd121868: dataIn1 = 32'd620
; 
32'd121869: dataIn1 = 32'd622
; 
32'd121870: dataIn1 = 32'd1322
; 
32'd121871: dataIn1 = 32'd1323
; 
32'd121872: dataIn1 = 32'd11498
; 
32'd121873: dataIn1 = 32'd11499
; 
32'd121874: dataIn1 = 32'd298
; 
32'd121875: dataIn1 = 32'd621
; 
32'd121876: dataIn1 = 32'd622
; 
32'd121877: dataIn1 = 32'd1322
; 
32'd121878: dataIn1 = 32'd1324
; 
32'd121879: dataIn1 = 32'd11501
; 
32'd121880: dataIn1 = 32'd11502
; 
32'd121881: dataIn1 = 32'd11503
; 
32'd121882: dataIn1 = 32'd298
; 
32'd121883: dataIn1 = 32'd308
; 
32'd121884: dataIn1 = 32'd620
; 
32'd121885: dataIn1 = 32'd621
; 
32'd121886: dataIn1 = 32'd622
; 
32'd121887: dataIn1 = 32'd1322
; 
32'd121888: dataIn1 = 32'd5552
; 
32'd121889: dataIn1 = 32'd5553
; 
32'd121890: dataIn1 = 32'd305
; 
32'd121891: dataIn1 = 32'd310
; 
32'd121892: dataIn1 = 32'd623
; 
32'd121893: dataIn1 = 32'd624
; 
32'd121894: dataIn1 = 32'd625
; 
32'd121895: dataIn1 = 32'd1325
; 
32'd121896: dataIn1 = 32'd5560
; 
32'd121897: dataIn1 = 32'd5561
; 
32'd121898: dataIn1 = 32'd310
; 
32'd121899: dataIn1 = 32'd623
; 
32'd121900: dataIn1 = 32'd624
; 
32'd121901: dataIn1 = 32'd1325
; 
32'd121902: dataIn1 = 32'd1326
; 
32'd121903: dataIn1 = 32'd11466
; 
32'd121904: dataIn1 = 32'd11467
; 
32'd121905: dataIn1 = 32'd11468
; 
32'd121906: dataIn1 = 32'd305
; 
32'd121907: dataIn1 = 32'd623
; 
32'd121908: dataIn1 = 32'd625
; 
32'd121909: dataIn1 = 32'd1325
; 
32'd121910: dataIn1 = 32'd1327
; 
32'd121911: dataIn1 = 32'd11470
; 
32'd121912: dataIn1 = 32'd11471
; 
32'd121913: dataIn1 = 32'd11472
; 
32'd121914: dataIn1 = 32'd310
; 
32'd121915: dataIn1 = 32'd626
; 
32'd121916: dataIn1 = 32'd634
; 
32'd121917: dataIn1 = 32'd1326
; 
32'd121918: dataIn1 = 32'd1332
; 
32'd121919: dataIn1 = 32'd11461
; 
32'd121920: dataIn1 = 32'd11462
; 
32'd121921: dataIn1 = 32'd11463
; 
32'd121922: dataIn1 = 32'd312
; 
32'd121923: dataIn1 = 32'd313
; 
32'd121924: dataIn1 = 32'd627
; 
32'd121925: dataIn1 = 32'd628
; 
32'd121926: dataIn1 = 32'd629
; 
32'd121927: dataIn1 = 32'd1328
; 
32'd121928: dataIn1 = 32'd5564
; 
32'd121929: dataIn1 = 32'd5565
; 
32'd121930: dataIn1 = 32'd313
; 
32'd121931: dataIn1 = 32'd627
; 
32'd121932: dataIn1 = 32'd628
; 
32'd121933: dataIn1 = 32'd1328
; 
32'd121934: dataIn1 = 32'd1329
; 
32'd121935: dataIn1 = 32'd11453
; 
32'd121936: dataIn1 = 32'd11454
; 
32'd121937: dataIn1 = 32'd11455
; 
32'd121938: dataIn1 = 32'd312
; 
32'd121939: dataIn1 = 32'd627
; 
32'd121940: dataIn1 = 32'd629
; 
32'd121941: dataIn1 = 32'd1328
; 
32'd121942: dataIn1 = 32'd1330
; 
32'd121943: dataIn1 = 32'd11449
; 
32'd121944: dataIn1 = 32'd11450
; 
32'd121945: dataIn1 = 32'd11451
; 
32'd121946: dataIn1 = 32'd313
; 
32'd121947: dataIn1 = 32'd630
; 
32'd121948: dataIn1 = 32'd634
; 
32'd121949: dataIn1 = 32'd1329
; 
32'd121950: dataIn1 = 32'd1332
; 
32'd121951: dataIn1 = 32'd11457
; 
32'd121952: dataIn1 = 32'd11458
; 
32'd121953: dataIn1 = 32'd11459
; 
32'd121954: dataIn1 = 32'd312
; 
32'd121955: dataIn1 = 32'd631
; 
32'd121956: dataIn1 = 32'd633
; 
32'd121957: dataIn1 = 32'd1330
; 
32'd121958: dataIn1 = 32'd1331
; 
32'd121959: dataIn1 = 32'd11445
; 
32'd121960: dataIn1 = 32'd11446
; 
32'd121961: dataIn1 = 32'd11447
; 
32'd121962: dataIn1 = 32'd314
; 
32'd121963: dataIn1 = 32'd632
; 
32'd121964: dataIn1 = 32'd633
; 
32'd121965: dataIn1 = 32'd1331
; 
32'd121966: dataIn1 = 32'd1340
; 
32'd121967: dataIn1 = 32'd11441
; 
32'd121968: dataIn1 = 32'd11442
; 
32'd121969: dataIn1 = 32'd11443
; 
32'd121970: dataIn1 = 32'd312
; 
32'd121971: dataIn1 = 32'd314
; 
32'd121972: dataIn1 = 32'd631
; 
32'd121973: dataIn1 = 32'd632
; 
32'd121974: dataIn1 = 32'd633
; 
32'd121975: dataIn1 = 32'd1331
; 
32'd121976: dataIn1 = 32'd5566
; 
32'd121977: dataIn1 = 32'd5567
; 
32'd121978: dataIn1 = 32'd310
; 
32'd121979: dataIn1 = 32'd313
; 
32'd121980: dataIn1 = 32'd626
; 
32'd121981: dataIn1 = 32'd630
; 
32'd121982: dataIn1 = 32'd634
; 
32'd121983: dataIn1 = 32'd1332
; 
32'd121984: dataIn1 = 32'd5562
; 
32'd121985: dataIn1 = 32'd5563
; 
32'd121986: dataIn1 = 32'd320
; 
32'd121987: dataIn1 = 32'd635
; 
32'd121988: dataIn1 = 32'd636
; 
32'd121989: dataIn1 = 32'd1333
; 
32'd121990: dataIn1 = 32'd1334
; 
32'd121991: dataIn1 = 32'd11421
; 
32'd121992: dataIn1 = 32'd11422
; 
32'd121993: dataIn1 = 32'd11423
; 
32'd121994: dataIn1 = 32'd319
; 
32'd121995: dataIn1 = 32'd320
; 
32'd121996: dataIn1 = 32'd635
; 
32'd121997: dataIn1 = 32'd636
; 
32'd121998: dataIn1 = 32'd637
; 
32'd121999: dataIn1 = 32'd1333
; 
32'd122000: dataIn1 = 32'd5572
; 
32'd122001: dataIn1 = 32'd5573
; 
32'd122002: dataIn1 = 32'd319
; 
32'd122003: dataIn1 = 32'd636
; 
32'd122004: dataIn1 = 32'd637
; 
32'd122005: dataIn1 = 32'd1333
; 
32'd122006: dataIn1 = 32'd1335
; 
32'd122007: dataIn1 = 32'd11417
; 
32'd122008: dataIn1 = 32'd11418
; 
32'd122009: dataIn1 = 32'd11419
; 
32'd122010: dataIn1 = 32'd320
; 
32'd122011: dataIn1 = 32'd638
; 
32'd122012: dataIn1 = 32'd642
; 
32'd122013: dataIn1 = 32'd1334
; 
32'd122014: dataIn1 = 32'd1337
; 
32'd122015: dataIn1 = 32'd11426
; 
32'd122016: dataIn1 = 32'd11427
; 
32'd122017: dataIn1 = 32'd11428
; 
32'd122018: dataIn1 = 32'd319
; 
32'd122019: dataIn1 = 32'd639
; 
32'd122020: dataIn1 = 32'd641
; 
32'd122021: dataIn1 = 32'd1335
; 
32'd122022: dataIn1 = 32'd1336
; 
32'd122023: dataIn1 = 32'd11414
; 
32'd122024: dataIn1 = 32'd11415
; 
32'd122025: dataIn1 = 32'd321
; 
32'd122026: dataIn1 = 32'd640
; 
32'd122027: dataIn1 = 32'd641
; 
32'd122028: dataIn1 = 32'd1336
; 
32'd122029: dataIn1 = 32'd1343
; 
32'd122030: dataIn1 = 32'd11409
; 
32'd122031: dataIn1 = 32'd11410
; 
32'd122032: dataIn1 = 32'd11411
; 
32'd122033: dataIn1 = 32'd319
; 
32'd122034: dataIn1 = 32'd321
; 
32'd122035: dataIn1 = 32'd639
; 
32'd122036: dataIn1 = 32'd640
; 
32'd122037: dataIn1 = 32'd641
; 
32'd122038: dataIn1 = 32'd1336
; 
32'd122039: dataIn1 = 32'd5574
; 
32'd122040: dataIn1 = 32'd5575
; 
32'd122041: dataIn1 = 32'd320
; 
32'd122042: dataIn1 = 32'd324
; 
32'd122043: dataIn1 = 32'd638
; 
32'd122044: dataIn1 = 32'd642
; 
32'd122045: dataIn1 = 32'd643
; 
32'd122046: dataIn1 = 32'd1337
; 
32'd122047: dataIn1 = 32'd5570
; 
32'd122048: dataIn1 = 32'd5571
; 
32'd122049: dataIn1 = 32'd324
; 
32'd122050: dataIn1 = 32'd642
; 
32'd122051: dataIn1 = 32'd643
; 
32'd122052: dataIn1 = 32'd1337
; 
32'd122053: dataIn1 = 32'd1339
; 
32'd122054: dataIn1 = 32'd11430
; 
32'd122055: dataIn1 = 32'd11431
; 
32'd122056: dataIn1 = 32'd324
; 
32'd122057: dataIn1 = 32'd644
; 
32'd122058: dataIn1 = 32'd646
; 
32'd122059: dataIn1 = 32'd1338
; 
32'd122060: dataIn1 = 32'd1339
; 
32'd122061: dataIn1 = 32'd11434
; 
32'd122062: dataIn1 = 32'd11435
; 
32'd122063: dataIn1 = 32'd11436
; 
32'd122064: dataIn1 = 32'd314
; 
32'd122065: dataIn1 = 32'd645
; 
32'd122066: dataIn1 = 32'd646
; 
32'd122067: dataIn1 = 32'd1338
; 
32'd122068: dataIn1 = 32'd1340
; 
32'd122069: dataIn1 = 32'd11438
; 
32'd122070: dataIn1 = 32'd11439
; 
32'd122071: dataIn1 = 32'd314
; 
32'd122072: dataIn1 = 32'd324
; 
32'd122073: dataIn1 = 32'd644
; 
32'd122074: dataIn1 = 32'd645
; 
32'd122075: dataIn1 = 32'd646
; 
32'd122076: dataIn1 = 32'd1338
; 
32'd122077: dataIn1 = 32'd5568
; 
32'd122078: dataIn1 = 32'd5569
; 
32'd122079: dataIn1 = 32'd321
; 
32'd122080: dataIn1 = 32'd326
; 
32'd122081: dataIn1 = 32'd647
; 
32'd122082: dataIn1 = 32'd648
; 
32'd122083: dataIn1 = 32'd649
; 
32'd122084: dataIn1 = 32'd1341
; 
32'd122085: dataIn1 = 32'd5576
; 
32'd122086: dataIn1 = 32'd5577
; 
32'd122087: dataIn1 = 32'd326
; 
32'd122088: dataIn1 = 32'd647
; 
32'd122089: dataIn1 = 32'd648
; 
32'd122090: dataIn1 = 32'd1341
; 
32'd122091: dataIn1 = 32'd1342
; 
32'd122092: dataIn1 = 32'd11402
; 
32'd122093: dataIn1 = 32'd11403
; 
32'd122094: dataIn1 = 32'd321
; 
32'd122095: dataIn1 = 32'd647
; 
32'd122096: dataIn1 = 32'd649
; 
32'd122097: dataIn1 = 32'd1341
; 
32'd122098: dataIn1 = 32'd1343
; 
32'd122099: dataIn1 = 32'd11405
; 
32'd122100: dataIn1 = 32'd11406
; 
32'd122101: dataIn1 = 32'd11407
; 
32'd122102: dataIn1 = 32'd326
; 
32'd122103: dataIn1 = 32'd650
; 
32'd122104: dataIn1 = 32'd658
; 
32'd122105: dataIn1 = 32'd1342
; 
32'd122106: dataIn1 = 32'd1348
; 
32'd122107: dataIn1 = 32'd11397
; 
32'd122108: dataIn1 = 32'd11398
; 
32'd122109: dataIn1 = 32'd11399
; 
32'd122110: dataIn1 = 32'd11400
; 
32'd122111: dataIn1 = 32'd328
; 
32'd122112: dataIn1 = 32'd329
; 
32'd122113: dataIn1 = 32'd651
; 
32'd122114: dataIn1 = 32'd652
; 
32'd122115: dataIn1 = 32'd653
; 
32'd122116: dataIn1 = 32'd1344
; 
32'd122117: dataIn1 = 32'd5580
; 
32'd122118: dataIn1 = 32'd5581
; 
32'd122119: dataIn1 = 32'd329
; 
32'd122120: dataIn1 = 32'd651
; 
32'd122121: dataIn1 = 32'd652
; 
32'd122122: dataIn1 = 32'd1344
; 
32'd122123: dataIn1 = 32'd1345
; 
32'd122124: dataIn1 = 32'd11389
; 
32'd122125: dataIn1 = 32'd11390
; 
32'd122126: dataIn1 = 32'd11391
; 
32'd122127: dataIn1 = 32'd328
; 
32'd122128: dataIn1 = 32'd651
; 
32'd122129: dataIn1 = 32'd653
; 
32'd122130: dataIn1 = 32'd1344
; 
32'd122131: dataIn1 = 32'd1346
; 
32'd122132: dataIn1 = 32'd11385
; 
32'd122133: dataIn1 = 32'd11386
; 
32'd122134: dataIn1 = 32'd11387
; 
32'd122135: dataIn1 = 32'd329
; 
32'd122136: dataIn1 = 32'd654
; 
32'd122137: dataIn1 = 32'd658
; 
32'd122138: dataIn1 = 32'd1345
; 
32'd122139: dataIn1 = 32'd1348
; 
32'd122140: dataIn1 = 32'd11394
; 
32'd122141: dataIn1 = 32'd11395
; 
32'd122142: dataIn1 = 32'd328
; 
32'd122143: dataIn1 = 32'd655
; 
32'd122144: dataIn1 = 32'd657
; 
32'd122145: dataIn1 = 32'd1346
; 
32'd122146: dataIn1 = 32'd1347
; 
32'd122147: dataIn1 = 32'd11381
; 
32'd122148: dataIn1 = 32'd11382
; 
32'd122149: dataIn1 = 32'd11383
; 
32'd122150: dataIn1 = 32'd11384
; 
32'd122151: dataIn1 = 32'd330
; 
32'd122152: dataIn1 = 32'd656
; 
32'd122153: dataIn1 = 32'd657
; 
32'd122154: dataIn1 = 32'd1347
; 
32'd122155: dataIn1 = 32'd1356
; 
32'd122156: dataIn1 = 32'd11378
; 
32'd122157: dataIn1 = 32'd11379
; 
32'd122158: dataIn1 = 32'd11380
; 
32'd122159: dataIn1 = 32'd328
; 
32'd122160: dataIn1 = 32'd330
; 
32'd122161: dataIn1 = 32'd655
; 
32'd122162: dataIn1 = 32'd656
; 
32'd122163: dataIn1 = 32'd657
; 
32'd122164: dataIn1 = 32'd1347
; 
32'd122165: dataIn1 = 32'd5582
; 
32'd122166: dataIn1 = 32'd5583
; 
32'd122167: dataIn1 = 32'd326
; 
32'd122168: dataIn1 = 32'd329
; 
32'd122169: dataIn1 = 32'd650
; 
32'd122170: dataIn1 = 32'd654
; 
32'd122171: dataIn1 = 32'd658
; 
32'd122172: dataIn1 = 32'd1348
; 
32'd122173: dataIn1 = 32'd5578
; 
32'd122174: dataIn1 = 32'd5579
; 
32'd122175: dataIn1 = 32'd336
; 
32'd122176: dataIn1 = 32'd659
; 
32'd122177: dataIn1 = 32'd660
; 
32'd122178: dataIn1 = 32'd1349
; 
32'd122179: dataIn1 = 32'd1350
; 
32'd122180: dataIn1 = 32'd11357
; 
32'd122181: dataIn1 = 32'd11358
; 
32'd122182: dataIn1 = 32'd11359
; 
32'd122183: dataIn1 = 32'd11360
; 
32'd122184: dataIn1 = 32'd335
; 
32'd122185: dataIn1 = 32'd336
; 
32'd122186: dataIn1 = 32'd659
; 
32'd122187: dataIn1 = 32'd660
; 
32'd122188: dataIn1 = 32'd661
; 
32'd122189: dataIn1 = 32'd1349
; 
32'd122190: dataIn1 = 32'd5588
; 
32'd122191: dataIn1 = 32'd5589
; 
32'd122192: dataIn1 = 32'd335
; 
32'd122193: dataIn1 = 32'd660
; 
32'd122194: dataIn1 = 32'd661
; 
32'd122195: dataIn1 = 32'd1349
; 
32'd122196: dataIn1 = 32'd1351
; 
32'd122197: dataIn1 = 32'd11354
; 
32'd122198: dataIn1 = 32'd11355
; 
32'd122199: dataIn1 = 32'd336
; 
32'd122200: dataIn1 = 32'd662
; 
32'd122201: dataIn1 = 32'd666
; 
32'd122202: dataIn1 = 32'd1350
; 
32'd122203: dataIn1 = 32'd1353
; 
32'd122204: dataIn1 = 32'd11362
; 
32'd122205: dataIn1 = 32'd11363
; 
32'd122206: dataIn1 = 32'd11364
; 
32'd122207: dataIn1 = 32'd335
; 
32'd122208: dataIn1 = 32'd663
; 
32'd122209: dataIn1 = 32'd665
; 
32'd122210: dataIn1 = 32'd1351
; 
32'd122211: dataIn1 = 32'd1352
; 
32'd122212: dataIn1 = 32'd11350
; 
32'd122213: dataIn1 = 32'd11351
; 
32'd122214: dataIn1 = 32'd337
; 
32'd122215: dataIn1 = 32'd664
; 
32'd122216: dataIn1 = 32'd665
; 
32'd122217: dataIn1 = 32'd1352
; 
32'd122218: dataIn1 = 32'd1359
; 
32'd122219: dataIn1 = 32'd11346
; 
32'd122220: dataIn1 = 32'd11347
; 
32'd122221: dataIn1 = 32'd335
; 
32'd122222: dataIn1 = 32'd337
; 
32'd122223: dataIn1 = 32'd663
; 
32'd122224: dataIn1 = 32'd664
; 
32'd122225: dataIn1 = 32'd665
; 
32'd122226: dataIn1 = 32'd1352
; 
32'd122227: dataIn1 = 32'd5590
; 
32'd122228: dataIn1 = 32'd5591
; 
32'd122229: dataIn1 = 32'd336
; 
32'd122230: dataIn1 = 32'd340
; 
32'd122231: dataIn1 = 32'd662
; 
32'd122232: dataIn1 = 32'd666
; 
32'd122233: dataIn1 = 32'd667
; 
32'd122234: dataIn1 = 32'd1353
; 
32'd122235: dataIn1 = 32'd5586
; 
32'd122236: dataIn1 = 32'd5587
; 
32'd122237: dataIn1 = 32'd340
; 
32'd122238: dataIn1 = 32'd666
; 
32'd122239: dataIn1 = 32'd667
; 
32'd122240: dataIn1 = 32'd1353
; 
32'd122241: dataIn1 = 32'd1355
; 
32'd122242: dataIn1 = 32'd11365
; 
32'd122243: dataIn1 = 32'd11366
; 
32'd122244: dataIn1 = 32'd11367
; 
32'd122245: dataIn1 = 32'd340
; 
32'd122246: dataIn1 = 32'd668
; 
32'd122247: dataIn1 = 32'd670
; 
32'd122248: dataIn1 = 32'd1354
; 
32'd122249: dataIn1 = 32'd1355
; 
32'd122250: dataIn1 = 32'd11370
; 
32'd122251: dataIn1 = 32'd11371
; 
32'd122252: dataIn1 = 32'd330
; 
32'd122253: dataIn1 = 32'd669
; 
32'd122254: dataIn1 = 32'd670
; 
32'd122255: dataIn1 = 32'd1354
; 
32'd122256: dataIn1 = 32'd1356
; 
32'd122257: dataIn1 = 32'd11374
; 
32'd122258: dataIn1 = 32'd11375
; 
32'd122259: dataIn1 = 32'd330
; 
32'd122260: dataIn1 = 32'd340
; 
32'd122261: dataIn1 = 32'd668
; 
32'd122262: dataIn1 = 32'd669
; 
32'd122263: dataIn1 = 32'd670
; 
32'd122264: dataIn1 = 32'd1354
; 
32'd122265: dataIn1 = 32'd5584
; 
32'd122266: dataIn1 = 32'd5585
; 
32'd122267: dataIn1 = 32'd337
; 
32'd122268: dataIn1 = 32'd342
; 
32'd122269: dataIn1 = 32'd671
; 
32'd122270: dataIn1 = 32'd672
; 
32'd122271: dataIn1 = 32'd673
; 
32'd122272: dataIn1 = 32'd1357
; 
32'd122273: dataIn1 = 32'd5592
; 
32'd122274: dataIn1 = 32'd5593
; 
32'd122275: dataIn1 = 32'd342
; 
32'd122276: dataIn1 = 32'd671
; 
32'd122277: dataIn1 = 32'd672
; 
32'd122278: dataIn1 = 32'd1357
; 
32'd122279: dataIn1 = 32'd1358
; 
32'd122280: dataIn1 = 32'd11337
; 
32'd122281: dataIn1 = 32'd11338
; 
32'd122282: dataIn1 = 32'd11339
; 
32'd122283: dataIn1 = 32'd11340
; 
32'd122284: dataIn1 = 32'd337
; 
32'd122285: dataIn1 = 32'd671
; 
32'd122286: dataIn1 = 32'd673
; 
32'd122287: dataIn1 = 32'd1357
; 
32'd122288: dataIn1 = 32'd1359
; 
32'd122289: dataIn1 = 32'd11342
; 
32'd122290: dataIn1 = 32'd11343
; 
32'd122291: dataIn1 = 32'd11344
; 
32'd122292: dataIn1 = 32'd342
; 
32'd122293: dataIn1 = 32'd674
; 
32'd122294: dataIn1 = 32'd682
; 
32'd122295: dataIn1 = 32'd1358
; 
32'd122296: dataIn1 = 32'd1364
; 
32'd122297: dataIn1 = 32'd11334
; 
32'd122298: dataIn1 = 32'd11335
; 
32'd122299: dataIn1 = 32'd344
; 
32'd122300: dataIn1 = 32'd345
; 
32'd122301: dataIn1 = 32'd675
; 
32'd122302: dataIn1 = 32'd676
; 
32'd122303: dataIn1 = 32'd677
; 
32'd122304: dataIn1 = 32'd1360
; 
32'd122305: dataIn1 = 32'd5596
; 
32'd122306: dataIn1 = 32'd5597
; 
32'd122307: dataIn1 = 32'd345
; 
32'd122308: dataIn1 = 32'd675
; 
32'd122309: dataIn1 = 32'd676
; 
32'd122310: dataIn1 = 32'd1360
; 
32'd122311: dataIn1 = 32'd1361
; 
32'd122312: dataIn1 = 32'd11326
; 
32'd122313: dataIn1 = 32'd11327
; 
32'd122314: dataIn1 = 32'd344
; 
32'd122315: dataIn1 = 32'd675
; 
32'd122316: dataIn1 = 32'd677
; 
32'd122317: dataIn1 = 32'd1360
; 
32'd122318: dataIn1 = 32'd1362
; 
32'd122319: dataIn1 = 32'd11322
; 
32'd122320: dataIn1 = 32'd11323
; 
32'd122321: dataIn1 = 32'd345
; 
32'd122322: dataIn1 = 32'd678
; 
32'd122323: dataIn1 = 32'd682
; 
32'd122324: dataIn1 = 32'd1361
; 
32'd122325: dataIn1 = 32'd1364
; 
32'd122326: dataIn1 = 32'd11330
; 
32'd122327: dataIn1 = 32'd11331
; 
32'd122328: dataIn1 = 32'd11332
; 
32'd122329: dataIn1 = 32'd344
; 
32'd122330: dataIn1 = 32'd679
; 
32'd122331: dataIn1 = 32'd681
; 
32'd122332: dataIn1 = 32'd1362
; 
32'd122333: dataIn1 = 32'd1363
; 
32'd122334: dataIn1 = 32'd11317
; 
32'd122335: dataIn1 = 32'd11318
; 
32'd122336: dataIn1 = 32'd11319
; 
32'd122337: dataIn1 = 32'd346
; 
32'd122338: dataIn1 = 32'd680
; 
32'd122339: dataIn1 = 32'd681
; 
32'd122340: dataIn1 = 32'd1363
; 
32'd122341: dataIn1 = 32'd1372
; 
32'd122342: dataIn1 = 32'd11313
; 
32'd122343: dataIn1 = 32'd11314
; 
32'd122344: dataIn1 = 32'd11315
; 
32'd122345: dataIn1 = 32'd344
; 
32'd122346: dataIn1 = 32'd346
; 
32'd122347: dataIn1 = 32'd679
; 
32'd122348: dataIn1 = 32'd680
; 
32'd122349: dataIn1 = 32'd681
; 
32'd122350: dataIn1 = 32'd1363
; 
32'd122351: dataIn1 = 32'd5598
; 
32'd122352: dataIn1 = 32'd5599
; 
32'd122353: dataIn1 = 32'd342
; 
32'd122354: dataIn1 = 32'd345
; 
32'd122355: dataIn1 = 32'd674
; 
32'd122356: dataIn1 = 32'd678
; 
32'd122357: dataIn1 = 32'd682
; 
32'd122358: dataIn1 = 32'd1364
; 
32'd122359: dataIn1 = 32'd5594
; 
32'd122360: dataIn1 = 32'd5595
; 
32'd122361: dataIn1 = 32'd352
; 
32'd122362: dataIn1 = 32'd683
; 
32'd122363: dataIn1 = 32'd684
; 
32'd122364: dataIn1 = 32'd1365
; 
32'd122365: dataIn1 = 32'd1366
; 
32'd122366: dataIn1 = 32'd11293
; 
32'd122367: dataIn1 = 32'd11294
; 
32'd122368: dataIn1 = 32'd11295
; 
32'd122369: dataIn1 = 32'd351
; 
32'd122370: dataIn1 = 32'd352
; 
32'd122371: dataIn1 = 32'd683
; 
32'd122372: dataIn1 = 32'd684
; 
32'd122373: dataIn1 = 32'd685
; 
32'd122374: dataIn1 = 32'd1365
; 
32'd122375: dataIn1 = 32'd5604
; 
32'd122376: dataIn1 = 32'd5605
; 
32'd122377: dataIn1 = 32'd351
; 
32'd122378: dataIn1 = 32'd684
; 
32'd122379: dataIn1 = 32'd685
; 
32'd122380: dataIn1 = 32'd1365
; 
32'd122381: dataIn1 = 32'd1367
; 
32'd122382: dataIn1 = 32'd11290
; 
32'd122383: dataIn1 = 32'd11291
; 
32'd122384: dataIn1 = 32'd352
; 
32'd122385: dataIn1 = 32'd686
; 
32'd122386: dataIn1 = 32'd690
; 
32'd122387: dataIn1 = 32'd1366
; 
32'd122388: dataIn1 = 32'd1369
; 
32'd122389: dataIn1 = 32'd11298
; 
32'd122390: dataIn1 = 32'd11299
; 
32'd122391: dataIn1 = 32'd351
; 
32'd122392: dataIn1 = 32'd687
; 
32'd122393: dataIn1 = 32'd689
; 
32'd122394: dataIn1 = 32'd1367
; 
32'd122395: dataIn1 = 32'd1368
; 
32'd122396: dataIn1 = 32'd11285
; 
32'd122397: dataIn1 = 32'd11286
; 
32'd122398: dataIn1 = 32'd11287
; 
32'd122399: dataIn1 = 32'd11288
; 
32'd122400: dataIn1 = 32'd353
; 
32'd122401: dataIn1 = 32'd688
; 
32'd122402: dataIn1 = 32'd689
; 
32'd122403: dataIn1 = 32'd1368
; 
32'd122404: dataIn1 = 32'd1375
; 
32'd122405: dataIn1 = 32'd11282
; 
32'd122406: dataIn1 = 32'd11283
; 
32'd122407: dataIn1 = 32'd351
; 
32'd122408: dataIn1 = 32'd353
; 
32'd122409: dataIn1 = 32'd687
; 
32'd122410: dataIn1 = 32'd688
; 
32'd122411: dataIn1 = 32'd689
; 
32'd122412: dataIn1 = 32'd1368
; 
32'd122413: dataIn1 = 32'd5606
; 
32'd122414: dataIn1 = 32'd5607
; 
32'd122415: dataIn1 = 32'd352
; 
32'd122416: dataIn1 = 32'd356
; 
32'd122417: dataIn1 = 32'd686
; 
32'd122418: dataIn1 = 32'd690
; 
32'd122419: dataIn1 = 32'd691
; 
32'd122420: dataIn1 = 32'd1369
; 
32'd122421: dataIn1 = 32'd5602
; 
32'd122422: dataIn1 = 32'd5603
; 
32'd122423: dataIn1 = 32'd356
; 
32'd122424: dataIn1 = 32'd690
; 
32'd122425: dataIn1 = 32'd691
; 
32'd122426: dataIn1 = 32'd1369
; 
32'd122427: dataIn1 = 32'd1371
; 
32'd122428: dataIn1 = 32'd11302
; 
32'd122429: dataIn1 = 32'd11303
; 
32'd122430: dataIn1 = 32'd356
; 
32'd122431: dataIn1 = 32'd692
; 
32'd122432: dataIn1 = 32'd694
; 
32'd122433: dataIn1 = 32'd1370
; 
32'd122434: dataIn1 = 32'd1371
; 
32'd122435: dataIn1 = 32'd11306
; 
32'd122436: dataIn1 = 32'd11307
; 
32'd122437: dataIn1 = 32'd346
; 
32'd122438: dataIn1 = 32'd693
; 
32'd122439: dataIn1 = 32'd694
; 
32'd122440: dataIn1 = 32'd1370
; 
32'd122441: dataIn1 = 32'd1372
; 
32'd122442: dataIn1 = 32'd11309
; 
32'd122443: dataIn1 = 32'd11310
; 
32'd122444: dataIn1 = 32'd11311
; 
32'd122445: dataIn1 = 32'd346
; 
32'd122446: dataIn1 = 32'd356
; 
32'd122447: dataIn1 = 32'd692
; 
32'd122448: dataIn1 = 32'd693
; 
32'd122449: dataIn1 = 32'd694
; 
32'd122450: dataIn1 = 32'd1370
; 
32'd122451: dataIn1 = 32'd5600
; 
32'd122452: dataIn1 = 32'd5601
; 
32'd122453: dataIn1 = 32'd353
; 
32'd122454: dataIn1 = 32'd358
; 
32'd122455: dataIn1 = 32'd695
; 
32'd122456: dataIn1 = 32'd696
; 
32'd122457: dataIn1 = 32'd697
; 
32'd122458: dataIn1 = 32'd1373
; 
32'd122459: dataIn1 = 32'd5608
; 
32'd122460: dataIn1 = 32'd5609
; 
32'd122461: dataIn1 = 32'd358
; 
32'd122462: dataIn1 = 32'd695
; 
32'd122463: dataIn1 = 32'd696
; 
32'd122464: dataIn1 = 32'd1373
; 
32'd122465: dataIn1 = 32'd1374
; 
32'd122466: dataIn1 = 32'd11274
; 
32'd122467: dataIn1 = 32'd11275
; 
32'd122468: dataIn1 = 32'd353
; 
32'd122469: dataIn1 = 32'd695
; 
32'd122470: dataIn1 = 32'd697
; 
32'd122471: dataIn1 = 32'd1373
; 
32'd122472: dataIn1 = 32'd1375
; 
32'd122473: dataIn1 = 32'd11278
; 
32'd122474: dataIn1 = 32'd11279
; 
32'd122475: dataIn1 = 32'd358
; 
32'd122476: dataIn1 = 32'd698
; 
32'd122477: dataIn1 = 32'd706
; 
32'd122478: dataIn1 = 32'd1374
; 
32'd122479: dataIn1 = 32'd1380
; 
32'd122480: dataIn1 = 32'd11270
; 
32'd122481: dataIn1 = 32'd11271
; 
32'd122482: dataIn1 = 32'd360
; 
32'd122483: dataIn1 = 32'd361
; 
32'd122484: dataIn1 = 32'd699
; 
32'd122485: dataIn1 = 32'd700
; 
32'd122486: dataIn1 = 32'd701
; 
32'd122487: dataIn1 = 32'd1376
; 
32'd122488: dataIn1 = 32'd5612
; 
32'd122489: dataIn1 = 32'd5613
; 
32'd122490: dataIn1 = 32'd361
; 
32'd122491: dataIn1 = 32'd699
; 
32'd122492: dataIn1 = 32'd700
; 
32'd122493: dataIn1 = 32'd1376
; 
32'd122494: dataIn1 = 32'd1377
; 
32'd122495: dataIn1 = 32'd11262
; 
32'd122496: dataIn1 = 32'd11263
; 
32'd122497: dataIn1 = 32'd11264
; 
32'd122498: dataIn1 = 32'd360
; 
32'd122499: dataIn1 = 32'd699
; 
32'd122500: dataIn1 = 32'd701
; 
32'd122501: dataIn1 = 32'd1376
; 
32'd122502: dataIn1 = 32'd1378
; 
32'd122503: dataIn1 = 32'd11258
; 
32'd122504: dataIn1 = 32'd11259
; 
32'd122505: dataIn1 = 32'd361
; 
32'd122506: dataIn1 = 32'd702
; 
32'd122507: dataIn1 = 32'd706
; 
32'd122508: dataIn1 = 32'd1377
; 
32'd122509: dataIn1 = 32'd1380
; 
32'd122510: dataIn1 = 32'd11265
; 
32'd122511: dataIn1 = 32'd11266
; 
32'd122512: dataIn1 = 32'd11267
; 
32'd122513: dataIn1 = 32'd11268
; 
32'd122514: dataIn1 = 32'd360
; 
32'd122515: dataIn1 = 32'd703
; 
32'd122516: dataIn1 = 32'd705
; 
32'd122517: dataIn1 = 32'd1378
; 
32'd122518: dataIn1 = 32'd1379
; 
32'd122519: dataIn1 = 32'd11254
; 
32'd122520: dataIn1 = 32'd11255
; 
32'd122521: dataIn1 = 32'd11256
; 
32'd122522: dataIn1 = 32'd362
; 
32'd122523: dataIn1 = 32'd704
; 
32'd122524: dataIn1 = 32'd705
; 
32'd122525: dataIn1 = 32'd1379
; 
32'd122526: dataIn1 = 32'd1388
; 
32'd122527: dataIn1 = 32'd11250
; 
32'd122528: dataIn1 = 32'd11251
; 
32'd122529: dataIn1 = 32'd360
; 
32'd122530: dataIn1 = 32'd362
; 
32'd122531: dataIn1 = 32'd703
; 
32'd122532: dataIn1 = 32'd704
; 
32'd122533: dataIn1 = 32'd705
; 
32'd122534: dataIn1 = 32'd1379
; 
32'd122535: dataIn1 = 32'd5614
; 
32'd122536: dataIn1 = 32'd5615
; 
32'd122537: dataIn1 = 32'd358
; 
32'd122538: dataIn1 = 32'd361
; 
32'd122539: dataIn1 = 32'd698
; 
32'd122540: dataIn1 = 32'd702
; 
32'd122541: dataIn1 = 32'd706
; 
32'd122542: dataIn1 = 32'd1380
; 
32'd122543: dataIn1 = 32'd5610
; 
32'd122544: dataIn1 = 32'd5611
; 
32'd122545: dataIn1 = 32'd368
; 
32'd122546: dataIn1 = 32'd707
; 
32'd122547: dataIn1 = 32'd708
; 
32'd122548: dataIn1 = 32'd1381
; 
32'd122549: dataIn1 = 32'd1382
; 
32'd122550: dataIn1 = 32'd11229
; 
32'd122551: dataIn1 = 32'd11230
; 
32'd122552: dataIn1 = 32'd11231
; 
32'd122553: dataIn1 = 32'd367
; 
32'd122554: dataIn1 = 32'd368
; 
32'd122555: dataIn1 = 32'd707
; 
32'd122556: dataIn1 = 32'd708
; 
32'd122557: dataIn1 = 32'd709
; 
32'd122558: dataIn1 = 32'd1381
; 
32'd122559: dataIn1 = 32'd5620
; 
32'd122560: dataIn1 = 32'd5621
; 
32'd122561: dataIn1 = 32'd367
; 
32'd122562: dataIn1 = 32'd708
; 
32'd122563: dataIn1 = 32'd709
; 
32'd122564: dataIn1 = 32'd1381
; 
32'd122565: dataIn1 = 32'd1383
; 
32'd122566: dataIn1 = 32'd11225
; 
32'd122567: dataIn1 = 32'd11226
; 
32'd122568: dataIn1 = 32'd11227
; 
32'd122569: dataIn1 = 32'd368
; 
32'd122570: dataIn1 = 32'd710
; 
32'd122571: dataIn1 = 32'd714
; 
32'd122572: dataIn1 = 32'd1382
; 
32'd122573: dataIn1 = 32'd1385
; 
32'd122574: dataIn1 = 32'd11234
; 
32'd122575: dataIn1 = 32'd11235
; 
32'd122576: dataIn1 = 32'd11236
; 
32'd122577: dataIn1 = 32'd367
; 
32'd122578: dataIn1 = 32'd711
; 
32'd122579: dataIn1 = 32'd713
; 
32'd122580: dataIn1 = 32'd1383
; 
32'd122581: dataIn1 = 32'd1384
; 
32'd122582: dataIn1 = 32'd11222
; 
32'd122583: dataIn1 = 32'd11223
; 
32'd122584: dataIn1 = 32'd369
; 
32'd122585: dataIn1 = 32'd712
; 
32'd122586: dataIn1 = 32'd713
; 
32'd122587: dataIn1 = 32'd1384
; 
32'd122588: dataIn1 = 32'd1391
; 
32'd122589: dataIn1 = 32'd11217
; 
32'd122590: dataIn1 = 32'd11218
; 
32'd122591: dataIn1 = 32'd11219
; 
32'd122592: dataIn1 = 32'd11220
; 
32'd122593: dataIn1 = 32'd367
; 
32'd122594: dataIn1 = 32'd369
; 
32'd122595: dataIn1 = 32'd711
; 
32'd122596: dataIn1 = 32'd712
; 
32'd122597: dataIn1 = 32'd713
; 
32'd122598: dataIn1 = 32'd1384
; 
32'd122599: dataIn1 = 32'd5622
; 
32'd122600: dataIn1 = 32'd5623
; 
32'd122601: dataIn1 = 32'd368
; 
32'd122602: dataIn1 = 32'd372
; 
32'd122603: dataIn1 = 32'd710
; 
32'd122604: dataIn1 = 32'd714
; 
32'd122605: dataIn1 = 32'd715
; 
32'd122606: dataIn1 = 32'd1385
; 
32'd122607: dataIn1 = 32'd5618
; 
32'd122608: dataIn1 = 32'd5619
; 
32'd122609: dataIn1 = 32'd372
; 
32'd122610: dataIn1 = 32'd714
; 
32'd122611: dataIn1 = 32'd715
; 
32'd122612: dataIn1 = 32'd1385
; 
32'd122613: dataIn1 = 32'd1387
; 
32'd122614: dataIn1 = 32'd11237
; 
32'd122615: dataIn1 = 32'd11238
; 
32'd122616: dataIn1 = 32'd11239
; 
32'd122617: dataIn1 = 32'd372
; 
32'd122618: dataIn1 = 32'd716
; 
32'd122619: dataIn1 = 32'd718
; 
32'd122620: dataIn1 = 32'd1386
; 
32'd122621: dataIn1 = 32'd1387
; 
32'd122622: dataIn1 = 32'd11241
; 
32'd122623: dataIn1 = 32'd11242
; 
32'd122624: dataIn1 = 32'd11243
; 
32'd122625: dataIn1 = 32'd362
; 
32'd122626: dataIn1 = 32'd717
; 
32'd122627: dataIn1 = 32'd718
; 
32'd122628: dataIn1 = 32'd1386
; 
32'd122629: dataIn1 = 32'd1388
; 
32'd122630: dataIn1 = 32'd11245
; 
32'd122631: dataIn1 = 32'd11246
; 
32'd122632: dataIn1 = 32'd11247
; 
32'd122633: dataIn1 = 32'd362
; 
32'd122634: dataIn1 = 32'd372
; 
32'd122635: dataIn1 = 32'd716
; 
32'd122636: dataIn1 = 32'd717
; 
32'd122637: dataIn1 = 32'd718
; 
32'd122638: dataIn1 = 32'd1386
; 
32'd122639: dataIn1 = 32'd5616
; 
32'd122640: dataIn1 = 32'd5617
; 
32'd122641: dataIn1 = 32'd369
; 
32'd122642: dataIn1 = 32'd374
; 
32'd122643: dataIn1 = 32'd719
; 
32'd122644: dataIn1 = 32'd720
; 
32'd122645: dataIn1 = 32'd721
; 
32'd122646: dataIn1 = 32'd1389
; 
32'd122647: dataIn1 = 32'd5624
; 
32'd122648: dataIn1 = 32'd5625
; 
32'd122649: dataIn1 = 32'd374
; 
32'd122650: dataIn1 = 32'd719
; 
32'd122651: dataIn1 = 32'd720
; 
32'd122652: dataIn1 = 32'd1389
; 
32'd122653: dataIn1 = 32'd1390
; 
32'd122654: dataIn1 = 32'd11210
; 
32'd122655: dataIn1 = 32'd11211
; 
32'd122656: dataIn1 = 32'd11212
; 
32'd122657: dataIn1 = 32'd369
; 
32'd122658: dataIn1 = 32'd719
; 
32'd122659: dataIn1 = 32'd721
; 
32'd122660: dataIn1 = 32'd1389
; 
32'd122661: dataIn1 = 32'd1391
; 
32'd122662: dataIn1 = 32'd11213
; 
32'd122663: dataIn1 = 32'd11214
; 
32'd122664: dataIn1 = 32'd11215
; 
32'd122665: dataIn1 = 32'd11216
; 
32'd122666: dataIn1 = 32'd374
; 
32'd122667: dataIn1 = 32'd722
; 
32'd122668: dataIn1 = 32'd730
; 
32'd122669: dataIn1 = 32'd1390
; 
32'd122670: dataIn1 = 32'd1396
; 
32'd122671: dataIn1 = 32'd11206
; 
32'd122672: dataIn1 = 32'd11207
; 
32'd122673: dataIn1 = 32'd11208
; 
32'd122674: dataIn1 = 32'd376
; 
32'd122675: dataIn1 = 32'd377
; 
32'd122676: dataIn1 = 32'd723
; 
32'd122677: dataIn1 = 32'd724
; 
32'd122678: dataIn1 = 32'd1392
; 
32'd122679: dataIn1 = 32'd1393
; 
32'd122680: dataIn1 = 32'd5628
; 
32'd122681: dataIn1 = 32'd5629
; 
32'd122682: dataIn1 = 32'd723
; 
32'd122683: dataIn1 = 32'd724
; 
32'd122684: dataIn1 = 32'd1392
; 
32'd122685: dataIn1 = 32'd1393
; 
32'd122686: dataIn1 = 32'd11203
; 
32'd122687: dataIn1 = 32'd11204
; 
32'd122688: dataIn1 = 32'd376
; 
32'd122689: dataIn1 = 32'd725
; 
32'd122690: dataIn1 = 32'd1392
; 
32'd122691: dataIn1 = 32'd1394
; 
32'd122692: dataIn1 = 32'd11201
; 
32'd122693: dataIn1 = 32'd11202
; 
32'd122694: dataIn1 = 32'd377
; 
32'd122695: dataIn1 = 32'd726
; 
32'd122696: dataIn1 = 32'd1393
; 
32'd122697: dataIn1 = 32'd1396
; 
32'd122698: dataIn1 = 32'd11205
; 
32'd122699: dataIn1 = 32'd11206
; 
32'd122700: dataIn1 = 32'd727
; 
32'd122701: dataIn1 = 32'd729
; 
32'd122702: dataIn1 = 32'd1394
; 
32'd122703: dataIn1 = 32'd1395
; 
32'd122704: dataIn1 = 32'd11198
; 
32'd122705: dataIn1 = 32'd11199
; 
32'd122706: dataIn1 = 32'd378
; 
32'd122707: dataIn1 = 32'd728
; 
32'd122708: dataIn1 = 32'd1395
; 
32'd122709: dataIn1 = 32'd10563
; 
32'd122710: dataIn1 = 32'd376
; 
32'd122711: dataIn1 = 32'd378
; 
32'd122712: dataIn1 = 32'd727
; 
32'd122713: dataIn1 = 32'd729
; 
32'd122714: dataIn1 = 32'd1394
; 
32'd122715: dataIn1 = 32'd1395
; 
32'd122716: dataIn1 = 32'd5630
; 
32'd122717: dataIn1 = 32'd5631
; 
32'd122718: dataIn1 = 32'd374
; 
32'd122719: dataIn1 = 32'd377
; 
32'd122720: dataIn1 = 32'd722
; 
32'd122721: dataIn1 = 32'd730
; 
32'd122722: dataIn1 = 32'd1396
; 
32'd122723: dataIn1 = 32'd5626
; 
32'd122724: dataIn1 = 32'd5627
; 
32'd122725: dataIn1 = 32'd731
; 
32'd122726: dataIn1 = 32'd1397
; 
32'd122727: dataIn1 = 32'd1398
; 
32'd122728: dataIn1 = 32'd1829
; 
32'd122729: dataIn1 = 32'd10750
; 
32'd122730: dataIn1 = 32'd10751
; 
32'd122731: dataIn1 = 32'd732
; 
32'd122732: dataIn1 = 32'd1399
; 
32'd122733: dataIn1 = 32'd1400
; 
32'd122734: dataIn1 = 32'd1831
; 
32'd122735: dataIn1 = 32'd10746
; 
32'd122736: dataIn1 = 32'd10747
; 
32'd122737: dataIn1 = 32'd733
; 
32'd122738: dataIn1 = 32'd1401
; 
32'd122739: dataIn1 = 32'd1402
; 
32'd122740: dataIn1 = 32'd1834
; 
32'd122741: dataIn1 = 32'd10754
; 
32'd122742: dataIn1 = 32'd10755
; 
32'd122743: dataIn1 = 32'd734
; 
32'd122744: dataIn1 = 32'd1403
; 
32'd122745: dataIn1 = 32'd1404
; 
32'd122746: dataIn1 = 32'd1835
; 
32'd122747: dataIn1 = 32'd10759
; 
32'd122748: dataIn1 = 32'd10760
; 
32'd122749: dataIn1 = 32'd735
; 
32'd122750: dataIn1 = 32'd1405
; 
32'd122751: dataIn1 = 32'd1406
; 
32'd122752: dataIn1 = 32'd1837
; 
32'd122753: dataIn1 = 32'd10738
; 
32'd122754: dataIn1 = 32'd10739
; 
32'd122755: dataIn1 = 32'd736
; 
32'd122756: dataIn1 = 32'd1407
; 
32'd122757: dataIn1 = 32'd1408
; 
32'd122758: dataIn1 = 32'd1840
; 
32'd122759: dataIn1 = 32'd10742
; 
32'd122760: dataIn1 = 32'd10743
; 
32'd122761: dataIn1 = 32'd737
; 
32'd122762: dataIn1 = 32'd1409
; 
32'd122763: dataIn1 = 32'd1410
; 
32'd122764: dataIn1 = 32'd1841
; 
32'd122765: dataIn1 = 32'd1842
; 
32'd122766: dataIn1 = 32'd10734
; 
32'd122767: dataIn1 = 32'd10735
; 
32'd122768: dataIn1 = 32'd738
; 
32'd122769: dataIn1 = 32'd1411
; 
32'd122770: dataIn1 = 32'd1412
; 
32'd122771: dataIn1 = 32'd1843
; 
32'd122772: dataIn1 = 32'd1844
; 
32'd122773: dataIn1 = 32'd10730
; 
32'd122774: dataIn1 = 32'd10731
; 
32'd122775: dataIn1 = 32'd739
; 
32'd122776: dataIn1 = 32'd1413
; 
32'd122777: dataIn1 = 32'd1414
; 
32'd122778: dataIn1 = 32'd1845
; 
32'd122779: dataIn1 = 32'd1846
; 
32'd122780: dataIn1 = 32'd10718
; 
32'd122781: dataIn1 = 32'd10719
; 
32'd122782: dataIn1 = 32'd740
; 
32'd122783: dataIn1 = 32'd1415
; 
32'd122784: dataIn1 = 32'd1416
; 
32'd122785: dataIn1 = 32'd1848
; 
32'd122786: dataIn1 = 32'd3446
; 
32'd122787: dataIn1 = 32'd10714
; 
32'd122788: dataIn1 = 32'd10715
; 
32'd122789: dataIn1 = 32'd741
; 
32'd122790: dataIn1 = 32'd1417
; 
32'd122791: dataIn1 = 32'd1418
; 
32'd122792: dataIn1 = 32'd1849
; 
32'd122793: dataIn1 = 32'd1850
; 
32'd122794: dataIn1 = 32'd10722
; 
32'd122795: dataIn1 = 32'd10723
; 
32'd122796: dataIn1 = 32'd742
; 
32'd122797: dataIn1 = 32'd1419
; 
32'd122798: dataIn1 = 32'd1420
; 
32'd122799: dataIn1 = 32'd1851
; 
32'd122800: dataIn1 = 32'd1852
; 
32'd122801: dataIn1 = 32'd10726
; 
32'd122802: dataIn1 = 32'd10727
; 
32'd122803: dataIn1 = 32'd743
; 
32'd122804: dataIn1 = 32'd1421
; 
32'd122805: dataIn1 = 32'd1424
; 
32'd122806: dataIn1 = 32'd3462
; 
32'd122807: dataIn1 = 32'd10707
; 
32'd122808: dataIn1 = 32'd11737
; 
32'd122809: dataIn1 = 32'd11738
; 
32'd122810: dataIn1 = 32'd744
; 
32'd122811: dataIn1 = 32'd750
; 
32'd122812: dataIn1 = 32'd1423
; 
32'd122813: dataIn1 = 32'd1432
; 
32'd122814: dataIn1 = 32'd11732
; 
32'd122815: dataIn1 = 32'd11733
; 
32'd122816: dataIn1 = 32'd11734
; 
32'd122817: dataIn1 = 32'd745
; 
32'd122818: dataIn1 = 32'd2041
; 
32'd122819: dataIn1 = 32'd3415
; 
32'd122820: dataIn1 = 32'd3416
; 
32'd122821: dataIn1 = 32'd3448
; 
32'd122822: dataIn1 = 32'd3462
; 
32'd122823: dataIn1 = 32'd3470
; 
32'd122824: dataIn1 = 32'd746
; 
32'd122825: dataIn1 = 32'd1424
; 
32'd122826: dataIn1 = 32'd1430
; 
32'd122827: dataIn1 = 32'd3448
; 
32'd122828: dataIn1 = 32'd10555
; 
32'd122829: dataIn1 = 32'd10556
; 
32'd122830: dataIn1 = 32'd10557
; 
32'd122831: dataIn1 = 32'd10558
; 
32'd122832: dataIn1 = 32'd10559
; 
32'd122833: dataIn1 = 32'd10560
; 
32'd122834: dataIn1 = 32'd747
; 
32'd122835: dataIn1 = 32'd1425
; 
32'd122836: dataIn1 = 32'd1426
; 
32'd122837: dataIn1 = 32'd3027
; 
32'd122838: dataIn1 = 32'd3029
; 
32'd122839: dataIn1 = 32'd10710
; 
32'd122840: dataIn1 = 32'd10711
; 
32'd122841: dataIn1 = 32'd392
; 
32'd122842: dataIn1 = 32'd748
; 
32'd122843: dataIn1 = 32'd761
; 
32'd122844: dataIn1 = 32'd1427
; 
32'd122845: dataIn1 = 32'd1428
; 
32'd122846: dataIn1 = 32'd1431
; 
32'd122847: dataIn1 = 32'd1450
; 
32'd122848: dataIn1 = 32'd392
; 
32'd122849: dataIn1 = 32'd749
; 
32'd122850: dataIn1 = 32'd1428
; 
32'd122851: dataIn1 = 32'd1429
; 
32'd122852: dataIn1 = 32'd3460
; 
32'd122853: dataIn1 = 32'd10271
; 
32'd122854: dataIn1 = 32'd10558
; 
32'd122855: dataIn1 = 32'd266
; 
32'd122856: dataIn1 = 32'd390
; 
32'd122857: dataIn1 = 32'd549
; 
32'd122858: dataIn1 = 32'd744
; 
32'd122859: dataIn1 = 32'd750
; 
32'd122860: dataIn1 = 32'd1423
; 
32'd122861: dataIn1 = 32'd1432
; 
32'd122862: dataIn1 = 32'd2041
; 
32'd122863: dataIn1 = 32'd2042
; 
32'd122864: dataIn1 = 32'd395
; 
32'd122865: dataIn1 = 32'd396
; 
32'd122866: dataIn1 = 32'd751
; 
32'd122867: dataIn1 = 32'd752
; 
32'd122868: dataIn1 = 32'd753
; 
32'd122869: dataIn1 = 32'd1433
; 
32'd122870: dataIn1 = 32'd4602
; 
32'd122871: dataIn1 = 32'd5426
; 
32'd122872: dataIn1 = 32'd396
; 
32'd122873: dataIn1 = 32'd751
; 
32'd122874: dataIn1 = 32'd752
; 
32'd122875: dataIn1 = 32'd1433
; 
32'd122876: dataIn1 = 32'd1435
; 
32'd122877: dataIn1 = 32'd1436
; 
32'd122878: dataIn1 = 32'd1438
; 
32'd122879: dataIn1 = 32'd395
; 
32'd122880: dataIn1 = 32'd751
; 
32'd122881: dataIn1 = 32'd753
; 
32'd122882: dataIn1 = 32'd1433
; 
32'd122883: dataIn1 = 32'd1434
; 
32'd122884: dataIn1 = 32'd1442
; 
32'd122885: dataIn1 = 32'd1443
; 
32'd122886: dataIn1 = 32'd396
; 
32'd122887: dataIn1 = 32'd754
; 
32'd122888: dataIn1 = 32'd761
; 
32'd122889: dataIn1 = 32'd1437
; 
32'd122890: dataIn1 = 32'd1438
; 
32'd122891: dataIn1 = 32'd1441
; 
32'd122892: dataIn1 = 32'd1450
; 
32'd122893: dataIn1 = 32'd755
; 
32'd122894: dataIn1 = 32'd1439
; 
32'd122895: dataIn1 = 32'd1440
; 
32'd122896: dataIn1 = 32'd3032
; 
32'd122897: dataIn1 = 32'd3033
; 
32'd122898: dataIn1 = 32'd10548
; 
32'd122899: dataIn1 = 32'd10549
; 
32'd122900: dataIn1 = 32'd10550
; 
32'd122901: dataIn1 = 32'd395
; 
32'd122902: dataIn1 = 32'd756
; 
32'd122903: dataIn1 = 32'd760
; 
32'd122904: dataIn1 = 32'd1443
; 
32'd122905: dataIn1 = 32'd1444
; 
32'd122906: dataIn1 = 32'd1446
; 
32'd122907: dataIn1 = 32'd1449
; 
32'd122908: dataIn1 = 32'd757
; 
32'd122909: dataIn1 = 32'd1445
; 
32'd122910: dataIn1 = 32'd1447
; 
32'd122911: dataIn1 = 32'd3447
; 
32'd122912: dataIn1 = 32'd10539
; 
32'd122913: dataIn1 = 32'd10540
; 
32'd122914: dataIn1 = 32'd10541
; 
32'd122915: dataIn1 = 32'd10542
; 
32'd122916: dataIn1 = 32'd10675
; 
32'd122917: dataIn1 = 32'd758
; 
32'd122918: dataIn1 = 32'd3411
; 
32'd122919: dataIn1 = 32'd3412
; 
32'd122920: dataIn1 = 32'd3447
; 
32'd122921: dataIn1 = 32'd3461
; 
32'd122922: dataIn1 = 32'd3469
; 
32'd122923: dataIn1 = 32'd10258
; 
32'd122924: dataIn1 = 32'd398
; 
32'd122925: dataIn1 = 32'd759
; 
32'd122926: dataIn1 = 32'd760
; 
32'd122927: dataIn1 = 32'd1448
; 
32'd122928: dataIn1 = 32'd1449
; 
32'd122929: dataIn1 = 32'd1478
; 
32'd122930: dataIn1 = 32'd1479
; 
32'd122931: dataIn1 = 32'd395
; 
32'd122932: dataIn1 = 32'd398
; 
32'd122933: dataIn1 = 32'd756
; 
32'd122934: dataIn1 = 32'd759
; 
32'd122935: dataIn1 = 32'd760
; 
32'd122936: dataIn1 = 32'd1449
; 
32'd122937: dataIn1 = 32'd5509
; 
32'd122938: dataIn1 = 32'd5510
; 
32'd122939: dataIn1 = 32'd392
; 
32'd122940: dataIn1 = 32'd396
; 
32'd122941: dataIn1 = 32'd748
; 
32'd122942: dataIn1 = 32'd754
; 
32'd122943: dataIn1 = 32'd761
; 
32'd122944: dataIn1 = 32'd1450
; 
32'd122945: dataIn1 = 32'd2289
; 
32'd122946: dataIn1 = 32'd2489
; 
32'd122947: dataIn1 = 32'd403
; 
32'd122948: dataIn1 = 32'd762
; 
32'd122949: dataIn1 = 32'd763
; 
32'd122950: dataIn1 = 32'd1452
; 
32'd122951: dataIn1 = 32'd1453
; 
32'd122952: dataIn1 = 32'd1455
; 
32'd122953: dataIn1 = 32'd1456
; 
32'd122954: dataIn1 = 32'd401
; 
32'd122955: dataIn1 = 32'd403
; 
32'd122956: dataIn1 = 32'd762
; 
32'd122957: dataIn1 = 32'd763
; 
32'd122958: dataIn1 = 32'd764
; 
32'd122959: dataIn1 = 32'd1452
; 
32'd122960: dataIn1 = 32'd2290
; 
32'd122961: dataIn1 = 32'd2291
; 
32'd122962: dataIn1 = 32'd401
; 
32'd122963: dataIn1 = 32'd763
; 
32'd122964: dataIn1 = 32'd764
; 
32'd122965: dataIn1 = 32'd767
; 
32'd122966: dataIn1 = 32'd1451
; 
32'd122967: dataIn1 = 32'd1452
; 
32'd122968: dataIn1 = 32'd1459
; 
32'd122969: dataIn1 = 32'd403
; 
32'd122970: dataIn1 = 32'd765
; 
32'd122971: dataIn1 = 32'd769
; 
32'd122972: dataIn1 = 32'd1454
; 
32'd122973: dataIn1 = 32'd1456
; 
32'd122974: dataIn1 = 32'd1457
; 
32'd122975: dataIn1 = 32'd1464
; 
32'd122976: dataIn1 = 32'd766
; 
32'd122977: dataIn1 = 32'd767
; 
32'd122978: dataIn1 = 32'd1459
; 
32'd122979: dataIn1 = 32'd1463
; 
32'd122980: dataIn1 = 32'd10526
; 
32'd122981: dataIn1 = 32'd10527
; 
32'd122982: dataIn1 = 32'd10528
; 
32'd122983: dataIn1 = 32'd10529
; 
32'd122984: dataIn1 = 32'd10684
; 
32'd122985: dataIn1 = 32'd207
; 
32'd122986: dataIn1 = 32'd401
; 
32'd122987: dataIn1 = 32'd764
; 
32'd122988: dataIn1 = 32'd766
; 
32'd122989: dataIn1 = 32'd767
; 
32'd122990: dataIn1 = 32'd1459
; 
32'd122991: dataIn1 = 32'd1463
; 
32'd122992: dataIn1 = 32'd1862
; 
32'd122993: dataIn1 = 32'd2045
; 
32'd122994: dataIn1 = 32'd768
; 
32'd122995: dataIn1 = 32'd1461
; 
32'd122996: dataIn1 = 32'd1462
; 
32'd122997: dataIn1 = 32'd1490
; 
32'd122998: dataIn1 = 32'd2758
; 
32'd122999: dataIn1 = 32'd10525
; 
32'd123000: dataIn1 = 32'd10526
; 
32'd123001: dataIn1 = 32'd403
; 
32'd123002: dataIn1 = 32'd405
; 
32'd123003: dataIn1 = 32'd765
; 
32'd123004: dataIn1 = 32'd769
; 
32'd123005: dataIn1 = 32'd770
; 
32'd123006: dataIn1 = 32'd1464
; 
32'd123007: dataIn1 = 32'd2292
; 
32'd123008: dataIn1 = 32'd2490
; 
32'd123009: dataIn1 = 32'd405
; 
32'd123010: dataIn1 = 32'd769
; 
32'd123011: dataIn1 = 32'd770
; 
32'd123012: dataIn1 = 32'd1464
; 
32'd123013: dataIn1 = 32'd1465
; 
32'd123014: dataIn1 = 32'd1475
; 
32'd123015: dataIn1 = 32'd1476
; 
32'd123016: dataIn1 = 32'd771
; 
32'd123017: dataIn1 = 32'd1467
; 
32'd123018: dataIn1 = 32'd1468
; 
32'd123019: dataIn1 = 32'd1469
; 
32'd123020: dataIn1 = 32'd1470
; 
32'd123021: dataIn1 = 32'd1859
; 
32'd123022: dataIn1 = 32'd10284
; 
32'd123023: dataIn1 = 32'd405
; 
32'd123024: dataIn1 = 32'd772
; 
32'd123025: dataIn1 = 32'd774
; 
32'd123026: dataIn1 = 32'd1473
; 
32'd123027: dataIn1 = 32'd1474
; 
32'd123028: dataIn1 = 32'd1476
; 
32'd123029: dataIn1 = 32'd1477
; 
32'd123030: dataIn1 = 32'd398
; 
32'd123031: dataIn1 = 32'd773
; 
32'd123032: dataIn1 = 32'd774
; 
32'd123033: dataIn1 = 32'd1472
; 
32'd123034: dataIn1 = 32'd1474
; 
32'd123035: dataIn1 = 32'd1478
; 
32'd123036: dataIn1 = 32'd1480
; 
32'd123037: dataIn1 = 32'd398
; 
32'd123038: dataIn1 = 32'd405
; 
32'd123039: dataIn1 = 32'd772
; 
32'd123040: dataIn1 = 32'd773
; 
32'd123041: dataIn1 = 32'd774
; 
32'd123042: dataIn1 = 32'd1474
; 
32'd123043: dataIn1 = 32'd4603
; 
32'd123044: dataIn1 = 32'd5427
; 
32'd123045: dataIn1 = 32'd775
; 
32'd123046: dataIn1 = 32'd2492
; 
32'd123047: dataIn1 = 32'd2493
; 
32'd123048: dataIn1 = 32'd2495
; 
32'd123049: dataIn1 = 32'd2496
; 
32'd123050: dataIn1 = 32'd3422
; 
32'd123051: dataIn1 = 32'd3423
; 
32'd123052: dataIn1 = 32'd776
; 
32'd123053: dataIn1 = 32'd1481
; 
32'd123054: dataIn1 = 32'd1482
; 
32'd123055: dataIn1 = 32'd2494
; 
32'd123056: dataIn1 = 32'd2496
; 
32'd123057: dataIn1 = 32'd10519
; 
32'd123058: dataIn1 = 32'd10520
; 
32'd123059: dataIn1 = 32'd777
; 
32'd123060: dataIn1 = 32'd1481
; 
32'd123061: dataIn1 = 32'd1485
; 
32'd123062: dataIn1 = 32'd2491
; 
32'd123063: dataIn1 = 32'd2492
; 
32'd123064: dataIn1 = 32'd10521
; 
32'd123065: dataIn1 = 32'd10522
; 
32'd123066: dataIn1 = 32'd778
; 
32'd123067: dataIn1 = 32'd1482
; 
32'd123068: dataIn1 = 32'd1491
; 
32'd123069: dataIn1 = 32'd2504
; 
32'd123070: dataIn1 = 32'd2505
; 
32'd123071: dataIn1 = 32'd10517
; 
32'd123072: dataIn1 = 32'd10518
; 
32'd123073: dataIn1 = 32'd779
; 
32'd123074: dataIn1 = 32'd1483
; 
32'd123075: dataIn1 = 32'd1484
; 
32'd123076: dataIn1 = 32'd1860
; 
32'd123077: dataIn1 = 32'd1861
; 
32'd123078: dataIn1 = 32'd10518
; 
32'd123079: dataIn1 = 32'd10519
; 
32'd123080: dataIn1 = 32'd780
; 
32'd123081: dataIn1 = 32'd1485
; 
32'd123082: dataIn1 = 32'd1490
; 
32'd123083: dataIn1 = 32'd2498
; 
32'd123084: dataIn1 = 32'd2499
; 
32'd123085: dataIn1 = 32'd10523
; 
32'd123086: dataIn1 = 32'd10524
; 
32'd123087: dataIn1 = 32'd781
; 
32'd123088: dataIn1 = 32'd1486
; 
32'd123089: dataIn1 = 32'd1487
; 
32'd123090: dataIn1 = 32'd1862
; 
32'd123091: dataIn1 = 32'd1863
; 
32'd123092: dataIn1 = 32'd10522
; 
32'd123093: dataIn1 = 32'd10523
; 
32'd123094: dataIn1 = 32'd270
; 
32'd123095: dataIn1 = 32'd782
; 
32'd123096: dataIn1 = 32'd976
; 
32'd123097: dataIn1 = 32'd1488
; 
32'd123098: dataIn1 = 32'd1489
; 
32'd123099: dataIn1 = 32'd3459
; 
32'd123100: dataIn1 = 32'd11665
; 
32'd123101: dataIn1 = 32'd11666
; 
32'd123102: dataIn1 = 32'd783
; 
32'd123103: dataIn1 = 32'd976
; 
32'd123104: dataIn1 = 32'd2497
; 
32'd123105: dataIn1 = 32'd2498
; 
32'd123106: dataIn1 = 32'd2758
; 
32'd123107: dataIn1 = 32'd3439
; 
32'd123108: dataIn1 = 32'd3459
; 
32'd123109: dataIn1 = 32'd784
; 
32'd123110: dataIn1 = 32'd2500
; 
32'd123111: dataIn1 = 32'd2502
; 
32'd123112: dataIn1 = 32'd2503
; 
32'd123113: dataIn1 = 32'd2505
; 
32'd123114: dataIn1 = 32'd3424
; 
32'd123115: dataIn1 = 32'd3425
; 
32'd123116: dataIn1 = 32'd785
; 
32'd123117: dataIn1 = 32'd1491
; 
32'd123118: dataIn1 = 32'd1493
; 
32'd123119: dataIn1 = 32'd2500
; 
32'd123120: dataIn1 = 32'd2501
; 
32'd123121: dataIn1 = 32'd10515
; 
32'd123122: dataIn1 = 32'd10516
; 
32'd123123: dataIn1 = 32'd786
; 
32'd123124: dataIn1 = 32'd2507
; 
32'd123125: dataIn1 = 32'd2508
; 
32'd123126: dataIn1 = 32'd2510
; 
32'd123127: dataIn1 = 32'd2511
; 
32'd123128: dataIn1 = 32'd3426
; 
32'd123129: dataIn1 = 32'd3427
; 
32'd123130: dataIn1 = 32'd787
; 
32'd123131: dataIn1 = 32'd1492
; 
32'd123132: dataIn1 = 32'd1493
; 
32'd123133: dataIn1 = 32'd2509
; 
32'd123134: dataIn1 = 32'd2511
; 
32'd123135: dataIn1 = 32'd10513
; 
32'd123136: dataIn1 = 32'd10514
; 
32'd123137: dataIn1 = 32'd788
; 
32'd123138: dataIn1 = 32'd1492
; 
32'd123139: dataIn1 = 32'd1496
; 
32'd123140: dataIn1 = 32'd2506
; 
32'd123141: dataIn1 = 32'd2507
; 
32'd123142: dataIn1 = 32'd10511
; 
32'd123143: dataIn1 = 32'd10512
; 
32'd123144: dataIn1 = 32'd789
; 
32'd123145: dataIn1 = 32'd1494
; 
32'd123146: dataIn1 = 32'd1495
; 
32'd123147: dataIn1 = 32'd1864
; 
32'd123148: dataIn1 = 32'd1865
; 
32'd123149: dataIn1 = 32'd10514
; 
32'd123150: dataIn1 = 32'd10515
; 
32'd123151: dataIn1 = 32'd790
; 
32'd123152: dataIn1 = 32'd1496
; 
32'd123153: dataIn1 = 32'd1513
; 
32'd123154: dataIn1 = 32'd2519
; 
32'd123155: dataIn1 = 32'd2520
; 
32'd123156: dataIn1 = 32'd10509
; 
32'd123157: dataIn1 = 32'd10510
; 
32'd123158: dataIn1 = 32'd791
; 
32'd123159: dataIn1 = 32'd1497
; 
32'd123160: dataIn1 = 32'd1498
; 
32'd123161: dataIn1 = 32'd1866
; 
32'd123162: dataIn1 = 32'd1867
; 
32'd123163: dataIn1 = 32'd10510
; 
32'd123164: dataIn1 = 32'd10511
; 
32'd123165: dataIn1 = 32'd792
; 
32'd123166: dataIn1 = 32'd1499
; 
32'd123167: dataIn1 = 32'd1500
; 
32'd123168: dataIn1 = 32'd10497
; 
32'd123169: dataIn1 = 32'd10498
; 
32'd123170: dataIn1 = 32'd10967
; 
32'd123171: dataIn1 = 32'd10968
; 
32'd123172: dataIn1 = 32'd793
; 
32'd123173: dataIn1 = 32'd1499
; 
32'd123174: dataIn1 = 32'd1503
; 
32'd123175: dataIn1 = 32'd10495
; 
32'd123176: dataIn1 = 32'd10496
; 
32'd123177: dataIn1 = 32'd10965
; 
32'd123178: dataIn1 = 32'd10966
; 
32'd123179: dataIn1 = 32'd794
; 
32'd123180: dataIn1 = 32'd1500
; 
32'd123181: dataIn1 = 32'd1515
; 
32'd123182: dataIn1 = 32'd10499
; 
32'd123183: dataIn1 = 32'd10500
; 
32'd123184: dataIn1 = 32'd10969
; 
32'd123185: dataIn1 = 32'd10970
; 
32'd123186: dataIn1 = 32'd795
; 
32'd123187: dataIn1 = 32'd1501
; 
32'd123188: dataIn1 = 32'd1502
; 
32'd123189: dataIn1 = 32'd3035
; 
32'd123190: dataIn1 = 32'd3036
; 
32'd123191: dataIn1 = 32'd10498
; 
32'd123192: dataIn1 = 32'd10499
; 
32'd123193: dataIn1 = 32'd796
; 
32'd123194: dataIn1 = 32'd1504
; 
32'd123195: dataIn1 = 32'd1505
; 
32'd123196: dataIn1 = 32'd1870
; 
32'd123197: dataIn1 = 32'd1871
; 
32'd123198: dataIn1 = 32'd10494
; 
32'd123199: dataIn1 = 32'd10495
; 
32'd123200: dataIn1 = 32'd797
; 
32'd123201: dataIn1 = 32'd1503
; 
32'd123202: dataIn1 = 32'd1526
; 
32'd123203: dataIn1 = 32'd10493
; 
32'd123204: dataIn1 = 32'd10494
; 
32'd123205: dataIn1 = 32'd10963
; 
32'd123206: dataIn1 = 32'd10964
; 
32'd123207: dataIn1 = 32'd798
; 
32'd123208: dataIn1 = 32'd1506
; 
32'd123209: dataIn1 = 32'd1507
; 
32'd123210: dataIn1 = 32'd1872
; 
32'd123211: dataIn1 = 32'd2759
; 
32'd123212: dataIn1 = 32'd10503
; 
32'd123213: dataIn1 = 32'd10504
; 
32'd123214: dataIn1 = 32'd799
; 
32'd123215: dataIn1 = 32'd1506
; 
32'd123216: dataIn1 = 32'd1510
; 
32'd123217: dataIn1 = 32'd2512
; 
32'd123218: dataIn1 = 32'd2514
; 
32'd123219: dataIn1 = 32'd10505
; 
32'd123220: dataIn1 = 32'd10506
; 
32'd123221: dataIn1 = 32'd800
; 
32'd123222: dataIn1 = 32'd2512
; 
32'd123223: dataIn1 = 32'd2513
; 
32'd123224: dataIn1 = 32'd2759
; 
32'd123225: dataIn1 = 32'd3040
; 
32'd123226: dataIn1 = 32'd3445
; 
32'd123227: dataIn1 = 32'd10251
; 
32'd123228: dataIn1 = 32'd801
; 
32'd123229: dataIn1 = 32'd1508
; 
32'd123230: dataIn1 = 32'd1509
; 
32'd123231: dataIn1 = 32'd1873
; 
32'd123232: dataIn1 = 32'd10285
; 
32'd123233: dataIn1 = 32'd10502
; 
32'd123234: dataIn1 = 32'd10503
; 
32'd123235: dataIn1 = 32'd802
; 
32'd123236: dataIn1 = 32'd1507
; 
32'd123237: dataIn1 = 32'd1515
; 
32'd123238: dataIn1 = 32'd1516
; 
32'd123239: dataIn1 = 32'd1517
; 
32'd123240: dataIn1 = 32'd10501
; 
32'd123241: dataIn1 = 32'd10502
; 
32'd123242: dataIn1 = 32'd803
; 
32'd123243: dataIn1 = 32'd1511
; 
32'd123244: dataIn1 = 32'd1512
; 
32'd123245: dataIn1 = 32'd1875
; 
32'd123246: dataIn1 = 32'd1876
; 
32'd123247: dataIn1 = 32'd10506
; 
32'd123248: dataIn1 = 32'd10507
; 
32'd123249: dataIn1 = 32'd804
; 
32'd123250: dataIn1 = 32'd1510
; 
32'd123251: dataIn1 = 32'd1513
; 
32'd123252: dataIn1 = 32'd2515
; 
32'd123253: dataIn1 = 32'd2516
; 
32'd123254: dataIn1 = 32'd10507
; 
32'd123255: dataIn1 = 32'd10508
; 
32'd123256: dataIn1 = 32'd805
; 
32'd123257: dataIn1 = 32'd2515
; 
32'd123258: dataIn1 = 32'd2517
; 
32'd123259: dataIn1 = 32'd2518
; 
32'd123260: dataIn1 = 32'd2520
; 
32'd123261: dataIn1 = 32'd3428
; 
32'd123262: dataIn1 = 32'd3429
; 
32'd123263: dataIn1 = 32'd806
; 
32'd123264: dataIn1 = 32'd2521
; 
32'd123265: dataIn1 = 32'd2522
; 
32'd123266: dataIn1 = 32'd2760
; 
32'd123267: dataIn1 = 32'd3440
; 
32'd123268: dataIn1 = 32'd3445
; 
32'd123269: dataIn1 = 32'd10252
; 
32'd123270: dataIn1 = 32'd807
; 
32'd123271: dataIn1 = 32'd1519
; 
32'd123272: dataIn1 = 32'd1520
; 
32'd123273: dataIn1 = 32'd10487
; 
32'd123274: dataIn1 = 32'd10488
; 
32'd123275: dataIn1 = 32'd10957
; 
32'd123276: dataIn1 = 32'd10958
; 
32'd123277: dataIn1 = 32'd808
; 
32'd123278: dataIn1 = 32'd1519
; 
32'd123279: dataIn1 = 32'd1523
; 
32'd123280: dataIn1 = 32'd10489
; 
32'd123281: dataIn1 = 32'd10490
; 
32'd123282: dataIn1 = 32'd10959
; 
32'd123283: dataIn1 = 32'd10960
; 
32'd123284: dataIn1 = 32'd809
; 
32'd123285: dataIn1 = 32'd1520
; 
32'd123286: dataIn1 = 32'd1527
; 
32'd123287: dataIn1 = 32'd10485
; 
32'd123288: dataIn1 = 32'd10486
; 
32'd123289: dataIn1 = 32'd10955
; 
32'd123290: dataIn1 = 32'd10956
; 
32'd123291: dataIn1 = 32'd810
; 
32'd123292: dataIn1 = 32'd1521
; 
32'd123293: dataIn1 = 32'd1522
; 
32'd123294: dataIn1 = 32'd1877
; 
32'd123295: dataIn1 = 32'd1878
; 
32'd123296: dataIn1 = 32'd10486
; 
32'd123297: dataIn1 = 32'd10487
; 
32'd123298: dataIn1 = 32'd811
; 
32'd123299: dataIn1 = 32'd1523
; 
32'd123300: dataIn1 = 32'd1526
; 
32'd123301: dataIn1 = 32'd10491
; 
32'd123302: dataIn1 = 32'd10492
; 
32'd123303: dataIn1 = 32'd10961
; 
32'd123304: dataIn1 = 32'd10962
; 
32'd123305: dataIn1 = 32'd812
; 
32'd123306: dataIn1 = 32'd1524
; 
32'd123307: dataIn1 = 32'd1525
; 
32'd123308: dataIn1 = 32'd1879
; 
32'd123309: dataIn1 = 32'd1880
; 
32'd123310: dataIn1 = 32'd10490
; 
32'd123311: dataIn1 = 32'd10491
; 
32'd123312: dataIn1 = 32'd813
; 
32'd123313: dataIn1 = 32'd1527
; 
32'd123314: dataIn1 = 32'd1529
; 
32'd123315: dataIn1 = 32'd10483
; 
32'd123316: dataIn1 = 32'd10484
; 
32'd123317: dataIn1 = 32'd10953
; 
32'd123318: dataIn1 = 32'd10954
; 
32'd123319: dataIn1 = 32'd814
; 
32'd123320: dataIn1 = 32'd1528
; 
32'd123321: dataIn1 = 32'd1529
; 
32'd123322: dataIn1 = 32'd10481
; 
32'd123323: dataIn1 = 32'd10482
; 
32'd123324: dataIn1 = 32'd10951
; 
32'd123325: dataIn1 = 32'd10952
; 
32'd123326: dataIn1 = 32'd815
; 
32'd123327: dataIn1 = 32'd1528
; 
32'd123328: dataIn1 = 32'd1532
; 
32'd123329: dataIn1 = 32'd10479
; 
32'd123330: dataIn1 = 32'd10480
; 
32'd123331: dataIn1 = 32'd10949
; 
32'd123332: dataIn1 = 32'd10950
; 
32'd123333: dataIn1 = 32'd816
; 
32'd123334: dataIn1 = 32'd1530
; 
32'd123335: dataIn1 = 32'd1531
; 
32'd123336: dataIn1 = 32'd1881
; 
32'd123337: dataIn1 = 32'd1882
; 
32'd123338: dataIn1 = 32'd10482
; 
32'd123339: dataIn1 = 32'd10483
; 
32'd123340: dataIn1 = 32'd817
; 
32'd123341: dataIn1 = 32'd1532
; 
32'd123342: dataIn1 = 32'd1549
; 
32'd123343: dataIn1 = 32'd10477
; 
32'd123344: dataIn1 = 32'd10478
; 
32'd123345: dataIn1 = 32'd10947
; 
32'd123346: dataIn1 = 32'd10948
; 
32'd123347: dataIn1 = 32'd818
; 
32'd123348: dataIn1 = 32'd1533
; 
32'd123349: dataIn1 = 32'd1534
; 
32'd123350: dataIn1 = 32'd1883
; 
32'd123351: dataIn1 = 32'd1884
; 
32'd123352: dataIn1 = 32'd10478
; 
32'd123353: dataIn1 = 32'd10479
; 
32'd123354: dataIn1 = 32'd819
; 
32'd123355: dataIn1 = 32'd1535
; 
32'd123356: dataIn1 = 32'd1536
; 
32'd123357: dataIn1 = 32'd10465
; 
32'd123358: dataIn1 = 32'd10466
; 
32'd123359: dataIn1 = 32'd10935
; 
32'd123360: dataIn1 = 32'd10936
; 
32'd123361: dataIn1 = 32'd820
; 
32'd123362: dataIn1 = 32'd1535
; 
32'd123363: dataIn1 = 32'd1539
; 
32'd123364: dataIn1 = 32'd10463
; 
32'd123365: dataIn1 = 32'd10464
; 
32'd123366: dataIn1 = 32'd10933
; 
32'd123367: dataIn1 = 32'd10934
; 
32'd123368: dataIn1 = 32'd821
; 
32'd123369: dataIn1 = 32'd1536
; 
32'd123370: dataIn1 = 32'd1550
; 
32'd123371: dataIn1 = 32'd10467
; 
32'd123372: dataIn1 = 32'd10468
; 
32'd123373: dataIn1 = 32'd10937
; 
32'd123374: dataIn1 = 32'd10938
; 
32'd123375: dataIn1 = 32'd822
; 
32'd123376: dataIn1 = 32'd1537
; 
32'd123377: dataIn1 = 32'd1538
; 
32'd123378: dataIn1 = 32'd1885
; 
32'd123379: dataIn1 = 32'd1886
; 
32'd123380: dataIn1 = 32'd10466
; 
32'd123381: dataIn1 = 32'd10467
; 
32'd123382: dataIn1 = 32'd823
; 
32'd123383: dataIn1 = 32'd1540
; 
32'd123384: dataIn1 = 32'd1541
; 
32'd123385: dataIn1 = 32'd1887
; 
32'd123386: dataIn1 = 32'd1888
; 
32'd123387: dataIn1 = 32'd10462
; 
32'd123388: dataIn1 = 32'd10463
; 
32'd123389: dataIn1 = 32'd824
; 
32'd123390: dataIn1 = 32'd1539
; 
32'd123391: dataIn1 = 32'd1558
; 
32'd123392: dataIn1 = 32'd10461
; 
32'd123393: dataIn1 = 32'd10462
; 
32'd123394: dataIn1 = 32'd10931
; 
32'd123395: dataIn1 = 32'd10932
; 
32'd123396: dataIn1 = 32'd825
; 
32'd123397: dataIn1 = 32'd1542
; 
32'd123398: dataIn1 = 32'd1543
; 
32'd123399: dataIn1 = 32'd10471
; 
32'd123400: dataIn1 = 32'd10472
; 
32'd123401: dataIn1 = 32'd10941
; 
32'd123402: dataIn1 = 32'd10942
; 
32'd123403: dataIn1 = 32'd826
; 
32'd123404: dataIn1 = 32'd1542
; 
32'd123405: dataIn1 = 32'd1546
; 
32'd123406: dataIn1 = 32'd10473
; 
32'd123407: dataIn1 = 32'd10474
; 
32'd123408: dataIn1 = 32'd10943
; 
32'd123409: dataIn1 = 32'd10944
; 
32'd123410: dataIn1 = 32'd827
; 
32'd123411: dataIn1 = 32'd1544
; 
32'd123412: dataIn1 = 32'd1545
; 
32'd123413: dataIn1 = 32'd1889
; 
32'd123414: dataIn1 = 32'd1890
; 
32'd123415: dataIn1 = 32'd10470
; 
32'd123416: dataIn1 = 32'd10471
; 
32'd123417: dataIn1 = 32'd828
; 
32'd123418: dataIn1 = 32'd1543
; 
32'd123419: dataIn1 = 32'd1550
; 
32'd123420: dataIn1 = 32'd10469
; 
32'd123421: dataIn1 = 32'd10470
; 
32'd123422: dataIn1 = 32'd10939
; 
32'd123423: dataIn1 = 32'd10940
; 
32'd123424: dataIn1 = 32'd829
; 
32'd123425: dataIn1 = 32'd1547
; 
32'd123426: dataIn1 = 32'd1548
; 
32'd123427: dataIn1 = 32'd1891
; 
32'd123428: dataIn1 = 32'd1892
; 
32'd123429: dataIn1 = 32'd10474
; 
32'd123430: dataIn1 = 32'd10475
; 
32'd123431: dataIn1 = 32'd830
; 
32'd123432: dataIn1 = 32'd1546
; 
32'd123433: dataIn1 = 32'd1549
; 
32'd123434: dataIn1 = 32'd10475
; 
32'd123435: dataIn1 = 32'd10476
; 
32'd123436: dataIn1 = 32'd10945
; 
32'd123437: dataIn1 = 32'd10946
; 
32'd123438: dataIn1 = 32'd831
; 
32'd123439: dataIn1 = 32'd1551
; 
32'd123440: dataIn1 = 32'd1552
; 
32'd123441: dataIn1 = 32'd10455
; 
32'd123442: dataIn1 = 32'd10456
; 
32'd123443: dataIn1 = 32'd10925
; 
32'd123444: dataIn1 = 32'd10926
; 
32'd123445: dataIn1 = 32'd832
; 
32'd123446: dataIn1 = 32'd1551
; 
32'd123447: dataIn1 = 32'd1555
; 
32'd123448: dataIn1 = 32'd10457
; 
32'd123449: dataIn1 = 32'd10458
; 
32'd123450: dataIn1 = 32'd10927
; 
32'd123451: dataIn1 = 32'd10928
; 
32'd123452: dataIn1 = 32'd833
; 
32'd123453: dataIn1 = 32'd1552
; 
32'd123454: dataIn1 = 32'd1559
; 
32'd123455: dataIn1 = 32'd10453
; 
32'd123456: dataIn1 = 32'd10454
; 
32'd123457: dataIn1 = 32'd10923
; 
32'd123458: dataIn1 = 32'd10924
; 
32'd123459: dataIn1 = 32'd834
; 
32'd123460: dataIn1 = 32'd1553
; 
32'd123461: dataIn1 = 32'd1554
; 
32'd123462: dataIn1 = 32'd1893
; 
32'd123463: dataIn1 = 32'd1894
; 
32'd123464: dataIn1 = 32'd10454
; 
32'd123465: dataIn1 = 32'd10455
; 
32'd123466: dataIn1 = 32'd835
; 
32'd123467: dataIn1 = 32'd1555
; 
32'd123468: dataIn1 = 32'd1558
; 
32'd123469: dataIn1 = 32'd10459
; 
32'd123470: dataIn1 = 32'd10460
; 
32'd123471: dataIn1 = 32'd10929
; 
32'd123472: dataIn1 = 32'd10930
; 
32'd123473: dataIn1 = 32'd836
; 
32'd123474: dataIn1 = 32'd1556
; 
32'd123475: dataIn1 = 32'd1557
; 
32'd123476: dataIn1 = 32'd1895
; 
32'd123477: dataIn1 = 32'd1896
; 
32'd123478: dataIn1 = 32'd10458
; 
32'd123479: dataIn1 = 32'd10459
; 
32'd123480: dataIn1 = 32'd837
; 
32'd123481: dataIn1 = 32'd1559
; 
32'd123482: dataIn1 = 32'd1561
; 
32'd123483: dataIn1 = 32'd10451
; 
32'd123484: dataIn1 = 32'd10452
; 
32'd123485: dataIn1 = 32'd10921
; 
32'd123486: dataIn1 = 32'd10922
; 
32'd123487: dataIn1 = 32'd838
; 
32'd123488: dataIn1 = 32'd1560
; 
32'd123489: dataIn1 = 32'd1561
; 
32'd123490: dataIn1 = 32'd10449
; 
32'd123491: dataIn1 = 32'd10450
; 
32'd123492: dataIn1 = 32'd10919
; 
32'd123493: dataIn1 = 32'd10920
; 
32'd123494: dataIn1 = 32'd839
; 
32'd123495: dataIn1 = 32'd1560
; 
32'd123496: dataIn1 = 32'd1564
; 
32'd123497: dataIn1 = 32'd10447
; 
32'd123498: dataIn1 = 32'd10448
; 
32'd123499: dataIn1 = 32'd10917
; 
32'd123500: dataIn1 = 32'd10918
; 
32'd123501: dataIn1 = 32'd840
; 
32'd123502: dataIn1 = 32'd1562
; 
32'd123503: dataIn1 = 32'd1563
; 
32'd123504: dataIn1 = 32'd1897
; 
32'd123505: dataIn1 = 32'd1898
; 
32'd123506: dataIn1 = 32'd10450
; 
32'd123507: dataIn1 = 32'd10451
; 
32'd123508: dataIn1 = 32'd841
; 
32'd123509: dataIn1 = 32'd1564
; 
32'd123510: dataIn1 = 32'd1581
; 
32'd123511: dataIn1 = 32'd10445
; 
32'd123512: dataIn1 = 32'd10446
; 
32'd123513: dataIn1 = 32'd10915
; 
32'd123514: dataIn1 = 32'd10916
; 
32'd123515: dataIn1 = 32'd842
; 
32'd123516: dataIn1 = 32'd1565
; 
32'd123517: dataIn1 = 32'd1566
; 
32'd123518: dataIn1 = 32'd1899
; 
32'd123519: dataIn1 = 32'd1900
; 
32'd123520: dataIn1 = 32'd10446
; 
32'd123521: dataIn1 = 32'd10447
; 
32'd123522: dataIn1 = 32'd843
; 
32'd123523: dataIn1 = 32'd1567
; 
32'd123524: dataIn1 = 32'd1568
; 
32'd123525: dataIn1 = 32'd10433
; 
32'd123526: dataIn1 = 32'd10434
; 
32'd123527: dataIn1 = 32'd10903
; 
32'd123528: dataIn1 = 32'd10904
; 
32'd123529: dataIn1 = 32'd844
; 
32'd123530: dataIn1 = 32'd1567
; 
32'd123531: dataIn1 = 32'd1571
; 
32'd123532: dataIn1 = 32'd10431
; 
32'd123533: dataIn1 = 32'd10432
; 
32'd123534: dataIn1 = 32'd10901
; 
32'd123535: dataIn1 = 32'd10902
; 
32'd123536: dataIn1 = 32'd845
; 
32'd123537: dataIn1 = 32'd1568
; 
32'd123538: dataIn1 = 32'd1582
; 
32'd123539: dataIn1 = 32'd10435
; 
32'd123540: dataIn1 = 32'd10436
; 
32'd123541: dataIn1 = 32'd10905
; 
32'd123542: dataIn1 = 32'd10906
; 
32'd123543: dataIn1 = 32'd846
; 
32'd123544: dataIn1 = 32'd1569
; 
32'd123545: dataIn1 = 32'd1570
; 
32'd123546: dataIn1 = 32'd1901
; 
32'd123547: dataIn1 = 32'd1902
; 
32'd123548: dataIn1 = 32'd10434
; 
32'd123549: dataIn1 = 32'd10435
; 
32'd123550: dataIn1 = 32'd847
; 
32'd123551: dataIn1 = 32'd1572
; 
32'd123552: dataIn1 = 32'd1573
; 
32'd123553: dataIn1 = 32'd1903
; 
32'd123554: dataIn1 = 32'd1904
; 
32'd123555: dataIn1 = 32'd10430
; 
32'd123556: dataIn1 = 32'd10431
; 
32'd123557: dataIn1 = 32'd848
; 
32'd123558: dataIn1 = 32'd1571
; 
32'd123559: dataIn1 = 32'd1590
; 
32'd123560: dataIn1 = 32'd10429
; 
32'd123561: dataIn1 = 32'd10430
; 
32'd123562: dataIn1 = 32'd10899
; 
32'd123563: dataIn1 = 32'd10900
; 
32'd123564: dataIn1 = 32'd849
; 
32'd123565: dataIn1 = 32'd1574
; 
32'd123566: dataIn1 = 32'd1575
; 
32'd123567: dataIn1 = 32'd10439
; 
32'd123568: dataIn1 = 32'd10440
; 
32'd123569: dataIn1 = 32'd10909
; 
32'd123570: dataIn1 = 32'd10910
; 
32'd123571: dataIn1 = 32'd850
; 
32'd123572: dataIn1 = 32'd1574
; 
32'd123573: dataIn1 = 32'd1578
; 
32'd123574: dataIn1 = 32'd10441
; 
32'd123575: dataIn1 = 32'd10442
; 
32'd123576: dataIn1 = 32'd10911
; 
32'd123577: dataIn1 = 32'd10912
; 
32'd123578: dataIn1 = 32'd851
; 
32'd123579: dataIn1 = 32'd1576
; 
32'd123580: dataIn1 = 32'd1577
; 
32'd123581: dataIn1 = 32'd1905
; 
32'd123582: dataIn1 = 32'd1906
; 
32'd123583: dataIn1 = 32'd10438
; 
32'd123584: dataIn1 = 32'd10439
; 
32'd123585: dataIn1 = 32'd852
; 
32'd123586: dataIn1 = 32'd1575
; 
32'd123587: dataIn1 = 32'd1582
; 
32'd123588: dataIn1 = 32'd10437
; 
32'd123589: dataIn1 = 32'd10438
; 
32'd123590: dataIn1 = 32'd10907
; 
32'd123591: dataIn1 = 32'd10908
; 
32'd123592: dataIn1 = 32'd853
; 
32'd123593: dataIn1 = 32'd1579
; 
32'd123594: dataIn1 = 32'd1580
; 
32'd123595: dataIn1 = 32'd1907
; 
32'd123596: dataIn1 = 32'd1908
; 
32'd123597: dataIn1 = 32'd10442
; 
32'd123598: dataIn1 = 32'd10443
; 
32'd123599: dataIn1 = 32'd854
; 
32'd123600: dataIn1 = 32'd1578
; 
32'd123601: dataIn1 = 32'd1581
; 
32'd123602: dataIn1 = 32'd10443
; 
32'd123603: dataIn1 = 32'd10444
; 
32'd123604: dataIn1 = 32'd10913
; 
32'd123605: dataIn1 = 32'd10914
; 
32'd123606: dataIn1 = 32'd855
; 
32'd123607: dataIn1 = 32'd1583
; 
32'd123608: dataIn1 = 32'd1584
; 
32'd123609: dataIn1 = 32'd10423
; 
32'd123610: dataIn1 = 32'd10424
; 
32'd123611: dataIn1 = 32'd10893
; 
32'd123612: dataIn1 = 32'd10894
; 
32'd123613: dataIn1 = 32'd856
; 
32'd123614: dataIn1 = 32'd1583
; 
32'd123615: dataIn1 = 32'd1587
; 
32'd123616: dataIn1 = 32'd10425
; 
32'd123617: dataIn1 = 32'd10426
; 
32'd123618: dataIn1 = 32'd10895
; 
32'd123619: dataIn1 = 32'd10896
; 
32'd123620: dataIn1 = 32'd857
; 
32'd123621: dataIn1 = 32'd1584
; 
32'd123622: dataIn1 = 32'd1591
; 
32'd123623: dataIn1 = 32'd10421
; 
32'd123624: dataIn1 = 32'd10422
; 
32'd123625: dataIn1 = 32'd10891
; 
32'd123626: dataIn1 = 32'd10892
; 
32'd123627: dataIn1 = 32'd858
; 
32'd123628: dataIn1 = 32'd1585
; 
32'd123629: dataIn1 = 32'd1586
; 
32'd123630: dataIn1 = 32'd1909
; 
32'd123631: dataIn1 = 32'd1910
; 
32'd123632: dataIn1 = 32'd10422
; 
32'd123633: dataIn1 = 32'd10423
; 
32'd123634: dataIn1 = 32'd859
; 
32'd123635: dataIn1 = 32'd1587
; 
32'd123636: dataIn1 = 32'd1590
; 
32'd123637: dataIn1 = 32'd10427
; 
32'd123638: dataIn1 = 32'd10428
; 
32'd123639: dataIn1 = 32'd10897
; 
32'd123640: dataIn1 = 32'd10898
; 
32'd123641: dataIn1 = 32'd860
; 
32'd123642: dataIn1 = 32'd1588
; 
32'd123643: dataIn1 = 32'd1589
; 
32'd123644: dataIn1 = 32'd1911
; 
32'd123645: dataIn1 = 32'd1912
; 
32'd123646: dataIn1 = 32'd10426
; 
32'd123647: dataIn1 = 32'd10427
; 
32'd123648: dataIn1 = 32'd861
; 
32'd123649: dataIn1 = 32'd1591
; 
32'd123650: dataIn1 = 32'd1593
; 
32'd123651: dataIn1 = 32'd10419
; 
32'd123652: dataIn1 = 32'd10420
; 
32'd123653: dataIn1 = 32'd10889
; 
32'd123654: dataIn1 = 32'd10890
; 
32'd123655: dataIn1 = 32'd862
; 
32'd123656: dataIn1 = 32'd1592
; 
32'd123657: dataIn1 = 32'd1593
; 
32'd123658: dataIn1 = 32'd10417
; 
32'd123659: dataIn1 = 32'd10418
; 
32'd123660: dataIn1 = 32'd10887
; 
32'd123661: dataIn1 = 32'd10888
; 
32'd123662: dataIn1 = 32'd863
; 
32'd123663: dataIn1 = 32'd1592
; 
32'd123664: dataIn1 = 32'd1596
; 
32'd123665: dataIn1 = 32'd10415
; 
32'd123666: dataIn1 = 32'd10416
; 
32'd123667: dataIn1 = 32'd10885
; 
32'd123668: dataIn1 = 32'd10886
; 
32'd123669: dataIn1 = 32'd864
; 
32'd123670: dataIn1 = 32'd1594
; 
32'd123671: dataIn1 = 32'd1595
; 
32'd123672: dataIn1 = 32'd1913
; 
32'd123673: dataIn1 = 32'd1914
; 
32'd123674: dataIn1 = 32'd10418
; 
32'd123675: dataIn1 = 32'd10419
; 
32'd123676: dataIn1 = 32'd865
; 
32'd123677: dataIn1 = 32'd1596
; 
32'd123678: dataIn1 = 32'd1613
; 
32'd123679: dataIn1 = 32'd10413
; 
32'd123680: dataIn1 = 32'd10414
; 
32'd123681: dataIn1 = 32'd10883
; 
32'd123682: dataIn1 = 32'd10884
; 
32'd123683: dataIn1 = 32'd866
; 
32'd123684: dataIn1 = 32'd1597
; 
32'd123685: dataIn1 = 32'd1598
; 
32'd123686: dataIn1 = 32'd1915
; 
32'd123687: dataIn1 = 32'd1916
; 
32'd123688: dataIn1 = 32'd10414
; 
32'd123689: dataIn1 = 32'd10415
; 
32'd123690: dataIn1 = 32'd867
; 
32'd123691: dataIn1 = 32'd1599
; 
32'd123692: dataIn1 = 32'd1600
; 
32'd123693: dataIn1 = 32'd10401
; 
32'd123694: dataIn1 = 32'd10402
; 
32'd123695: dataIn1 = 32'd10871
; 
32'd123696: dataIn1 = 32'd10872
; 
32'd123697: dataIn1 = 32'd868
; 
32'd123698: dataIn1 = 32'd1599
; 
32'd123699: dataIn1 = 32'd1603
; 
32'd123700: dataIn1 = 32'd10399
; 
32'd123701: dataIn1 = 32'd10400
; 
32'd123702: dataIn1 = 32'd10869
; 
32'd123703: dataIn1 = 32'd10870
; 
32'd123704: dataIn1 = 32'd869
; 
32'd123705: dataIn1 = 32'd1600
; 
32'd123706: dataIn1 = 32'd1614
; 
32'd123707: dataIn1 = 32'd10403
; 
32'd123708: dataIn1 = 32'd10404
; 
32'd123709: dataIn1 = 32'd10873
; 
32'd123710: dataIn1 = 32'd10874
; 
32'd123711: dataIn1 = 32'd870
; 
32'd123712: dataIn1 = 32'd1601
; 
32'd123713: dataIn1 = 32'd1602
; 
32'd123714: dataIn1 = 32'd1917
; 
32'd123715: dataIn1 = 32'd1918
; 
32'd123716: dataIn1 = 32'd10402
; 
32'd123717: dataIn1 = 32'd10403
; 
32'd123718: dataIn1 = 32'd871
; 
32'd123719: dataIn1 = 32'd1604
; 
32'd123720: dataIn1 = 32'd1605
; 
32'd123721: dataIn1 = 32'd1919
; 
32'd123722: dataIn1 = 32'd1920
; 
32'd123723: dataIn1 = 32'd10398
; 
32'd123724: dataIn1 = 32'd10399
; 
32'd123725: dataIn1 = 32'd872
; 
32'd123726: dataIn1 = 32'd1603
; 
32'd123727: dataIn1 = 32'd1622
; 
32'd123728: dataIn1 = 32'd10397
; 
32'd123729: dataIn1 = 32'd10398
; 
32'd123730: dataIn1 = 32'd10867
; 
32'd123731: dataIn1 = 32'd10868
; 
32'd123732: dataIn1 = 32'd873
; 
32'd123733: dataIn1 = 32'd1606
; 
32'd123734: dataIn1 = 32'd1607
; 
32'd123735: dataIn1 = 32'd10407
; 
32'd123736: dataIn1 = 32'd10408
; 
32'd123737: dataIn1 = 32'd10877
; 
32'd123738: dataIn1 = 32'd10878
; 
32'd123739: dataIn1 = 32'd874
; 
32'd123740: dataIn1 = 32'd1606
; 
32'd123741: dataIn1 = 32'd1610
; 
32'd123742: dataIn1 = 32'd10409
; 
32'd123743: dataIn1 = 32'd10410
; 
32'd123744: dataIn1 = 32'd10879
; 
32'd123745: dataIn1 = 32'd10880
; 
32'd123746: dataIn1 = 32'd875
; 
32'd123747: dataIn1 = 32'd1608
; 
32'd123748: dataIn1 = 32'd1609
; 
32'd123749: dataIn1 = 32'd1921
; 
32'd123750: dataIn1 = 32'd1922
; 
32'd123751: dataIn1 = 32'd10406
; 
32'd123752: dataIn1 = 32'd10407
; 
32'd123753: dataIn1 = 32'd876
; 
32'd123754: dataIn1 = 32'd1607
; 
32'd123755: dataIn1 = 32'd1614
; 
32'd123756: dataIn1 = 32'd10405
; 
32'd123757: dataIn1 = 32'd10406
; 
32'd123758: dataIn1 = 32'd10875
; 
32'd123759: dataIn1 = 32'd10876
; 
32'd123760: dataIn1 = 32'd877
; 
32'd123761: dataIn1 = 32'd1611
; 
32'd123762: dataIn1 = 32'd1612
; 
32'd123763: dataIn1 = 32'd1923
; 
32'd123764: dataIn1 = 32'd1924
; 
32'd123765: dataIn1 = 32'd10410
; 
32'd123766: dataIn1 = 32'd10411
; 
32'd123767: dataIn1 = 32'd878
; 
32'd123768: dataIn1 = 32'd1610
; 
32'd123769: dataIn1 = 32'd1613
; 
32'd123770: dataIn1 = 32'd10411
; 
32'd123771: dataIn1 = 32'd10412
; 
32'd123772: dataIn1 = 32'd10881
; 
32'd123773: dataIn1 = 32'd10882
; 
32'd123774: dataIn1 = 32'd879
; 
32'd123775: dataIn1 = 32'd1615
; 
32'd123776: dataIn1 = 32'd1616
; 
32'd123777: dataIn1 = 32'd10391
; 
32'd123778: dataIn1 = 32'd10392
; 
32'd123779: dataIn1 = 32'd10861
; 
32'd123780: dataIn1 = 32'd10862
; 
32'd123781: dataIn1 = 32'd880
; 
32'd123782: dataIn1 = 32'd1615
; 
32'd123783: dataIn1 = 32'd1619
; 
32'd123784: dataIn1 = 32'd10393
; 
32'd123785: dataIn1 = 32'd10394
; 
32'd123786: dataIn1 = 32'd10863
; 
32'd123787: dataIn1 = 32'd10864
; 
32'd123788: dataIn1 = 32'd881
; 
32'd123789: dataIn1 = 32'd1616
; 
32'd123790: dataIn1 = 32'd1623
; 
32'd123791: dataIn1 = 32'd10389
; 
32'd123792: dataIn1 = 32'd10390
; 
32'd123793: dataIn1 = 32'd10859
; 
32'd123794: dataIn1 = 32'd10860
; 
32'd123795: dataIn1 = 32'd882
; 
32'd123796: dataIn1 = 32'd1617
; 
32'd123797: dataIn1 = 32'd1618
; 
32'd123798: dataIn1 = 32'd1925
; 
32'd123799: dataIn1 = 32'd1926
; 
32'd123800: dataIn1 = 32'd10390
; 
32'd123801: dataIn1 = 32'd10391
; 
32'd123802: dataIn1 = 32'd883
; 
32'd123803: dataIn1 = 32'd1619
; 
32'd123804: dataIn1 = 32'd1622
; 
32'd123805: dataIn1 = 32'd10395
; 
32'd123806: dataIn1 = 32'd10396
; 
32'd123807: dataIn1 = 32'd10865
; 
32'd123808: dataIn1 = 32'd10866
; 
32'd123809: dataIn1 = 32'd884
; 
32'd123810: dataIn1 = 32'd1620
; 
32'd123811: dataIn1 = 32'd1621
; 
32'd123812: dataIn1 = 32'd1927
; 
32'd123813: dataIn1 = 32'd1928
; 
32'd123814: dataIn1 = 32'd10394
; 
32'd123815: dataIn1 = 32'd10395
; 
32'd123816: dataIn1 = 32'd885
; 
32'd123817: dataIn1 = 32'd1623
; 
32'd123818: dataIn1 = 32'd1625
; 
32'd123819: dataIn1 = 32'd10387
; 
32'd123820: dataIn1 = 32'd10388
; 
32'd123821: dataIn1 = 32'd10857
; 
32'd123822: dataIn1 = 32'd10858
; 
32'd123823: dataIn1 = 32'd886
; 
32'd123824: dataIn1 = 32'd1624
; 
32'd123825: dataIn1 = 32'd1625
; 
32'd123826: dataIn1 = 32'd10385
; 
32'd123827: dataIn1 = 32'd10386
; 
32'd123828: dataIn1 = 32'd10855
; 
32'd123829: dataIn1 = 32'd10856
; 
32'd123830: dataIn1 = 32'd887
; 
32'd123831: dataIn1 = 32'd1624
; 
32'd123832: dataIn1 = 32'd1628
; 
32'd123833: dataIn1 = 32'd10383
; 
32'd123834: dataIn1 = 32'd10384
; 
32'd123835: dataIn1 = 32'd10853
; 
32'd123836: dataIn1 = 32'd10854
; 
32'd123837: dataIn1 = 32'd888
; 
32'd123838: dataIn1 = 32'd1626
; 
32'd123839: dataIn1 = 32'd1627
; 
32'd123840: dataIn1 = 32'd1929
; 
32'd123841: dataIn1 = 32'd1930
; 
32'd123842: dataIn1 = 32'd10386
; 
32'd123843: dataIn1 = 32'd10387
; 
32'd123844: dataIn1 = 32'd889
; 
32'd123845: dataIn1 = 32'd1628
; 
32'd123846: dataIn1 = 32'd1645
; 
32'd123847: dataIn1 = 32'd10381
; 
32'd123848: dataIn1 = 32'd10382
; 
32'd123849: dataIn1 = 32'd10851
; 
32'd123850: dataIn1 = 32'd10852
; 
32'd123851: dataIn1 = 32'd890
; 
32'd123852: dataIn1 = 32'd1629
; 
32'd123853: dataIn1 = 32'd1630
; 
32'd123854: dataIn1 = 32'd1931
; 
32'd123855: dataIn1 = 32'd1932
; 
32'd123856: dataIn1 = 32'd10382
; 
32'd123857: dataIn1 = 32'd10383
; 
32'd123858: dataIn1 = 32'd891
; 
32'd123859: dataIn1 = 32'd1631
; 
32'd123860: dataIn1 = 32'd1632
; 
32'd123861: dataIn1 = 32'd10369
; 
32'd123862: dataIn1 = 32'd10370
; 
32'd123863: dataIn1 = 32'd10839
; 
32'd123864: dataIn1 = 32'd10840
; 
32'd123865: dataIn1 = 32'd892
; 
32'd123866: dataIn1 = 32'd1631
; 
32'd123867: dataIn1 = 32'd1635
; 
32'd123868: dataIn1 = 32'd10367
; 
32'd123869: dataIn1 = 32'd10368
; 
32'd123870: dataIn1 = 32'd10837
; 
32'd123871: dataIn1 = 32'd10838
; 
32'd123872: dataIn1 = 32'd893
; 
32'd123873: dataIn1 = 32'd1632
; 
32'd123874: dataIn1 = 32'd1646
; 
32'd123875: dataIn1 = 32'd10371
; 
32'd123876: dataIn1 = 32'd10372
; 
32'd123877: dataIn1 = 32'd10841
; 
32'd123878: dataIn1 = 32'd10842
; 
32'd123879: dataIn1 = 32'd894
; 
32'd123880: dataIn1 = 32'd1633
; 
32'd123881: dataIn1 = 32'd1634
; 
32'd123882: dataIn1 = 32'd1933
; 
32'd123883: dataIn1 = 32'd1934
; 
32'd123884: dataIn1 = 32'd10370
; 
32'd123885: dataIn1 = 32'd10371
; 
32'd123886: dataIn1 = 32'd895
; 
32'd123887: dataIn1 = 32'd1636
; 
32'd123888: dataIn1 = 32'd1637
; 
32'd123889: dataIn1 = 32'd1935
; 
32'd123890: dataIn1 = 32'd1936
; 
32'd123891: dataIn1 = 32'd10366
; 
32'd123892: dataIn1 = 32'd10367
; 
32'd123893: dataIn1 = 32'd896
; 
32'd123894: dataIn1 = 32'd1635
; 
32'd123895: dataIn1 = 32'd1654
; 
32'd123896: dataIn1 = 32'd10365
; 
32'd123897: dataIn1 = 32'd10366
; 
32'd123898: dataIn1 = 32'd10835
; 
32'd123899: dataIn1 = 32'd10836
; 
32'd123900: dataIn1 = 32'd897
; 
32'd123901: dataIn1 = 32'd1638
; 
32'd123902: dataIn1 = 32'd1639
; 
32'd123903: dataIn1 = 32'd10375
; 
32'd123904: dataIn1 = 32'd10376
; 
32'd123905: dataIn1 = 32'd10845
; 
32'd123906: dataIn1 = 32'd10846
; 
32'd123907: dataIn1 = 32'd898
; 
32'd123908: dataIn1 = 32'd1638
; 
32'd123909: dataIn1 = 32'd1642
; 
32'd123910: dataIn1 = 32'd10377
; 
32'd123911: dataIn1 = 32'd10378
; 
32'd123912: dataIn1 = 32'd10847
; 
32'd123913: dataIn1 = 32'd10848
; 
32'd123914: dataIn1 = 32'd899
; 
32'd123915: dataIn1 = 32'd1640
; 
32'd123916: dataIn1 = 32'd1641
; 
32'd123917: dataIn1 = 32'd1937
; 
32'd123918: dataIn1 = 32'd1938
; 
32'd123919: dataIn1 = 32'd10374
; 
32'd123920: dataIn1 = 32'd10375
; 
32'd123921: dataIn1 = 32'd900
; 
32'd123922: dataIn1 = 32'd1639
; 
32'd123923: dataIn1 = 32'd1646
; 
32'd123924: dataIn1 = 32'd10373
; 
32'd123925: dataIn1 = 32'd10374
; 
32'd123926: dataIn1 = 32'd10843
; 
32'd123927: dataIn1 = 32'd10844
; 
32'd123928: dataIn1 = 32'd901
; 
32'd123929: dataIn1 = 32'd1643
; 
32'd123930: dataIn1 = 32'd1644
; 
32'd123931: dataIn1 = 32'd1939
; 
32'd123932: dataIn1 = 32'd1940
; 
32'd123933: dataIn1 = 32'd10378
; 
32'd123934: dataIn1 = 32'd10379
; 
32'd123935: dataIn1 = 32'd902
; 
32'd123936: dataIn1 = 32'd1642
; 
32'd123937: dataIn1 = 32'd1645
; 
32'd123938: dataIn1 = 32'd10379
; 
32'd123939: dataIn1 = 32'd10380
; 
32'd123940: dataIn1 = 32'd10849
; 
32'd123941: dataIn1 = 32'd10850
; 
32'd123942: dataIn1 = 32'd903
; 
32'd123943: dataIn1 = 32'd1647
; 
32'd123944: dataIn1 = 32'd1648
; 
32'd123945: dataIn1 = 32'd10359
; 
32'd123946: dataIn1 = 32'd10360
; 
32'd123947: dataIn1 = 32'd10829
; 
32'd123948: dataIn1 = 32'd10830
; 
32'd123949: dataIn1 = 32'd904
; 
32'd123950: dataIn1 = 32'd1647
; 
32'd123951: dataIn1 = 32'd1651
; 
32'd123952: dataIn1 = 32'd10361
; 
32'd123953: dataIn1 = 32'd10362
; 
32'd123954: dataIn1 = 32'd10831
; 
32'd123955: dataIn1 = 32'd10832
; 
32'd123956: dataIn1 = 32'd905
; 
32'd123957: dataIn1 = 32'd1648
; 
32'd123958: dataIn1 = 32'd1655
; 
32'd123959: dataIn1 = 32'd10357
; 
32'd123960: dataIn1 = 32'd10358
; 
32'd123961: dataIn1 = 32'd10827
; 
32'd123962: dataIn1 = 32'd10828
; 
32'd123963: dataIn1 = 32'd906
; 
32'd123964: dataIn1 = 32'd1649
; 
32'd123965: dataIn1 = 32'd1650
; 
32'd123966: dataIn1 = 32'd1941
; 
32'd123967: dataIn1 = 32'd1942
; 
32'd123968: dataIn1 = 32'd10358
; 
32'd123969: dataIn1 = 32'd10359
; 
32'd123970: dataIn1 = 32'd907
; 
32'd123971: dataIn1 = 32'd1651
; 
32'd123972: dataIn1 = 32'd1654
; 
32'd123973: dataIn1 = 32'd10363
; 
32'd123974: dataIn1 = 32'd10364
; 
32'd123975: dataIn1 = 32'd10833
; 
32'd123976: dataIn1 = 32'd10834
; 
32'd123977: dataIn1 = 32'd908
; 
32'd123978: dataIn1 = 32'd1652
; 
32'd123979: dataIn1 = 32'd1653
; 
32'd123980: dataIn1 = 32'd1943
; 
32'd123981: dataIn1 = 32'd1944
; 
32'd123982: dataIn1 = 32'd10362
; 
32'd123983: dataIn1 = 32'd10363
; 
32'd123984: dataIn1 = 32'd909
; 
32'd123985: dataIn1 = 32'd1655
; 
32'd123986: dataIn1 = 32'd1657
; 
32'd123987: dataIn1 = 32'd10355
; 
32'd123988: dataIn1 = 32'd10356
; 
32'd123989: dataIn1 = 32'd10825
; 
32'd123990: dataIn1 = 32'd10826
; 
32'd123991: dataIn1 = 32'd910
; 
32'd123992: dataIn1 = 32'd1656
; 
32'd123993: dataIn1 = 32'd1657
; 
32'd123994: dataIn1 = 32'd10353
; 
32'd123995: dataIn1 = 32'd10354
; 
32'd123996: dataIn1 = 32'd10823
; 
32'd123997: dataIn1 = 32'd10824
; 
32'd123998: dataIn1 = 32'd911
; 
32'd123999: dataIn1 = 32'd1656
; 
32'd124000: dataIn1 = 32'd1660
; 
32'd124001: dataIn1 = 32'd10351
; 
32'd124002: dataIn1 = 32'd10352
; 
32'd124003: dataIn1 = 32'd10821
; 
32'd124004: dataIn1 = 32'd10822
; 
32'd124005: dataIn1 = 32'd912
; 
32'd124006: dataIn1 = 32'd1658
; 
32'd124007: dataIn1 = 32'd1659
; 
32'd124008: dataIn1 = 32'd1945
; 
32'd124009: dataIn1 = 32'd1946
; 
32'd124010: dataIn1 = 32'd10354
; 
32'd124011: dataIn1 = 32'd10355
; 
32'd124012: dataIn1 = 32'd913
; 
32'd124013: dataIn1 = 32'd1660
; 
32'd124014: dataIn1 = 32'd1677
; 
32'd124015: dataIn1 = 32'd10349
; 
32'd124016: dataIn1 = 32'd10350
; 
32'd124017: dataIn1 = 32'd10819
; 
32'd124018: dataIn1 = 32'd10820
; 
32'd124019: dataIn1 = 32'd914
; 
32'd124020: dataIn1 = 32'd1661
; 
32'd124021: dataIn1 = 32'd1662
; 
32'd124022: dataIn1 = 32'd1947
; 
32'd124023: dataIn1 = 32'd1948
; 
32'd124024: dataIn1 = 32'd10350
; 
32'd124025: dataIn1 = 32'd10351
; 
32'd124026: dataIn1 = 32'd915
; 
32'd124027: dataIn1 = 32'd1663
; 
32'd124028: dataIn1 = 32'd1664
; 
32'd124029: dataIn1 = 32'd10337
; 
32'd124030: dataIn1 = 32'd10338
; 
32'd124031: dataIn1 = 32'd10807
; 
32'd124032: dataIn1 = 32'd10808
; 
32'd124033: dataIn1 = 32'd916
; 
32'd124034: dataIn1 = 32'd1663
; 
32'd124035: dataIn1 = 32'd1667
; 
32'd124036: dataIn1 = 32'd10335
; 
32'd124037: dataIn1 = 32'd10336
; 
32'd124038: dataIn1 = 32'd10805
; 
32'd124039: dataIn1 = 32'd10806
; 
32'd124040: dataIn1 = 32'd917
; 
32'd124041: dataIn1 = 32'd1664
; 
32'd124042: dataIn1 = 32'd1678
; 
32'd124043: dataIn1 = 32'd10339
; 
32'd124044: dataIn1 = 32'd10340
; 
32'd124045: dataIn1 = 32'd10809
; 
32'd124046: dataIn1 = 32'd10810
; 
32'd124047: dataIn1 = 32'd918
; 
32'd124048: dataIn1 = 32'd1665
; 
32'd124049: dataIn1 = 32'd1666
; 
32'd124050: dataIn1 = 32'd1949
; 
32'd124051: dataIn1 = 32'd1950
; 
32'd124052: dataIn1 = 32'd10338
; 
32'd124053: dataIn1 = 32'd10339
; 
32'd124054: dataIn1 = 32'd919
; 
32'd124055: dataIn1 = 32'd1668
; 
32'd124056: dataIn1 = 32'd1669
; 
32'd124057: dataIn1 = 32'd1951
; 
32'd124058: dataIn1 = 32'd1952
; 
32'd124059: dataIn1 = 32'd10334
; 
32'd124060: dataIn1 = 32'd10335
; 
32'd124061: dataIn1 = 32'd920
; 
32'd124062: dataIn1 = 32'd1667
; 
32'd124063: dataIn1 = 32'd1686
; 
32'd124064: dataIn1 = 32'd10333
; 
32'd124065: dataIn1 = 32'd10334
; 
32'd124066: dataIn1 = 32'd10803
; 
32'd124067: dataIn1 = 32'd10804
; 
32'd124068: dataIn1 = 32'd921
; 
32'd124069: dataIn1 = 32'd1670
; 
32'd124070: dataIn1 = 32'd1671
; 
32'd124071: dataIn1 = 32'd10343
; 
32'd124072: dataIn1 = 32'd10344
; 
32'd124073: dataIn1 = 32'd10813
; 
32'd124074: dataIn1 = 32'd10814
; 
32'd124075: dataIn1 = 32'd922
; 
32'd124076: dataIn1 = 32'd1670
; 
32'd124077: dataIn1 = 32'd1674
; 
32'd124078: dataIn1 = 32'd10345
; 
32'd124079: dataIn1 = 32'd10346
; 
32'd124080: dataIn1 = 32'd10815
; 
32'd124081: dataIn1 = 32'd10816
; 
32'd124082: dataIn1 = 32'd923
; 
32'd124083: dataIn1 = 32'd1672
; 
32'd124084: dataIn1 = 32'd1673
; 
32'd124085: dataIn1 = 32'd1953
; 
32'd124086: dataIn1 = 32'd1954
; 
32'd124087: dataIn1 = 32'd10342
; 
32'd124088: dataIn1 = 32'd10343
; 
32'd124089: dataIn1 = 32'd924
; 
32'd124090: dataIn1 = 32'd1671
; 
32'd124091: dataIn1 = 32'd1678
; 
32'd124092: dataIn1 = 32'd10341
; 
32'd124093: dataIn1 = 32'd10342
; 
32'd124094: dataIn1 = 32'd10811
; 
32'd124095: dataIn1 = 32'd10812
; 
32'd124096: dataIn1 = 32'd925
; 
32'd124097: dataIn1 = 32'd1675
; 
32'd124098: dataIn1 = 32'd1676
; 
32'd124099: dataIn1 = 32'd1955
; 
32'd124100: dataIn1 = 32'd1956
; 
32'd124101: dataIn1 = 32'd10346
; 
32'd124102: dataIn1 = 32'd10347
; 
32'd124103: dataIn1 = 32'd926
; 
32'd124104: dataIn1 = 32'd1674
; 
32'd124105: dataIn1 = 32'd1677
; 
32'd124106: dataIn1 = 32'd10347
; 
32'd124107: dataIn1 = 32'd10348
; 
32'd124108: dataIn1 = 32'd10817
; 
32'd124109: dataIn1 = 32'd10818
; 
32'd124110: dataIn1 = 32'd927
; 
32'd124111: dataIn1 = 32'd1679
; 
32'd124112: dataIn1 = 32'd1680
; 
32'd124113: dataIn1 = 32'd10327
; 
32'd124114: dataIn1 = 32'd10328
; 
32'd124115: dataIn1 = 32'd10797
; 
32'd124116: dataIn1 = 32'd10798
; 
32'd124117: dataIn1 = 32'd928
; 
32'd124118: dataIn1 = 32'd1679
; 
32'd124119: dataIn1 = 32'd1683
; 
32'd124120: dataIn1 = 32'd10329
; 
32'd124121: dataIn1 = 32'd10330
; 
32'd124122: dataIn1 = 32'd10799
; 
32'd124123: dataIn1 = 32'd10800
; 
32'd124124: dataIn1 = 32'd929
; 
32'd124125: dataIn1 = 32'd1680
; 
32'd124126: dataIn1 = 32'd1687
; 
32'd124127: dataIn1 = 32'd10325
; 
32'd124128: dataIn1 = 32'd10326
; 
32'd124129: dataIn1 = 32'd10795
; 
32'd124130: dataIn1 = 32'd10796
; 
32'd124131: dataIn1 = 32'd930
; 
32'd124132: dataIn1 = 32'd1681
; 
32'd124133: dataIn1 = 32'd1682
; 
32'd124134: dataIn1 = 32'd1957
; 
32'd124135: dataIn1 = 32'd1958
; 
32'd124136: dataIn1 = 32'd10326
; 
32'd124137: dataIn1 = 32'd10327
; 
32'd124138: dataIn1 = 32'd931
; 
32'd124139: dataIn1 = 32'd1683
; 
32'd124140: dataIn1 = 32'd1686
; 
32'd124141: dataIn1 = 32'd10331
; 
32'd124142: dataIn1 = 32'd10332
; 
32'd124143: dataIn1 = 32'd10801
; 
32'd124144: dataIn1 = 32'd10802
; 
32'd124145: dataIn1 = 32'd932
; 
32'd124146: dataIn1 = 32'd1684
; 
32'd124147: dataIn1 = 32'd1685
; 
32'd124148: dataIn1 = 32'd1959
; 
32'd124149: dataIn1 = 32'd1960
; 
32'd124150: dataIn1 = 32'd10330
; 
32'd124151: dataIn1 = 32'd10331
; 
32'd124152: dataIn1 = 32'd933
; 
32'd124153: dataIn1 = 32'd1687
; 
32'd124154: dataIn1 = 32'd1689
; 
32'd124155: dataIn1 = 32'd10323
; 
32'd124156: dataIn1 = 32'd10324
; 
32'd124157: dataIn1 = 32'd10793
; 
32'd124158: dataIn1 = 32'd10794
; 
32'd124159: dataIn1 = 32'd934
; 
32'd124160: dataIn1 = 32'd1688
; 
32'd124161: dataIn1 = 32'd1689
; 
32'd124162: dataIn1 = 32'd10321
; 
32'd124163: dataIn1 = 32'd10322
; 
32'd124164: dataIn1 = 32'd10791
; 
32'd124165: dataIn1 = 32'd10792
; 
32'd124166: dataIn1 = 32'd935
; 
32'd124167: dataIn1 = 32'd1688
; 
32'd124168: dataIn1 = 32'd1692
; 
32'd124169: dataIn1 = 32'd10319
; 
32'd124170: dataIn1 = 32'd10320
; 
32'd124171: dataIn1 = 32'd10789
; 
32'd124172: dataIn1 = 32'd10790
; 
32'd124173: dataIn1 = 32'd936
; 
32'd124174: dataIn1 = 32'd1690
; 
32'd124175: dataIn1 = 32'd1691
; 
32'd124176: dataIn1 = 32'd1961
; 
32'd124177: dataIn1 = 32'd1962
; 
32'd124178: dataIn1 = 32'd10322
; 
32'd124179: dataIn1 = 32'd10323
; 
32'd124180: dataIn1 = 32'd937
; 
32'd124181: dataIn1 = 32'd1692
; 
32'd124182: dataIn1 = 32'd1709
; 
32'd124183: dataIn1 = 32'd10317
; 
32'd124184: dataIn1 = 32'd10318
; 
32'd124185: dataIn1 = 32'd10787
; 
32'd124186: dataIn1 = 32'd10788
; 
32'd124187: dataIn1 = 32'd938
; 
32'd124188: dataIn1 = 32'd1693
; 
32'd124189: dataIn1 = 32'd1694
; 
32'd124190: dataIn1 = 32'd1963
; 
32'd124191: dataIn1 = 32'd1964
; 
32'd124192: dataIn1 = 32'd10318
; 
32'd124193: dataIn1 = 32'd10319
; 
32'd124194: dataIn1 = 32'd939
; 
32'd124195: dataIn1 = 32'd1695
; 
32'd124196: dataIn1 = 32'd1696
; 
32'd124197: dataIn1 = 32'd10305
; 
32'd124198: dataIn1 = 32'd10306
; 
32'd124199: dataIn1 = 32'd10775
; 
32'd124200: dataIn1 = 32'd10776
; 
32'd124201: dataIn1 = 32'd940
; 
32'd124202: dataIn1 = 32'd1695
; 
32'd124203: dataIn1 = 32'd1699
; 
32'd124204: dataIn1 = 32'd10303
; 
32'd124205: dataIn1 = 32'd10304
; 
32'd124206: dataIn1 = 32'd10773
; 
32'd124207: dataIn1 = 32'd10774
; 
32'd124208: dataIn1 = 32'd941
; 
32'd124209: dataIn1 = 32'd1696
; 
32'd124210: dataIn1 = 32'd1710
; 
32'd124211: dataIn1 = 32'd10308
; 
32'd124212: dataIn1 = 32'd10309
; 
32'd124213: dataIn1 = 32'd10777
; 
32'd124214: dataIn1 = 32'd10778
; 
32'd124215: dataIn1 = 32'd942
; 
32'd124216: dataIn1 = 32'd1697
; 
32'd124217: dataIn1 = 32'd1698
; 
32'd124218: dataIn1 = 32'd1966
; 
32'd124219: dataIn1 = 32'd10306
; 
32'd124220: dataIn1 = 32'd10307
; 
32'd124221: dataIn1 = 32'd943
; 
32'd124222: dataIn1 = 32'd1700
; 
32'd124223: dataIn1 = 32'd1701
; 
32'd124224: dataIn1 = 32'd1968
; 
32'd124225: dataIn1 = 32'd10302
; 
32'd124226: dataIn1 = 32'd10303
; 
32'd124227: dataIn1 = 32'd944
; 
32'd124228: dataIn1 = 32'd1699
; 
32'd124229: dataIn1 = 32'd1718
; 
32'd124230: dataIn1 = 32'd10301
; 
32'd124231: dataIn1 = 32'd10302
; 
32'd124232: dataIn1 = 32'd10771
; 
32'd124233: dataIn1 = 32'd10772
; 
32'd124234: dataIn1 = 32'd945
; 
32'd124235: dataIn1 = 32'd1702
; 
32'd124236: dataIn1 = 32'd1703
; 
32'd124237: dataIn1 = 32'd10311
; 
32'd124238: dataIn1 = 32'd10312
; 
32'd124239: dataIn1 = 32'd10313
; 
32'd124240: dataIn1 = 32'd10781
; 
32'd124241: dataIn1 = 32'd10782
; 
32'd124242: dataIn1 = 32'd946
; 
32'd124243: dataIn1 = 32'd1702
; 
32'd124244: dataIn1 = 32'd1706
; 
32'd124245: dataIn1 = 32'd10314
; 
32'd124246: dataIn1 = 32'd10315
; 
32'd124247: dataIn1 = 32'd10783
; 
32'd124248: dataIn1 = 32'd10784
; 
32'd124249: dataIn1 = 32'd947
; 
32'd124250: dataIn1 = 32'd1704
; 
32'd124251: dataIn1 = 32'd1705
; 
32'd124252: dataIn1 = 32'd1969
; 
32'd124253: dataIn1 = 32'd10310
; 
32'd124254: dataIn1 = 32'd10311
; 
32'd124255: dataIn1 = 32'd948
; 
32'd124256: dataIn1 = 32'd1703
; 
32'd124257: dataIn1 = 32'd1710
; 
32'd124258: dataIn1 = 32'd10309
; 
32'd124259: dataIn1 = 32'd10310
; 
32'd124260: dataIn1 = 32'd10779
; 
32'd124261: dataIn1 = 32'd10780
; 
32'd124262: dataIn1 = 32'd949
; 
32'd124263: dataIn1 = 32'd1707
; 
32'd124264: dataIn1 = 32'd1708
; 
32'd124265: dataIn1 = 32'd1972
; 
32'd124266: dataIn1 = 32'd10313
; 
32'd124267: dataIn1 = 32'd10314
; 
32'd124268: dataIn1 = 32'd950
; 
32'd124269: dataIn1 = 32'd1706
; 
32'd124270: dataIn1 = 32'd1709
; 
32'd124271: dataIn1 = 32'd10316
; 
32'd124272: dataIn1 = 32'd10785
; 
32'd124273: dataIn1 = 32'd10786
; 
32'd124274: dataIn1 = 32'd951
; 
32'd124275: dataIn1 = 32'd1711
; 
32'd124276: dataIn1 = 32'd1712
; 
32'd124277: dataIn1 = 32'd10295
; 
32'd124278: dataIn1 = 32'd10296
; 
32'd124279: dataIn1 = 32'd10765
; 
32'd124280: dataIn1 = 32'd10766
; 
32'd124281: dataIn1 = 32'd952
; 
32'd124282: dataIn1 = 32'd1711
; 
32'd124283: dataIn1 = 32'd1715
; 
32'd124284: dataIn1 = 32'd10297
; 
32'd124285: dataIn1 = 32'd10298
; 
32'd124286: dataIn1 = 32'd10767
; 
32'd124287: dataIn1 = 32'd10768
; 
32'd124288: dataIn1 = 32'd953
; 
32'd124289: dataIn1 = 32'd1712
; 
32'd124290: dataIn1 = 32'd1719
; 
32'd124291: dataIn1 = 32'd10294
; 
32'd124292: dataIn1 = 32'd10762
; 
32'd124293: dataIn1 = 32'd10763
; 
32'd124294: dataIn1 = 32'd10764
; 
32'd124295: dataIn1 = 32'd954
; 
32'd124296: dataIn1 = 32'd1713
; 
32'd124297: dataIn1 = 32'd1714
; 
32'd124298: dataIn1 = 32'd1974
; 
32'd124299: dataIn1 = 32'd10293
; 
32'd124300: dataIn1 = 32'd10294
; 
32'd124301: dataIn1 = 32'd10295
; 
32'd124302: dataIn1 = 32'd955
; 
32'd124303: dataIn1 = 32'd1715
; 
32'd124304: dataIn1 = 32'd1718
; 
32'd124305: dataIn1 = 32'd10299
; 
32'd124306: dataIn1 = 32'd10300
; 
32'd124307: dataIn1 = 32'd10769
; 
32'd124308: dataIn1 = 32'd10770
; 
32'd124309: dataIn1 = 32'd956
; 
32'd124310: dataIn1 = 32'd1716
; 
32'd124311: dataIn1 = 32'd1717
; 
32'd124312: dataIn1 = 32'd1975
; 
32'd124313: dataIn1 = 32'd10298
; 
32'd124314: dataIn1 = 32'd10299
; 
32'd124315: dataIn1 = 32'd957
; 
32'd124316: dataIn1 = 32'd1719
; 
32'd124317: dataIn1 = 32'd10292
; 
32'd124318: dataIn1 = 32'd10293
; 
32'd124319: dataIn1 = 32'd10562
; 
32'd124320: dataIn1 = 32'd266
; 
32'd124321: dataIn1 = 32'd958
; 
32'd124322: dataIn1 = 32'd959
; 
32'd124323: dataIn1 = 32'd10249
; 
32'd124324: dataIn1 = 32'd10250
; 
32'd124325: dataIn1 = 32'd10253
; 
32'd124326: dataIn1 = 32'd10269
; 
32'd124327: dataIn1 = 32'd1
; 
32'd124328: dataIn1 = 32'd266
; 
32'd124329: dataIn1 = 32'd550
; 
32'd124330: dataIn1 = 32'd958
; 
32'd124331: dataIn1 = 32'd959
; 
32'd124332: dataIn1 = 32'd1265
; 
32'd124333: dataIn1 = 32'd1859
; 
32'd124334: dataIn1 = 32'd2042
; 
32'd124335: dataIn1 = 32'd10253
; 
32'd124336: dataIn1 = 32'd268
; 
32'd124337: dataIn1 = 32'd270
; 
32'd124338: dataIn1 = 32'd556
; 
32'd124339: dataIn1 = 32'd558
; 
32'd124340: dataIn1 = 32'd960
; 
32'd124341: dataIn1 = 32'd3450
; 
32'd124342: dataIn1 = 32'd3463
; 
32'd124343: dataIn1 = 32'd10254
; 
32'd124344: dataIn1 = 32'd961
; 
32'd124345: dataIn1 = 32'd1035
; 
32'd124346: dataIn1 = 32'd1831
; 
32'd124347: dataIn1 = 32'd1832
; 
32'd124348: dataIn1 = 32'd2030
; 
32'd124349: dataIn1 = 32'd2031
; 
32'd124350: dataIn1 = 32'd195
; 
32'd124351: dataIn1 = 32'd962
; 
32'd124352: dataIn1 = 32'd1829
; 
32'd124353: dataIn1 = 32'd1830
; 
32'd124354: dataIn1 = 32'd2029
; 
32'd124355: dataIn1 = 32'd2030
; 
32'd124356: dataIn1 = 32'd123
; 
32'd124357: dataIn1 = 32'd963
; 
32'd124358: dataIn1 = 32'd1835
; 
32'd124359: dataIn1 = 32'd1836
; 
32'd124360: dataIn1 = 32'd2032
; 
32'd124361: dataIn1 = 32'd964
; 
32'd124362: dataIn1 = 32'd1034
; 
32'd124363: dataIn1 = 32'd1833
; 
32'd124364: dataIn1 = 32'd1834
; 
32'd124365: dataIn1 = 32'd2029
; 
32'd124366: dataIn1 = 32'd2032
; 
32'd124367: dataIn1 = 32'd122
; 
32'd124368: dataIn1 = 32'd965
; 
32'd124369: dataIn1 = 32'd1839
; 
32'd124370: dataIn1 = 32'd1840
; 
32'd124371: dataIn1 = 32'd2031
; 
32'd124372: dataIn1 = 32'd2033
; 
32'd124373: dataIn1 = 32'd122
; 
32'd124374: dataIn1 = 32'd966
; 
32'd124375: dataIn1 = 32'd1036
; 
32'd124376: dataIn1 = 32'd1837
; 
32'd124377: dataIn1 = 32'd1838
; 
32'd124378: dataIn1 = 32'd2033
; 
32'd124379: dataIn1 = 32'd2034
; 
32'd124380: dataIn1 = 32'd199
; 
32'd124381: dataIn1 = 32'd967
; 
32'd124382: dataIn1 = 32'd1037
; 
32'd124383: dataIn1 = 32'd1843
; 
32'd124384: dataIn1 = 32'd1844
; 
32'd124385: dataIn1 = 32'd2035
; 
32'd124386: dataIn1 = 32'd2036
; 
32'd124387: dataIn1 = 32'd199
; 
32'd124388: dataIn1 = 32'd968
; 
32'd124389: dataIn1 = 32'd1036
; 
32'd124390: dataIn1 = 32'd1841
; 
32'd124391: dataIn1 = 32'd1842
; 
32'd124392: dataIn1 = 32'd2034
; 
32'd124393: dataIn1 = 32'd2035
; 
32'd124394: dataIn1 = 32'd202
; 
32'd124395: dataIn1 = 32'd969
; 
32'd124396: dataIn1 = 32'd1847
; 
32'd124397: dataIn1 = 32'd1848
; 
32'd124398: dataIn1 = 32'd2038
; 
32'd124399: dataIn1 = 32'd2039
; 
32'd124400: dataIn1 = 32'd2534
; 
32'd124401: dataIn1 = 32'd3405
; 
32'd124402: dataIn1 = 32'd202
; 
32'd124403: dataIn1 = 32'd970
; 
32'd124404: dataIn1 = 32'd1038
; 
32'd124405: dataIn1 = 32'd1845
; 
32'd124406: dataIn1 = 32'd1846
; 
32'd124407: dataIn1 = 32'd2037
; 
32'd124408: dataIn1 = 32'd2038
; 
32'd124409: dataIn1 = 32'd125
; 
32'd124410: dataIn1 = 32'd971
; 
32'd124411: dataIn1 = 32'd1037
; 
32'd124412: dataIn1 = 32'd1851
; 
32'd124413: dataIn1 = 32'd1852
; 
32'd124414: dataIn1 = 32'd2036
; 
32'd124415: dataIn1 = 32'd2040
; 
32'd124416: dataIn1 = 32'd125
; 
32'd124417: dataIn1 = 32'd972
; 
32'd124418: dataIn1 = 32'd1038
; 
32'd124419: dataIn1 = 32'd1849
; 
32'd124420: dataIn1 = 32'd1850
; 
32'd124421: dataIn1 = 32'd2037
; 
32'd124422: dataIn1 = 32'd2040
; 
32'd124423: dataIn1 = 32'd973
; 
32'd124424: dataIn1 = 32'd1862
; 
32'd124425: dataIn1 = 32'd1863
; 
32'd124426: dataIn1 = 32'd2043
; 
32'd124427: dataIn1 = 32'd2045
; 
32'd124428: dataIn1 = 32'd2523
; 
32'd124429: dataIn1 = 32'd2526
; 
32'd124430: dataIn1 = 32'd974
; 
32'd124431: dataIn1 = 32'd2523
; 
32'd124432: dataIn1 = 32'd2524
; 
32'd124433: dataIn1 = 32'd2527
; 
32'd124434: dataIn1 = 32'd5716
; 
32'd124435: dataIn1 = 32'd5717
; 
32'd124436: dataIn1 = 32'd5724
; 
32'd124437: dataIn1 = 32'd975
; 
32'd124438: dataIn1 = 32'd1860
; 
32'd124439: dataIn1 = 32'd1861
; 
32'd124440: dataIn1 = 32'd2043
; 
32'd124441: dataIn1 = 32'd2044
; 
32'd124442: dataIn1 = 32'd2528
; 
32'd124443: dataIn1 = 32'd2537
; 
32'd124444: dataIn1 = 32'd270
; 
32'd124445: dataIn1 = 32'd407
; 
32'd124446: dataIn1 = 32'd782
; 
32'd124447: dataIn1 = 32'd783
; 
32'd124448: dataIn1 = 32'd976
; 
32'd124449: dataIn1 = 32'd2497
; 
32'd124450: dataIn1 = 32'd3423
; 
32'd124451: dataIn1 = 32'd3450
; 
32'd124452: dataIn1 = 32'd3459
; 
32'd124453: dataIn1 = 32'd977
; 
32'd124454: dataIn1 = 32'd1866
; 
32'd124455: dataIn1 = 32'd1867
; 
32'd124456: dataIn1 = 32'd2046
; 
32'd124457: dataIn1 = 32'd2047
; 
32'd124458: dataIn1 = 32'd2530
; 
32'd124459: dataIn1 = 32'd2540
; 
32'd124460: dataIn1 = 32'd978
; 
32'd124461: dataIn1 = 32'd1864
; 
32'd124462: dataIn1 = 32'd1865
; 
32'd124463: dataIn1 = 32'd2044
; 
32'd124464: dataIn1 = 32'd2046
; 
32'd124465: dataIn1 = 32'd2529
; 
32'd124466: dataIn1 = 32'd2536
; 
32'd124467: dataIn1 = 32'd979
; 
32'd124468: dataIn1 = 32'd1043
; 
32'd124469: dataIn1 = 32'd1870
; 
32'd124470: dataIn1 = 32'd1871
; 
32'd124471: dataIn1 = 32'd2049
; 
32'd124472: dataIn1 = 32'd2050
; 
32'd124473: dataIn1 = 32'd5511
; 
32'd124474: dataIn1 = 32'd980
; 
32'd124475: dataIn1 = 32'd2049
; 
32'd124476: dataIn1 = 32'd3038
; 
32'd124477: dataIn1 = 32'd3039
; 
32'd124478: dataIn1 = 32'd3417
; 
32'd124479: dataIn1 = 32'd5307
; 
32'd124480: dataIn1 = 32'd5428
; 
32'd124481: dataIn1 = 32'd981
; 
32'd124482: dataIn1 = 32'd3429
; 
32'd124483: dataIn1 = 32'd3454
; 
32'd124484: dataIn1 = 32'd10251
; 
32'd124485: dataIn1 = 32'd10252
; 
32'd124486: dataIn1 = 32'd10264
; 
32'd124487: dataIn1 = 32'd10265
; 
32'd124488: dataIn1 = 32'd982
; 
32'd124489: dataIn1 = 32'd1875
; 
32'd124490: dataIn1 = 32'd1876
; 
32'd124491: dataIn1 = 32'd2047
; 
32'd124492: dataIn1 = 32'd2051
; 
32'd124493: dataIn1 = 32'd2532
; 
32'd124494: dataIn1 = 32'd2541
; 
32'd124495: dataIn1 = 32'd4618
; 
32'd124496: dataIn1 = 32'd983
; 
32'd124497: dataIn1 = 32'd1873
; 
32'd124498: dataIn1 = 32'd2051
; 
32'd124499: dataIn1 = 32'd4628
; 
32'd124500: dataIn1 = 32'd4629
; 
32'd124501: dataIn1 = 32'd4634
; 
32'd124502: dataIn1 = 32'd10273
; 
32'd124503: dataIn1 = 32'd132
; 
32'd124504: dataIn1 = 32'd984
; 
32'd124505: dataIn1 = 32'd1043
; 
32'd124506: dataIn1 = 32'd1879
; 
32'd124507: dataIn1 = 32'd1880
; 
32'd124508: dataIn1 = 32'd2050
; 
32'd124509: dataIn1 = 32'd2052
; 
32'd124510: dataIn1 = 32'd132
; 
32'd124511: dataIn1 = 32'd985
; 
32'd124512: dataIn1 = 32'd1044
; 
32'd124513: dataIn1 = 32'd1877
; 
32'd124514: dataIn1 = 32'd1878
; 
32'd124515: dataIn1 = 32'd2052
; 
32'd124516: dataIn1 = 32'd2053
; 
32'd124517: dataIn1 = 32'd215
; 
32'd124518: dataIn1 = 32'd986
; 
32'd124519: dataIn1 = 32'd1045
; 
32'd124520: dataIn1 = 32'd1883
; 
32'd124521: dataIn1 = 32'd1884
; 
32'd124522: dataIn1 = 32'd2054
; 
32'd124523: dataIn1 = 32'd2055
; 
32'd124524: dataIn1 = 32'd215
; 
32'd124525: dataIn1 = 32'd987
; 
32'd124526: dataIn1 = 32'd1044
; 
32'd124527: dataIn1 = 32'd1881
; 
32'd124528: dataIn1 = 32'd1882
; 
32'd124529: dataIn1 = 32'd2053
; 
32'd124530: dataIn1 = 32'd2054
; 
32'd124531: dataIn1 = 32'd218
; 
32'd124532: dataIn1 = 32'd988
; 
32'd124533: dataIn1 = 32'd1047
; 
32'd124534: dataIn1 = 32'd1887
; 
32'd124535: dataIn1 = 32'd1888
; 
32'd124536: dataIn1 = 32'd2057
; 
32'd124537: dataIn1 = 32'd2058
; 
32'd124538: dataIn1 = 32'd218
; 
32'd124539: dataIn1 = 32'd989
; 
32'd124540: dataIn1 = 32'd1046
; 
32'd124541: dataIn1 = 32'd1885
; 
32'd124542: dataIn1 = 32'd1886
; 
32'd124543: dataIn1 = 32'd2056
; 
32'd124544: dataIn1 = 32'd2057
; 
32'd124545: dataIn1 = 32'd134
; 
32'd124546: dataIn1 = 32'd990
; 
32'd124547: dataIn1 = 32'd1045
; 
32'd124548: dataIn1 = 32'd1891
; 
32'd124549: dataIn1 = 32'd1892
; 
32'd124550: dataIn1 = 32'd2055
; 
32'd124551: dataIn1 = 32'd2059
; 
32'd124552: dataIn1 = 32'd134
; 
32'd124553: dataIn1 = 32'd991
; 
32'd124554: dataIn1 = 32'd1046
; 
32'd124555: dataIn1 = 32'd1889
; 
32'd124556: dataIn1 = 32'd1890
; 
32'd124557: dataIn1 = 32'd2056
; 
32'd124558: dataIn1 = 32'd2059
; 
32'd124559: dataIn1 = 32'd135
; 
32'd124560: dataIn1 = 32'd992
; 
32'd124561: dataIn1 = 32'd1047
; 
32'd124562: dataIn1 = 32'd1895
; 
32'd124563: dataIn1 = 32'd1896
; 
32'd124564: dataIn1 = 32'd2058
; 
32'd124565: dataIn1 = 32'd2060
; 
32'd124566: dataIn1 = 32'd135
; 
32'd124567: dataIn1 = 32'd993
; 
32'd124568: dataIn1 = 32'd1048
; 
32'd124569: dataIn1 = 32'd1893
; 
32'd124570: dataIn1 = 32'd1894
; 
32'd124571: dataIn1 = 32'd2060
; 
32'd124572: dataIn1 = 32'd2061
; 
32'd124573: dataIn1 = 32'd221
; 
32'd124574: dataIn1 = 32'd994
; 
32'd124575: dataIn1 = 32'd1049
; 
32'd124576: dataIn1 = 32'd1899
; 
32'd124577: dataIn1 = 32'd1900
; 
32'd124578: dataIn1 = 32'd2062
; 
32'd124579: dataIn1 = 32'd2063
; 
32'd124580: dataIn1 = 32'd221
; 
32'd124581: dataIn1 = 32'd995
; 
32'd124582: dataIn1 = 32'd1048
; 
32'd124583: dataIn1 = 32'd1897
; 
32'd124584: dataIn1 = 32'd1898
; 
32'd124585: dataIn1 = 32'd2061
; 
32'd124586: dataIn1 = 32'd2062
; 
32'd124587: dataIn1 = 32'd224
; 
32'd124588: dataIn1 = 32'd996
; 
32'd124589: dataIn1 = 32'd1051
; 
32'd124590: dataIn1 = 32'd1903
; 
32'd124591: dataIn1 = 32'd1904
; 
32'd124592: dataIn1 = 32'd2065
; 
32'd124593: dataIn1 = 32'd2066
; 
32'd124594: dataIn1 = 32'd224
; 
32'd124595: dataIn1 = 32'd997
; 
32'd124596: dataIn1 = 32'd1050
; 
32'd124597: dataIn1 = 32'd1901
; 
32'd124598: dataIn1 = 32'd1902
; 
32'd124599: dataIn1 = 32'd2064
; 
32'd124600: dataIn1 = 32'd2065
; 
32'd124601: dataIn1 = 32'd137
; 
32'd124602: dataIn1 = 32'd998
; 
32'd124603: dataIn1 = 32'd1049
; 
32'd124604: dataIn1 = 32'd1907
; 
32'd124605: dataIn1 = 32'd1908
; 
32'd124606: dataIn1 = 32'd2063
; 
32'd124607: dataIn1 = 32'd2067
; 
32'd124608: dataIn1 = 32'd137
; 
32'd124609: dataIn1 = 32'd999
; 
32'd124610: dataIn1 = 32'd1050
; 
32'd124611: dataIn1 = 32'd1905
; 
32'd124612: dataIn1 = 32'd1906
; 
32'd124613: dataIn1 = 32'd2064
; 
32'd124614: dataIn1 = 32'd2067
; 
32'd124615: dataIn1 = 32'd138
; 
32'd124616: dataIn1 = 32'd1000
; 
32'd124617: dataIn1 = 32'd1051
; 
32'd124618: dataIn1 = 32'd1911
; 
32'd124619: dataIn1 = 32'd1912
; 
32'd124620: dataIn1 = 32'd2066
; 
32'd124621: dataIn1 = 32'd2068
; 
32'd124622: dataIn1 = 32'd138
; 
32'd124623: dataIn1 = 32'd1001
; 
32'd124624: dataIn1 = 32'd1052
; 
32'd124625: dataIn1 = 32'd1909
; 
32'd124626: dataIn1 = 32'd1910
; 
32'd124627: dataIn1 = 32'd2068
; 
32'd124628: dataIn1 = 32'd2069
; 
32'd124629: dataIn1 = 32'd227
; 
32'd124630: dataIn1 = 32'd1002
; 
32'd124631: dataIn1 = 32'd1053
; 
32'd124632: dataIn1 = 32'd1915
; 
32'd124633: dataIn1 = 32'd1916
; 
32'd124634: dataIn1 = 32'd2070
; 
32'd124635: dataIn1 = 32'd2071
; 
32'd124636: dataIn1 = 32'd227
; 
32'd124637: dataIn1 = 32'd1003
; 
32'd124638: dataIn1 = 32'd1052
; 
32'd124639: dataIn1 = 32'd1913
; 
32'd124640: dataIn1 = 32'd1914
; 
32'd124641: dataIn1 = 32'd2069
; 
32'd124642: dataIn1 = 32'd2070
; 
32'd124643: dataIn1 = 32'd230
; 
32'd124644: dataIn1 = 32'd1004
; 
32'd124645: dataIn1 = 32'd1055
; 
32'd124646: dataIn1 = 32'd1919
; 
32'd124647: dataIn1 = 32'd1920
; 
32'd124648: dataIn1 = 32'd2073
; 
32'd124649: dataIn1 = 32'd2074
; 
32'd124650: dataIn1 = 32'd230
; 
32'd124651: dataIn1 = 32'd1005
; 
32'd124652: dataIn1 = 32'd1054
; 
32'd124653: dataIn1 = 32'd1917
; 
32'd124654: dataIn1 = 32'd1918
; 
32'd124655: dataIn1 = 32'd2072
; 
32'd124656: dataIn1 = 32'd2073
; 
32'd124657: dataIn1 = 32'd140
; 
32'd124658: dataIn1 = 32'd1006
; 
32'd124659: dataIn1 = 32'd1053
; 
32'd124660: dataIn1 = 32'd1923
; 
32'd124661: dataIn1 = 32'd1924
; 
32'd124662: dataIn1 = 32'd2071
; 
32'd124663: dataIn1 = 32'd2075
; 
32'd124664: dataIn1 = 32'd140
; 
32'd124665: dataIn1 = 32'd1007
; 
32'd124666: dataIn1 = 32'd1054
; 
32'd124667: dataIn1 = 32'd1921
; 
32'd124668: dataIn1 = 32'd1922
; 
32'd124669: dataIn1 = 32'd2072
; 
32'd124670: dataIn1 = 32'd2075
; 
32'd124671: dataIn1 = 32'd141
; 
32'd124672: dataIn1 = 32'd1008
; 
32'd124673: dataIn1 = 32'd1055
; 
32'd124674: dataIn1 = 32'd1927
; 
32'd124675: dataIn1 = 32'd1928
; 
32'd124676: dataIn1 = 32'd2074
; 
32'd124677: dataIn1 = 32'd2076
; 
32'd124678: dataIn1 = 32'd141
; 
32'd124679: dataIn1 = 32'd1009
; 
32'd124680: dataIn1 = 32'd1056
; 
32'd124681: dataIn1 = 32'd1925
; 
32'd124682: dataIn1 = 32'd1926
; 
32'd124683: dataIn1 = 32'd2076
; 
32'd124684: dataIn1 = 32'd2077
; 
32'd124685: dataIn1 = 32'd233
; 
32'd124686: dataIn1 = 32'd1010
; 
32'd124687: dataIn1 = 32'd1057
; 
32'd124688: dataIn1 = 32'd1931
; 
32'd124689: dataIn1 = 32'd1932
; 
32'd124690: dataIn1 = 32'd2078
; 
32'd124691: dataIn1 = 32'd2079
; 
32'd124692: dataIn1 = 32'd233
; 
32'd124693: dataIn1 = 32'd1011
; 
32'd124694: dataIn1 = 32'd1056
; 
32'd124695: dataIn1 = 32'd1929
; 
32'd124696: dataIn1 = 32'd1930
; 
32'd124697: dataIn1 = 32'd2077
; 
32'd124698: dataIn1 = 32'd2078
; 
32'd124699: dataIn1 = 32'd236
; 
32'd124700: dataIn1 = 32'd1012
; 
32'd124701: dataIn1 = 32'd1059
; 
32'd124702: dataIn1 = 32'd1935
; 
32'd124703: dataIn1 = 32'd1936
; 
32'd124704: dataIn1 = 32'd2081
; 
32'd124705: dataIn1 = 32'd2082
; 
32'd124706: dataIn1 = 32'd236
; 
32'd124707: dataIn1 = 32'd1013
; 
32'd124708: dataIn1 = 32'd1058
; 
32'd124709: dataIn1 = 32'd1933
; 
32'd124710: dataIn1 = 32'd1934
; 
32'd124711: dataIn1 = 32'd2080
; 
32'd124712: dataIn1 = 32'd2081
; 
32'd124713: dataIn1 = 32'd143
; 
32'd124714: dataIn1 = 32'd1014
; 
32'd124715: dataIn1 = 32'd1057
; 
32'd124716: dataIn1 = 32'd1939
; 
32'd124717: dataIn1 = 32'd1940
; 
32'd124718: dataIn1 = 32'd2079
; 
32'd124719: dataIn1 = 32'd2083
; 
32'd124720: dataIn1 = 32'd143
; 
32'd124721: dataIn1 = 32'd1015
; 
32'd124722: dataIn1 = 32'd1058
; 
32'd124723: dataIn1 = 32'd1937
; 
32'd124724: dataIn1 = 32'd1938
; 
32'd124725: dataIn1 = 32'd2080
; 
32'd124726: dataIn1 = 32'd2083
; 
32'd124727: dataIn1 = 32'd144
; 
32'd124728: dataIn1 = 32'd1016
; 
32'd124729: dataIn1 = 32'd1059
; 
32'd124730: dataIn1 = 32'd1943
; 
32'd124731: dataIn1 = 32'd1944
; 
32'd124732: dataIn1 = 32'd2082
; 
32'd124733: dataIn1 = 32'd2084
; 
32'd124734: dataIn1 = 32'd144
; 
32'd124735: dataIn1 = 32'd1017
; 
32'd124736: dataIn1 = 32'd1060
; 
32'd124737: dataIn1 = 32'd1941
; 
32'd124738: dataIn1 = 32'd1942
; 
32'd124739: dataIn1 = 32'd2084
; 
32'd124740: dataIn1 = 32'd2085
; 
32'd124741: dataIn1 = 32'd239
; 
32'd124742: dataIn1 = 32'd1018
; 
32'd124743: dataIn1 = 32'd1061
; 
32'd124744: dataIn1 = 32'd1947
; 
32'd124745: dataIn1 = 32'd1948
; 
32'd124746: dataIn1 = 32'd2086
; 
32'd124747: dataIn1 = 32'd2087
; 
32'd124748: dataIn1 = 32'd239
; 
32'd124749: dataIn1 = 32'd1019
; 
32'd124750: dataIn1 = 32'd1060
; 
32'd124751: dataIn1 = 32'd1945
; 
32'd124752: dataIn1 = 32'd1946
; 
32'd124753: dataIn1 = 32'd2085
; 
32'd124754: dataIn1 = 32'd2086
; 
32'd124755: dataIn1 = 32'd242
; 
32'd124756: dataIn1 = 32'd1020
; 
32'd124757: dataIn1 = 32'd1063
; 
32'd124758: dataIn1 = 32'd1951
; 
32'd124759: dataIn1 = 32'd1952
; 
32'd124760: dataIn1 = 32'd2089
; 
32'd124761: dataIn1 = 32'd2090
; 
32'd124762: dataIn1 = 32'd242
; 
32'd124763: dataIn1 = 32'd1021
; 
32'd124764: dataIn1 = 32'd1062
; 
32'd124765: dataIn1 = 32'd1949
; 
32'd124766: dataIn1 = 32'd1950
; 
32'd124767: dataIn1 = 32'd2088
; 
32'd124768: dataIn1 = 32'd2089
; 
32'd124769: dataIn1 = 32'd146
; 
32'd124770: dataIn1 = 32'd1022
; 
32'd124771: dataIn1 = 32'd1061
; 
32'd124772: dataIn1 = 32'd1955
; 
32'd124773: dataIn1 = 32'd1956
; 
32'd124774: dataIn1 = 32'd2087
; 
32'd124775: dataIn1 = 32'd2091
; 
32'd124776: dataIn1 = 32'd146
; 
32'd124777: dataIn1 = 32'd1023
; 
32'd124778: dataIn1 = 32'd1062
; 
32'd124779: dataIn1 = 32'd1953
; 
32'd124780: dataIn1 = 32'd1954
; 
32'd124781: dataIn1 = 32'd2088
; 
32'd124782: dataIn1 = 32'd2091
; 
32'd124783: dataIn1 = 32'd147
; 
32'd124784: dataIn1 = 32'd1024
; 
32'd124785: dataIn1 = 32'd1063
; 
32'd124786: dataIn1 = 32'd1959
; 
32'd124787: dataIn1 = 32'd1960
; 
32'd124788: dataIn1 = 32'd2090
; 
32'd124789: dataIn1 = 32'd2092
; 
32'd124790: dataIn1 = 32'd147
; 
32'd124791: dataIn1 = 32'd1025
; 
32'd124792: dataIn1 = 32'd1064
; 
32'd124793: dataIn1 = 32'd1957
; 
32'd124794: dataIn1 = 32'd1958
; 
32'd124795: dataIn1 = 32'd2092
; 
32'd124796: dataIn1 = 32'd2093
; 
32'd124797: dataIn1 = 32'd245
; 
32'd124798: dataIn1 = 32'd1026
; 
32'd124799: dataIn1 = 32'd1065
; 
32'd124800: dataIn1 = 32'd1963
; 
32'd124801: dataIn1 = 32'd1964
; 
32'd124802: dataIn1 = 32'd2094
; 
32'd124803: dataIn1 = 32'd2095
; 
32'd124804: dataIn1 = 32'd245
; 
32'd124805: dataIn1 = 32'd1027
; 
32'd124806: dataIn1 = 32'd1064
; 
32'd124807: dataIn1 = 32'd1961
; 
32'd124808: dataIn1 = 32'd1962
; 
32'd124809: dataIn1 = 32'd2093
; 
32'd124810: dataIn1 = 32'd2094
; 
32'd124811: dataIn1 = 32'd248
; 
32'd124812: dataIn1 = 32'd1028
; 
32'd124813: dataIn1 = 32'd1967
; 
32'd124814: dataIn1 = 32'd1968
; 
32'd124815: dataIn1 = 32'd2097
; 
32'd124816: dataIn1 = 32'd2098
; 
32'd124817: dataIn1 = 32'd1029
; 
32'd124818: dataIn1 = 32'd1066
; 
32'd124819: dataIn1 = 32'd1965
; 
32'd124820: dataIn1 = 32'd1966
; 
32'd124821: dataIn1 = 32'd2096
; 
32'd124822: dataIn1 = 32'd2097
; 
32'd124823: dataIn1 = 32'd149
; 
32'd124824: dataIn1 = 32'd1030
; 
32'd124825: dataIn1 = 32'd1065
; 
32'd124826: dataIn1 = 32'd1971
; 
32'd124827: dataIn1 = 32'd1972
; 
32'd124828: dataIn1 = 32'd2095
; 
32'd124829: dataIn1 = 32'd2099
; 
32'd124830: dataIn1 = 32'd149
; 
32'd124831: dataIn1 = 32'd1031
; 
32'd124832: dataIn1 = 32'd1969
; 
32'd124833: dataIn1 = 32'd1970
; 
32'd124834: dataIn1 = 32'd2096
; 
32'd124835: dataIn1 = 32'd2099
; 
32'd124836: dataIn1 = 32'd1032
; 
32'd124837: dataIn1 = 32'd1067
; 
32'd124838: dataIn1 = 32'd1975
; 
32'd124839: dataIn1 = 32'd1976
; 
32'd124840: dataIn1 = 32'd2098
; 
32'd124841: dataIn1 = 32'd2100
; 
32'd124842: dataIn1 = 32'd150
; 
32'd124843: dataIn1 = 32'd1033
; 
32'd124844: dataIn1 = 32'd1973
; 
32'd124845: dataIn1 = 32'd1974
; 
32'd124846: dataIn1 = 32'd2100
; 
32'd124847: dataIn1 = 32'd123
; 
32'd124848: dataIn1 = 32'd195
; 
32'd124849: dataIn1 = 32'd964
; 
32'd124850: dataIn1 = 32'd1034
; 
32'd124851: dataIn1 = 32'd2029
; 
32'd124852: dataIn1 = 32'd2032
; 
32'd124853: dataIn1 = 32'd3492
; 
32'd124854: dataIn1 = 32'd3496
; 
32'd124855: dataIn1 = 32'd122
; 
32'd124856: dataIn1 = 32'd195
; 
32'd124857: dataIn1 = 32'd961
; 
32'd124858: dataIn1 = 32'd1035
; 
32'd124859: dataIn1 = 32'd2030
; 
32'd124860: dataIn1 = 32'd2031
; 
32'd124861: dataIn1 = 32'd3484
; 
32'd124862: dataIn1 = 32'd3488
; 
32'd124863: dataIn1 = 32'd122
; 
32'd124864: dataIn1 = 32'd199
; 
32'd124865: dataIn1 = 32'd966
; 
32'd124866: dataIn1 = 32'd968
; 
32'd124867: dataIn1 = 32'd1036
; 
32'd124868: dataIn1 = 32'd2034
; 
32'd124869: dataIn1 = 32'd3476
; 
32'd124870: dataIn1 = 32'd3480
; 
32'd124871: dataIn1 = 32'd125
; 
32'd124872: dataIn1 = 32'd199
; 
32'd124873: dataIn1 = 32'd967
; 
32'd124874: dataIn1 = 32'd971
; 
32'd124875: dataIn1 = 32'd1037
; 
32'd124876: dataIn1 = 32'd2036
; 
32'd124877: dataIn1 = 32'd3465
; 
32'd124878: dataIn1 = 32'd3472
; 
32'd124879: dataIn1 = 32'd125
; 
32'd124880: dataIn1 = 32'd202
; 
32'd124881: dataIn1 = 32'd970
; 
32'd124882: dataIn1 = 32'd972
; 
32'd124883: dataIn1 = 32'd1038
; 
32'd124884: dataIn1 = 32'd2037
; 
32'd124885: dataIn1 = 32'd3430
; 
32'd124886: dataIn1 = 32'd3455
; 
32'd124887: dataIn1 = 32'd202
; 
32'd124888: dataIn1 = 32'd1039
; 
32'd124889: dataIn1 = 32'd2533
; 
32'd124890: dataIn1 = 32'd2534
; 
32'd124891: dataIn1 = 32'd2535
; 
32'd124892: dataIn1 = 32'd2553
; 
32'd124893: dataIn1 = 32'd4609
; 
32'd124894: dataIn1 = 32'd4642
; 
32'd124895: dataIn1 = 32'd1040
; 
32'd124896: dataIn1 = 32'd2536
; 
32'd124897: dataIn1 = 32'd2537
; 
32'd124898: dataIn1 = 32'd5924
; 
32'd124899: dataIn1 = 32'd5926
; 
32'd124900: dataIn1 = 32'd5931
; 
32'd124901: dataIn1 = 32'd5935
; 
32'd124902: dataIn1 = 32'd1041
; 
32'd124903: dataIn1 = 32'd4613
; 
32'd124904: dataIn1 = 32'd4614
; 
32'd124905: dataIn1 = 32'd4616
; 
32'd124906: dataIn1 = 32'd4622
; 
32'd124907: dataIn1 = 32'd5914
; 
32'd124908: dataIn1 = 32'd5915
; 
32'd124909: dataIn1 = 32'd1042
; 
32'd124910: dataIn1 = 32'd4626
; 
32'd124911: dataIn1 = 32'd4627
; 
32'd124912: dataIn1 = 32'd4633
; 
32'd124913: dataIn1 = 32'd4683
; 
32'd124914: dataIn1 = 32'd5429
; 
32'd124915: dataIn1 = 32'd10267
; 
32'd124916: dataIn1 = 32'd132
; 
32'd124917: dataIn1 = 32'd212
; 
32'd124918: dataIn1 = 32'd979
; 
32'd124919: dataIn1 = 32'd984
; 
32'd124920: dataIn1 = 32'd1043
; 
32'd124921: dataIn1 = 32'd2050
; 
32'd124922: dataIn1 = 32'd2565
; 
32'd124923: dataIn1 = 32'd3431
; 
32'd124924: dataIn1 = 32'd5511
; 
32'd124925: dataIn1 = 32'd132
; 
32'd124926: dataIn1 = 32'd215
; 
32'd124927: dataIn1 = 32'd985
; 
32'd124928: dataIn1 = 32'd987
; 
32'd124929: dataIn1 = 32'd1044
; 
32'd124930: dataIn1 = 32'd2053
; 
32'd124931: dataIn1 = 32'd3432
; 
32'd124932: dataIn1 = 32'd3456
; 
32'd124933: dataIn1 = 32'd134
; 
32'd124934: dataIn1 = 32'd215
; 
32'd124935: dataIn1 = 32'd986
; 
32'd124936: dataIn1 = 32'd990
; 
32'd124937: dataIn1 = 32'd1045
; 
32'd124938: dataIn1 = 32'd2055
; 
32'd124939: dataIn1 = 32'd3466
; 
32'd124940: dataIn1 = 32'd3473
; 
32'd124941: dataIn1 = 32'd134
; 
32'd124942: dataIn1 = 32'd218
; 
32'd124943: dataIn1 = 32'd989
; 
32'd124944: dataIn1 = 32'd991
; 
32'd124945: dataIn1 = 32'd1046
; 
32'd124946: dataIn1 = 32'd2056
; 
32'd124947: dataIn1 = 32'd3477
; 
32'd124948: dataIn1 = 32'd3481
; 
32'd124949: dataIn1 = 32'd135
; 
32'd124950: dataIn1 = 32'd218
; 
32'd124951: dataIn1 = 32'd988
; 
32'd124952: dataIn1 = 32'd992
; 
32'd124953: dataIn1 = 32'd1047
; 
32'd124954: dataIn1 = 32'd2058
; 
32'd124955: dataIn1 = 32'd3485
; 
32'd124956: dataIn1 = 32'd3489
; 
32'd124957: dataIn1 = 32'd135
; 
32'd124958: dataIn1 = 32'd221
; 
32'd124959: dataIn1 = 32'd993
; 
32'd124960: dataIn1 = 32'd995
; 
32'd124961: dataIn1 = 32'd1048
; 
32'd124962: dataIn1 = 32'd2061
; 
32'd124963: dataIn1 = 32'd3493
; 
32'd124964: dataIn1 = 32'd3497
; 
32'd124965: dataIn1 = 32'd137
; 
32'd124966: dataIn1 = 32'd221
; 
32'd124967: dataIn1 = 32'd994
; 
32'd124968: dataIn1 = 32'd998
; 
32'd124969: dataIn1 = 32'd1049
; 
32'd124970: dataIn1 = 32'd2063
; 
32'd124971: dataIn1 = 32'd3500
; 
32'd124972: dataIn1 = 32'd3503
; 
32'd124973: dataIn1 = 32'd137
; 
32'd124974: dataIn1 = 32'd224
; 
32'd124975: dataIn1 = 32'd997
; 
32'd124976: dataIn1 = 32'd999
; 
32'd124977: dataIn1 = 32'd1050
; 
32'd124978: dataIn1 = 32'd2064
; 
32'd124979: dataIn1 = 32'd3505
; 
32'd124980: dataIn1 = 32'd3507
; 
32'd124981: dataIn1 = 32'd138
; 
32'd124982: dataIn1 = 32'd224
; 
32'd124983: dataIn1 = 32'd996
; 
32'd124984: dataIn1 = 32'd1000
; 
32'd124985: dataIn1 = 32'd1051
; 
32'd124986: dataIn1 = 32'd2066
; 
32'd124987: dataIn1 = 32'd3509
; 
32'd124988: dataIn1 = 32'd3511
; 
32'd124989: dataIn1 = 32'd138
; 
32'd124990: dataIn1 = 32'd227
; 
32'd124991: dataIn1 = 32'd1001
; 
32'd124992: dataIn1 = 32'd1003
; 
32'd124993: dataIn1 = 32'd1052
; 
32'd124994: dataIn1 = 32'd2069
; 
32'd124995: dataIn1 = 32'd3513
; 
32'd124996: dataIn1 = 32'd3515
; 
32'd124997: dataIn1 = 32'd140
; 
32'd124998: dataIn1 = 32'd227
; 
32'd124999: dataIn1 = 32'd1002
; 
32'd125000: dataIn1 = 32'd1006
; 
32'd125001: dataIn1 = 32'd1053
; 
32'd125002: dataIn1 = 32'd2071
; 
32'd125003: dataIn1 = 32'd3517
; 
32'd125004: dataIn1 = 32'd3519
; 
32'd125005: dataIn1 = 32'd140
; 
32'd125006: dataIn1 = 32'd230
; 
32'd125007: dataIn1 = 32'd1005
; 
32'd125008: dataIn1 = 32'd1007
; 
32'd125009: dataIn1 = 32'd1054
; 
32'd125010: dataIn1 = 32'd2072
; 
32'd125011: dataIn1 = 32'd3521
; 
32'd125012: dataIn1 = 32'd3523
; 
32'd125013: dataIn1 = 32'd141
; 
32'd125014: dataIn1 = 32'd230
; 
32'd125015: dataIn1 = 32'd1004
; 
32'd125016: dataIn1 = 32'd1008
; 
32'd125017: dataIn1 = 32'd1055
; 
32'd125018: dataIn1 = 32'd2074
; 
32'd125019: dataIn1 = 32'd3525
; 
32'd125020: dataIn1 = 32'd3527
; 
32'd125021: dataIn1 = 32'd141
; 
32'd125022: dataIn1 = 32'd233
; 
32'd125023: dataIn1 = 32'd1009
; 
32'd125024: dataIn1 = 32'd1011
; 
32'd125025: dataIn1 = 32'd1056
; 
32'd125026: dataIn1 = 32'd2077
; 
32'd125027: dataIn1 = 32'd3529
; 
32'd125028: dataIn1 = 32'd3531
; 
32'd125029: dataIn1 = 32'd143
; 
32'd125030: dataIn1 = 32'd233
; 
32'd125031: dataIn1 = 32'd1010
; 
32'd125032: dataIn1 = 32'd1014
; 
32'd125033: dataIn1 = 32'd1057
; 
32'd125034: dataIn1 = 32'd2079
; 
32'd125035: dataIn1 = 32'd3533
; 
32'd125036: dataIn1 = 32'd3535
; 
32'd125037: dataIn1 = 32'd143
; 
32'd125038: dataIn1 = 32'd236
; 
32'd125039: dataIn1 = 32'd1013
; 
32'd125040: dataIn1 = 32'd1015
; 
32'd125041: dataIn1 = 32'd1058
; 
32'd125042: dataIn1 = 32'd2080
; 
32'd125043: dataIn1 = 32'd3537
; 
32'd125044: dataIn1 = 32'd3539
; 
32'd125045: dataIn1 = 32'd144
; 
32'd125046: dataIn1 = 32'd236
; 
32'd125047: dataIn1 = 32'd1012
; 
32'd125048: dataIn1 = 32'd1016
; 
32'd125049: dataIn1 = 32'd1059
; 
32'd125050: dataIn1 = 32'd2082
; 
32'd125051: dataIn1 = 32'd3541
; 
32'd125052: dataIn1 = 32'd3543
; 
32'd125053: dataIn1 = 32'd144
; 
32'd125054: dataIn1 = 32'd239
; 
32'd125055: dataIn1 = 32'd1017
; 
32'd125056: dataIn1 = 32'd1019
; 
32'd125057: dataIn1 = 32'd1060
; 
32'd125058: dataIn1 = 32'd2085
; 
32'd125059: dataIn1 = 32'd3545
; 
32'd125060: dataIn1 = 32'd3547
; 
32'd125061: dataIn1 = 32'd146
; 
32'd125062: dataIn1 = 32'd239
; 
32'd125063: dataIn1 = 32'd1018
; 
32'd125064: dataIn1 = 32'd1022
; 
32'd125065: dataIn1 = 32'd1061
; 
32'd125066: dataIn1 = 32'd2087
; 
32'd125067: dataIn1 = 32'd3549
; 
32'd125068: dataIn1 = 32'd3551
; 
32'd125069: dataIn1 = 32'd146
; 
32'd125070: dataIn1 = 32'd242
; 
32'd125071: dataIn1 = 32'd1021
; 
32'd125072: dataIn1 = 32'd1023
; 
32'd125073: dataIn1 = 32'd1062
; 
32'd125074: dataIn1 = 32'd2088
; 
32'd125075: dataIn1 = 32'd3553
; 
32'd125076: dataIn1 = 32'd3555
; 
32'd125077: dataIn1 = 32'd147
; 
32'd125078: dataIn1 = 32'd242
; 
32'd125079: dataIn1 = 32'd1020
; 
32'd125080: dataIn1 = 32'd1024
; 
32'd125081: dataIn1 = 32'd1063
; 
32'd125082: dataIn1 = 32'd2090
; 
32'd125083: dataIn1 = 32'd3557
; 
32'd125084: dataIn1 = 32'd3559
; 
32'd125085: dataIn1 = 32'd147
; 
32'd125086: dataIn1 = 32'd245
; 
32'd125087: dataIn1 = 32'd1025
; 
32'd125088: dataIn1 = 32'd1027
; 
32'd125089: dataIn1 = 32'd1064
; 
32'd125090: dataIn1 = 32'd2093
; 
32'd125091: dataIn1 = 32'd3561
; 
32'd125092: dataIn1 = 32'd3563
; 
32'd125093: dataIn1 = 32'd149
; 
32'd125094: dataIn1 = 32'd245
; 
32'd125095: dataIn1 = 32'd1026
; 
32'd125096: dataIn1 = 32'd1030
; 
32'd125097: dataIn1 = 32'd1065
; 
32'd125098: dataIn1 = 32'd2095
; 
32'd125099: dataIn1 = 32'd3565
; 
32'd125100: dataIn1 = 32'd3567
; 
32'd125101: dataIn1 = 32'd149
; 
32'd125102: dataIn1 = 32'd248
; 
32'd125103: dataIn1 = 32'd1029
; 
32'd125104: dataIn1 = 32'd1066
; 
32'd125105: dataIn1 = 32'd2096
; 
32'd125106: dataIn1 = 32'd2097
; 
32'd125107: dataIn1 = 32'd3569
; 
32'd125108: dataIn1 = 32'd3571
; 
32'd125109: dataIn1 = 32'd150
; 
32'd125110: dataIn1 = 32'd248
; 
32'd125111: dataIn1 = 32'd1032
; 
32'd125112: dataIn1 = 32'd1067
; 
32'd125113: dataIn1 = 32'd2098
; 
32'd125114: dataIn1 = 32'd2100
; 
32'd125115: dataIn1 = 32'd3573
; 
32'd125116: dataIn1 = 32'd3575
; 
32'd125117: dataIn1 = 32'd1068
; 
32'd125118: dataIn1 = 32'd2548
; 
32'd125119: dataIn1 = 32'd2549
; 
32'd125120: dataIn1 = 32'd3492
; 
32'd125121: dataIn1 = 32'd3496
; 
32'd125122: dataIn1 = 32'd4637
; 
32'd125123: dataIn1 = 32'd1069
; 
32'd125124: dataIn1 = 32'd2547
; 
32'd125125: dataIn1 = 32'd2548
; 
32'd125126: dataIn1 = 32'd2608
; 
32'd125127: dataIn1 = 32'd2609
; 
32'd125128: dataIn1 = 32'd3484
; 
32'd125129: dataIn1 = 32'd3488
; 
32'd125130: dataIn1 = 32'd4800
; 
32'd125131: dataIn1 = 32'd1070
; 
32'd125132: dataIn1 = 32'd2550
; 
32'd125133: dataIn1 = 32'd2552
; 
32'd125134: dataIn1 = 32'd2607
; 
32'd125135: dataIn1 = 32'd2609
; 
32'd125136: dataIn1 = 32'd3476
; 
32'd125137: dataIn1 = 32'd3480
; 
32'd125138: dataIn1 = 32'd4796
; 
32'd125139: dataIn1 = 32'd1071
; 
32'd125140: dataIn1 = 32'd2550
; 
32'd125141: dataIn1 = 32'd2551
; 
32'd125142: dataIn1 = 32'd2612
; 
32'd125143: dataIn1 = 32'd2613
; 
32'd125144: dataIn1 = 32'd3465
; 
32'd125145: dataIn1 = 32'd3472
; 
32'd125146: dataIn1 = 32'd4810
; 
32'd125147: dataIn1 = 32'd1072
; 
32'd125148: dataIn1 = 32'd2556
; 
32'd125149: dataIn1 = 32'd2557
; 
32'd125150: dataIn1 = 32'd2613
; 
32'd125151: dataIn1 = 32'd2614
; 
32'd125152: dataIn1 = 32'd3430
; 
32'd125153: dataIn1 = 32'd3455
; 
32'd125154: dataIn1 = 32'd4813
; 
32'd125155: dataIn1 = 32'd1073
; 
32'd125156: dataIn1 = 32'd2553
; 
32'd125157: dataIn1 = 32'd2556
; 
32'd125158: dataIn1 = 32'd4821
; 
32'd125159: dataIn1 = 32'd4822
; 
32'd125160: dataIn1 = 32'd4835
; 
32'd125161: dataIn1 = 32'd5512
; 
32'd125162: dataIn1 = 32'd1074
; 
32'd125163: dataIn1 = 32'd4652
; 
32'd125164: dataIn1 = 32'd4671
; 
32'd125165: dataIn1 = 32'd5909
; 
32'd125166: dataIn1 = 32'd5910
; 
32'd125167: dataIn1 = 32'd6697
; 
32'd125168: dataIn1 = 32'd6702
; 
32'd125169: dataIn1 = 32'd1075
; 
32'd125170: dataIn1 = 32'd4654
; 
32'd125171: dataIn1 = 32'd4655
; 
32'd125172: dataIn1 = 32'd4662
; 
32'd125173: dataIn1 = 32'd4667
; 
32'd125174: dataIn1 = 32'd4846
; 
32'd125175: dataIn1 = 32'd4847
; 
32'd125176: dataIn1 = 32'd1076
; 
32'd125177: dataIn1 = 32'd4676
; 
32'd125178: dataIn1 = 32'd4677
; 
32'd125179: dataIn1 = 32'd4842
; 
32'd125180: dataIn1 = 32'd4843
; 
32'd125181: dataIn1 = 32'd4856
; 
32'd125182: dataIn1 = 32'd10268
; 
32'd125183: dataIn1 = 32'd1077
; 
32'd125184: dataIn1 = 32'd2565
; 
32'd125185: dataIn1 = 32'd3431
; 
32'd125186: dataIn1 = 32'd4680
; 
32'd125187: dataIn1 = 32'd4681
; 
32'd125188: dataIn1 = 32'd4887
; 
32'd125189: dataIn1 = 32'd4888
; 
32'd125190: dataIn1 = 32'd1078
; 
32'd125191: dataIn1 = 32'd3432
; 
32'd125192: dataIn1 = 32'd3456
; 
32'd125193: dataIn1 = 32'd4689
; 
32'd125194: dataIn1 = 32'd4690
; 
32'd125195: dataIn1 = 32'd4889
; 
32'd125196: dataIn1 = 32'd4890
; 
32'd125197: dataIn1 = 32'd1079
; 
32'd125198: dataIn1 = 32'd3466
; 
32'd125199: dataIn1 = 32'd3473
; 
32'd125200: dataIn1 = 32'd4691
; 
32'd125201: dataIn1 = 32'd4692
; 
32'd125202: dataIn1 = 32'd4910
; 
32'd125203: dataIn1 = 32'd4911
; 
32'd125204: dataIn1 = 32'd1080
; 
32'd125205: dataIn1 = 32'd3477
; 
32'd125206: dataIn1 = 32'd3481
; 
32'd125207: dataIn1 = 32'd4696
; 
32'd125208: dataIn1 = 32'd4697
; 
32'd125209: dataIn1 = 32'd4906
; 
32'd125210: dataIn1 = 32'd4907
; 
32'd125211: dataIn1 = 32'd1081
; 
32'd125212: dataIn1 = 32'd3485
; 
32'd125213: dataIn1 = 32'd3489
; 
32'd125214: dataIn1 = 32'd4700
; 
32'd125215: dataIn1 = 32'd4701
; 
32'd125216: dataIn1 = 32'd4925
; 
32'd125217: dataIn1 = 32'd4926
; 
32'd125218: dataIn1 = 32'd1082
; 
32'd125219: dataIn1 = 32'd3493
; 
32'd125220: dataIn1 = 32'd3497
; 
32'd125221: dataIn1 = 32'd4707
; 
32'd125222: dataIn1 = 32'd4708
; 
32'd125223: dataIn1 = 32'd4927
; 
32'd125224: dataIn1 = 32'd4928
; 
32'd125225: dataIn1 = 32'd1083
; 
32'd125226: dataIn1 = 32'd3500
; 
32'd125227: dataIn1 = 32'd3503
; 
32'd125228: dataIn1 = 32'd4709
; 
32'd125229: dataIn1 = 32'd4710
; 
32'd125230: dataIn1 = 32'd4948
; 
32'd125231: dataIn1 = 32'd4949
; 
32'd125232: dataIn1 = 32'd1084
; 
32'd125233: dataIn1 = 32'd3505
; 
32'd125234: dataIn1 = 32'd3507
; 
32'd125235: dataIn1 = 32'd4714
; 
32'd125236: dataIn1 = 32'd4715
; 
32'd125237: dataIn1 = 32'd4944
; 
32'd125238: dataIn1 = 32'd4945
; 
32'd125239: dataIn1 = 32'd1085
; 
32'd125240: dataIn1 = 32'd3509
; 
32'd125241: dataIn1 = 32'd3511
; 
32'd125242: dataIn1 = 32'd4718
; 
32'd125243: dataIn1 = 32'd4719
; 
32'd125244: dataIn1 = 32'd4963
; 
32'd125245: dataIn1 = 32'd4964
; 
32'd125246: dataIn1 = 32'd1086
; 
32'd125247: dataIn1 = 32'd3513
; 
32'd125248: dataIn1 = 32'd3515
; 
32'd125249: dataIn1 = 32'd4725
; 
32'd125250: dataIn1 = 32'd4726
; 
32'd125251: dataIn1 = 32'd4965
; 
32'd125252: dataIn1 = 32'd4966
; 
32'd125253: dataIn1 = 32'd1087
; 
32'd125254: dataIn1 = 32'd3517
; 
32'd125255: dataIn1 = 32'd3519
; 
32'd125256: dataIn1 = 32'd4727
; 
32'd125257: dataIn1 = 32'd4728
; 
32'd125258: dataIn1 = 32'd4986
; 
32'd125259: dataIn1 = 32'd4987
; 
32'd125260: dataIn1 = 32'd1088
; 
32'd125261: dataIn1 = 32'd3521
; 
32'd125262: dataIn1 = 32'd3523
; 
32'd125263: dataIn1 = 32'd4732
; 
32'd125264: dataIn1 = 32'd4733
; 
32'd125265: dataIn1 = 32'd4982
; 
32'd125266: dataIn1 = 32'd4983
; 
32'd125267: dataIn1 = 32'd1089
; 
32'd125268: dataIn1 = 32'd3525
; 
32'd125269: dataIn1 = 32'd3527
; 
32'd125270: dataIn1 = 32'd4736
; 
32'd125271: dataIn1 = 32'd4737
; 
32'd125272: dataIn1 = 32'd5001
; 
32'd125273: dataIn1 = 32'd5002
; 
32'd125274: dataIn1 = 32'd1090
; 
32'd125275: dataIn1 = 32'd3529
; 
32'd125276: dataIn1 = 32'd3531
; 
32'd125277: dataIn1 = 32'd4743
; 
32'd125278: dataIn1 = 32'd4744
; 
32'd125279: dataIn1 = 32'd5003
; 
32'd125280: dataIn1 = 32'd5004
; 
32'd125281: dataIn1 = 32'd1091
; 
32'd125282: dataIn1 = 32'd3533
; 
32'd125283: dataIn1 = 32'd3535
; 
32'd125284: dataIn1 = 32'd4745
; 
32'd125285: dataIn1 = 32'd4746
; 
32'd125286: dataIn1 = 32'd5024
; 
32'd125287: dataIn1 = 32'd5025
; 
32'd125288: dataIn1 = 32'd1092
; 
32'd125289: dataIn1 = 32'd3537
; 
32'd125290: dataIn1 = 32'd3539
; 
32'd125291: dataIn1 = 32'd4750
; 
32'd125292: dataIn1 = 32'd4751
; 
32'd125293: dataIn1 = 32'd5020
; 
32'd125294: dataIn1 = 32'd5021
; 
32'd125295: dataIn1 = 32'd1093
; 
32'd125296: dataIn1 = 32'd3541
; 
32'd125297: dataIn1 = 32'd3543
; 
32'd125298: dataIn1 = 32'd4754
; 
32'd125299: dataIn1 = 32'd4755
; 
32'd125300: dataIn1 = 32'd5039
; 
32'd125301: dataIn1 = 32'd5040
; 
32'd125302: dataIn1 = 32'd1094
; 
32'd125303: dataIn1 = 32'd3545
; 
32'd125304: dataIn1 = 32'd3547
; 
32'd125305: dataIn1 = 32'd4761
; 
32'd125306: dataIn1 = 32'd4762
; 
32'd125307: dataIn1 = 32'd5041
; 
32'd125308: dataIn1 = 32'd5042
; 
32'd125309: dataIn1 = 32'd1095
; 
32'd125310: dataIn1 = 32'd3549
; 
32'd125311: dataIn1 = 32'd3551
; 
32'd125312: dataIn1 = 32'd4763
; 
32'd125313: dataIn1 = 32'd4764
; 
32'd125314: dataIn1 = 32'd5062
; 
32'd125315: dataIn1 = 32'd5063
; 
32'd125316: dataIn1 = 32'd1096
; 
32'd125317: dataIn1 = 32'd3553
; 
32'd125318: dataIn1 = 32'd3555
; 
32'd125319: dataIn1 = 32'd4768
; 
32'd125320: dataIn1 = 32'd4769
; 
32'd125321: dataIn1 = 32'd5058
; 
32'd125322: dataIn1 = 32'd5059
; 
32'd125323: dataIn1 = 32'd1097
; 
32'd125324: dataIn1 = 32'd3557
; 
32'd125325: dataIn1 = 32'd3559
; 
32'd125326: dataIn1 = 32'd4772
; 
32'd125327: dataIn1 = 32'd4773
; 
32'd125328: dataIn1 = 32'd5077
; 
32'd125329: dataIn1 = 32'd5078
; 
32'd125330: dataIn1 = 32'd1098
; 
32'd125331: dataIn1 = 32'd3561
; 
32'd125332: dataIn1 = 32'd3563
; 
32'd125333: dataIn1 = 32'd4779
; 
32'd125334: dataIn1 = 32'd4780
; 
32'd125335: dataIn1 = 32'd5079
; 
32'd125336: dataIn1 = 32'd5080
; 
32'd125337: dataIn1 = 32'd1099
; 
32'd125338: dataIn1 = 32'd3565
; 
32'd125339: dataIn1 = 32'd3567
; 
32'd125340: dataIn1 = 32'd4781
; 
32'd125341: dataIn1 = 32'd4782
; 
32'd125342: dataIn1 = 32'd5100
; 
32'd125343: dataIn1 = 32'd5101
; 
32'd125344: dataIn1 = 32'd1100
; 
32'd125345: dataIn1 = 32'd3569
; 
32'd125346: dataIn1 = 32'd3571
; 
32'd125347: dataIn1 = 32'd4786
; 
32'd125348: dataIn1 = 32'd4787
; 
32'd125349: dataIn1 = 32'd5096
; 
32'd125350: dataIn1 = 32'd5097
; 
32'd125351: dataIn1 = 32'd1101
; 
32'd125352: dataIn1 = 32'd3575
; 
32'd125353: dataIn1 = 32'd4790
; 
32'd125354: dataIn1 = 32'd4791
; 
32'd125355: dataIn1 = 32'd1102
; 
32'd125356: dataIn1 = 32'd4792
; 
32'd125357: dataIn1 = 32'd4793
; 
32'd125358: dataIn1 = 32'd9680
; 
32'd125359: dataIn1 = 32'd9681
; 
32'd125360: dataIn1 = 32'd9696
; 
32'd125361: dataIn1 = 32'd9709
; 
32'd125362: dataIn1 = 32'd1103
; 
32'd125363: dataIn1 = 32'd4805
; 
32'd125364: dataIn1 = 32'd4807
; 
32'd125365: dataIn1 = 32'd9711
; 
32'd125366: dataIn1 = 32'd9712
; 
32'd125367: dataIn1 = 32'd9719
; 
32'd125368: dataIn1 = 32'd9729
; 
32'd125369: dataIn1 = 32'd1104
; 
32'd125370: dataIn1 = 32'd4825
; 
32'd125371: dataIn1 = 32'd4826
; 
32'd125372: dataIn1 = 32'd4837
; 
32'd125373: dataIn1 = 32'd6935
; 
32'd125374: dataIn1 = 32'd6936
; 
32'd125375: dataIn1 = 32'd6971
; 
32'd125376: dataIn1 = 32'd1105
; 
32'd125377: dataIn1 = 32'd5958
; 
32'd125378: dataIn1 = 32'd5959
; 
32'd125379: dataIn1 = 32'd5977
; 
32'd125380: dataIn1 = 32'd5990
; 
32'd125381: dataIn1 = 32'd7294
; 
32'd125382: dataIn1 = 32'd7295
; 
32'd125383: dataIn1 = 32'd1106
; 
32'd125384: dataIn1 = 32'd6019
; 
32'd125385: dataIn1 = 32'd6020
; 
32'd125386: dataIn1 = 32'd6042
; 
32'd125387: dataIn1 = 32'd6060
; 
32'd125388: dataIn1 = 32'd7254
; 
32'd125389: dataIn1 = 32'd7255
; 
32'd125390: dataIn1 = 32'd1107
; 
32'd125391: dataIn1 = 32'd7447
; 
32'd125392: dataIn1 = 32'd7448
; 
32'd125393: dataIn1 = 32'd7472
; 
32'd125394: dataIn1 = 32'd7494
; 
32'd125395: dataIn1 = 32'd9611
; 
32'd125396: dataIn1 = 32'd9612
; 
32'd125397: dataIn1 = 32'd1108
; 
32'd125398: dataIn1 = 32'd7524
; 
32'd125399: dataIn1 = 32'd7525
; 
32'd125400: dataIn1 = 32'd7571
; 
32'd125401: dataIn1 = 32'd7593
; 
32'd125402: dataIn1 = 32'd9623
; 
32'd125403: dataIn1 = 32'd9625
; 
32'd125404: dataIn1 = 32'd1109
; 
32'd125405: dataIn1 = 32'd7698
; 
32'd125406: dataIn1 = 32'd7699
; 
32'd125407: dataIn1 = 32'd7725
; 
32'd125408: dataIn1 = 32'd7747
; 
32'd125409: dataIn1 = 32'd9644
; 
32'd125410: dataIn1 = 32'd9645
; 
32'd125411: dataIn1 = 32'd1110
; 
32'd125412: dataIn1 = 32'd4946
; 
32'd125413: dataIn1 = 32'd4947
; 
32'd125414: dataIn1 = 32'd7777
; 
32'd125415: dataIn1 = 32'd7778
; 
32'd125416: dataIn1 = 32'd7824
; 
32'd125417: dataIn1 = 32'd7846
; 
32'd125418: dataIn1 = 32'd1111
; 
32'd125419: dataIn1 = 32'd4967
; 
32'd125420: dataIn1 = 32'd4968
; 
32'd125421: dataIn1 = 32'd7951
; 
32'd125422: dataIn1 = 32'd7952
; 
32'd125423: dataIn1 = 32'd7978
; 
32'd125424: dataIn1 = 32'd8000
; 
32'd125425: dataIn1 = 32'd1112
; 
32'd125426: dataIn1 = 32'd4984
; 
32'd125427: dataIn1 = 32'd4985
; 
32'd125428: dataIn1 = 32'd8030
; 
32'd125429: dataIn1 = 32'd8031
; 
32'd125430: dataIn1 = 32'd8077
; 
32'd125431: dataIn1 = 32'd8099
; 
32'd125432: dataIn1 = 32'd1113
; 
32'd125433: dataIn1 = 32'd5005
; 
32'd125434: dataIn1 = 32'd5006
; 
32'd125435: dataIn1 = 32'd8204
; 
32'd125436: dataIn1 = 32'd8205
; 
32'd125437: dataIn1 = 32'd8231
; 
32'd125438: dataIn1 = 32'd8253
; 
32'd125439: dataIn1 = 32'd1114
; 
32'd125440: dataIn1 = 32'd5022
; 
32'd125441: dataIn1 = 32'd5023
; 
32'd125442: dataIn1 = 32'd8283
; 
32'd125443: dataIn1 = 32'd8284
; 
32'd125444: dataIn1 = 32'd8329
; 
32'd125445: dataIn1 = 32'd8351
; 
32'd125446: dataIn1 = 32'd1115
; 
32'd125447: dataIn1 = 32'd5043
; 
32'd125448: dataIn1 = 32'd5044
; 
32'd125449: dataIn1 = 32'd8456
; 
32'd125450: dataIn1 = 32'd8457
; 
32'd125451: dataIn1 = 32'd8483
; 
32'd125452: dataIn1 = 32'd8505
; 
32'd125453: dataIn1 = 32'd1116
; 
32'd125454: dataIn1 = 32'd5060
; 
32'd125455: dataIn1 = 32'd5061
; 
32'd125456: dataIn1 = 32'd8535
; 
32'd125457: dataIn1 = 32'd8536
; 
32'd125458: dataIn1 = 32'd8582
; 
32'd125459: dataIn1 = 32'd8604
; 
32'd125460: dataIn1 = 32'd1117
; 
32'd125461: dataIn1 = 32'd5081
; 
32'd125462: dataIn1 = 32'd5082
; 
32'd125463: dataIn1 = 32'd8709
; 
32'd125464: dataIn1 = 32'd8710
; 
32'd125465: dataIn1 = 32'd8736
; 
32'd125466: dataIn1 = 32'd8758
; 
32'd125467: dataIn1 = 32'd1118
; 
32'd125468: dataIn1 = 32'd5098
; 
32'd125469: dataIn1 = 32'd5099
; 
32'd125470: dataIn1 = 32'd8788
; 
32'd125471: dataIn1 = 32'd8789
; 
32'd125472: dataIn1 = 32'd8834
; 
32'd125473: dataIn1 = 32'd8856
; 
32'd125474: dataIn1 = 32'd1119
; 
32'd125475: dataIn1 = 32'd6079
; 
32'd125476: dataIn1 = 32'd6080
; 
32'd125477: dataIn1 = 32'd6131
; 
32'd125478: dataIn1 = 32'd6594
; 
32'd125479: dataIn1 = 32'd6705
; 
32'd125480: dataIn1 = 32'd6719
; 
32'd125481: dataIn1 = 32'd1120
; 
32'd125482: dataIn1 = 32'd6095
; 
32'd125483: dataIn1 = 32'd6096
; 
32'd125484: dataIn1 = 32'd6118
; 
32'd125485: dataIn1 = 32'd6706
; 
32'd125486: dataIn1 = 32'd6820
; 
32'd125487: dataIn1 = 32'd9262
; 
32'd125488: dataIn1 = 32'd1121
; 
32'd125489: dataIn1 = 32'd2702
; 
32'd125490: dataIn1 = 32'd2744
; 
32'd125491: dataIn1 = 32'd5134
; 
32'd125492: dataIn1 = 32'd5135
; 
32'd125493: dataIn1 = 32'd5148
; 
32'd125494: dataIn1 = 32'd5278
; 
32'd125495: dataIn1 = 32'd6177
; 
32'd125496: dataIn1 = 32'd1122
; 
32'd125497: dataIn1 = 32'd2701
; 
32'd125498: dataIn1 = 32'd2740
; 
32'd125499: dataIn1 = 32'd5138
; 
32'd125500: dataIn1 = 32'd5139
; 
32'd125501: dataIn1 = 32'd5144
; 
32'd125502: dataIn1 = 32'd5272
; 
32'd125503: dataIn1 = 32'd1123
; 
32'd125504: dataIn1 = 32'd6752
; 
32'd125505: dataIn1 = 32'd6753
; 
32'd125506: dataIn1 = 32'd9237
; 
32'd125507: dataIn1 = 32'd9239
; 
32'd125508: dataIn1 = 32'd9288
; 
32'd125509: dataIn1 = 32'd9291
; 
32'd125510: dataIn1 = 32'd1124
; 
32'd125511: dataIn1 = 32'd6750
; 
32'd125512: dataIn1 = 32'd6751
; 
32'd125513: dataIn1 = 32'd9238
; 
32'd125514: dataIn1 = 32'd9289
; 
32'd125515: dataIn1 = 32'd9322
; 
32'd125516: dataIn1 = 32'd9337
; 
32'd125517: dataIn1 = 32'd1125
; 
32'd125518: dataIn1 = 32'd6762
; 
32'd125519: dataIn1 = 32'd6763
; 
32'd125520: dataIn1 = 32'd9242
; 
32'd125521: dataIn1 = 32'd9245
; 
32'd125522: dataIn1 = 32'd9281
; 
32'd125523: dataIn1 = 32'd9294
; 
32'd125524: dataIn1 = 32'd1126
; 
32'd125525: dataIn1 = 32'd6760
; 
32'd125526: dataIn1 = 32'd6761
; 
32'd125527: dataIn1 = 32'd9243
; 
32'd125528: dataIn1 = 32'd9244
; 
32'd125529: dataIn1 = 32'd9295
; 
32'd125530: dataIn1 = 32'd9297
; 
32'd125531: dataIn1 = 32'd1127
; 
32'd125532: dataIn1 = 32'd6319
; 
32'd125533: dataIn1 = 32'd6320
; 
32'd125534: dataIn1 = 32'd6373
; 
32'd125535: dataIn1 = 32'd6659
; 
32'd125536: dataIn1 = 32'd6709
; 
32'd125537: dataIn1 = 32'd6726
; 
32'd125538: dataIn1 = 32'd1128
; 
32'd125539: dataIn1 = 32'd6336
; 
32'd125540: dataIn1 = 32'd6337
; 
32'd125541: dataIn1 = 32'd6360
; 
32'd125542: dataIn1 = 32'd6637
; 
32'd125543: dataIn1 = 32'd6710
; 
32'd125544: dataIn1 = 32'd6721
; 
32'd125545: dataIn1 = 32'd1129
; 
32'd125546: dataIn1 = 32'd6395
; 
32'd125547: dataIn1 = 32'd6396
; 
32'd125548: dataIn1 = 32'd6443
; 
32'd125549: dataIn1 = 32'd6678
; 
32'd125550: dataIn1 = 32'd9750
; 
32'd125551: dataIn1 = 32'd10138
; 
32'd125552: dataIn1 = 32'd10222
; 
32'd125553: dataIn1 = 32'd10282
; 
32'd125554: dataIn1 = 32'd1130
; 
32'd125555: dataIn1 = 32'd6715
; 
32'd125556: dataIn1 = 32'd6723
; 
32'd125557: dataIn1 = 32'd6764
; 
32'd125558: dataIn1 = 32'd6765
; 
32'd125559: dataIn1 = 32'd9233
; 
32'd125560: dataIn1 = 32'd9234
; 
32'd125561: dataIn1 = 32'd1131
; 
32'd125562: dataIn1 = 32'd6774
; 
32'd125563: dataIn1 = 32'd6775
; 
32'd125564: dataIn1 = 32'd9248
; 
32'd125565: dataIn1 = 32'd9251
; 
32'd125566: dataIn1 = 32'd9300
; 
32'd125567: dataIn1 = 32'd9303
; 
32'd125568: dataIn1 = 32'd1132
; 
32'd125569: dataIn1 = 32'd6772
; 
32'd125570: dataIn1 = 32'd6773
; 
32'd125571: dataIn1 = 32'd9249
; 
32'd125572: dataIn1 = 32'd9250
; 
32'd125573: dataIn1 = 32'd9283
; 
32'd125574: dataIn1 = 32'd9301
; 
32'd125575: dataIn1 = 32'd1133
; 
32'd125576: dataIn1 = 32'd6784
; 
32'd125577: dataIn1 = 32'd6785
; 
32'd125578: dataIn1 = 32'd9254
; 
32'd125579: dataIn1 = 32'd9257
; 
32'd125580: dataIn1 = 32'd9268
; 
32'd125581: dataIn1 = 32'd9306
; 
32'd125582: dataIn1 = 32'd1134
; 
32'd125583: dataIn1 = 32'd6782
; 
32'd125584: dataIn1 = 32'd6783
; 
32'd125585: dataIn1 = 32'd9255
; 
32'd125586: dataIn1 = 32'd9256
; 
32'd125587: dataIn1 = 32'd9307
; 
32'd125588: dataIn1 = 32'd9309
; 
32'd125589: dataIn1 = 32'd1135
; 
32'd125590: dataIn1 = 32'd2735
; 
32'd125591: dataIn1 = 32'd2736
; 
32'd125592: dataIn1 = 32'd2737
; 
32'd125593: dataIn1 = 32'd3433
; 
32'd125594: dataIn1 = 32'd3434
; 
32'd125595: dataIn1 = 32'd5513
; 
32'd125596: dataIn1 = 32'd6741
; 
32'd125597: dataIn1 = 32'd1136
; 
32'd125598: dataIn1 = 32'd2739
; 
32'd125599: dataIn1 = 32'd2740
; 
32'd125600: dataIn1 = 32'd2741
; 
32'd125601: dataIn1 = 32'd2742
; 
32'd125602: dataIn1 = 32'd3435
; 
32'd125603: dataIn1 = 32'd3436
; 
32'd125604: dataIn1 = 32'd1137
; 
32'd125605: dataIn1 = 32'd2744
; 
32'd125606: dataIn1 = 32'd2745
; 
32'd125607: dataIn1 = 32'd2746
; 
32'd125608: dataIn1 = 32'd3419
; 
32'd125609: dataIn1 = 32'd3437
; 
32'd125610: dataIn1 = 32'd5515
; 
32'd125611: dataIn1 = 32'd1138
; 
32'd125612: dataIn1 = 32'd2108
; 
32'd125613: dataIn1 = 32'd2748
; 
32'd125614: dataIn1 = 32'd5445
; 
32'd125615: dataIn1 = 32'd5446
; 
32'd125616: dataIn1 = 32'd5514
; 
32'd125617: dataIn1 = 32'd5517
; 
32'd125618: dataIn1 = 32'd9329
; 
32'd125619: dataIn1 = 32'd1139
; 
32'd125620: dataIn1 = 32'd2107
; 
32'd125621: dataIn1 = 32'd2109
; 
32'd125622: dataIn1 = 32'd5447
; 
32'd125623: dataIn1 = 32'd5448
; 
32'd125624: dataIn1 = 32'd5516
; 
32'd125625: dataIn1 = 32'd5519
; 
32'd125626: dataIn1 = 32'd9323
; 
32'd125627: dataIn1 = 32'd1140
; 
32'd125628: dataIn1 = 32'd2111
; 
32'd125629: dataIn1 = 32'd5449
; 
32'd125630: dataIn1 = 32'd5450
; 
32'd125631: dataIn1 = 32'd5518
; 
32'd125632: dataIn1 = 32'd5521
; 
32'd125633: dataIn1 = 32'd6743
; 
32'd125634: dataIn1 = 32'd9676
; 
32'd125635: dataIn1 = 32'd1141
; 
32'd125636: dataIn1 = 32'd5523
; 
32'd125637: dataIn1 = 32'd10154
; 
32'd125638: dataIn1 = 32'd10276
; 
32'd125639: dataIn1 = 32'd10277
; 
32'd125640: dataIn1 = 32'd10281
; 
32'd125641: dataIn1 = 32'd10283
; 
32'd125642: dataIn1 = 32'd1142
; 
32'd125643: dataIn1 = 32'd2117
; 
32'd125644: dataIn1 = 32'd2118
; 
32'd125645: dataIn1 = 32'd5453
; 
32'd125646: dataIn1 = 32'd5454
; 
32'd125647: dataIn1 = 32'd5522
; 
32'd125648: dataIn1 = 32'd5524
; 
32'd125649: dataIn1 = 32'd9334
; 
32'd125650: dataIn1 = 32'd504
; 
32'd125651: dataIn1 = 32'd1143
; 
32'd125652: dataIn1 = 32'd1144
; 
32'd125653: dataIn1 = 32'd1145
; 
32'd125654: dataIn1 = 32'd1146
; 
32'd125655: dataIn1 = 32'd10578
; 
32'd125656: dataIn1 = 32'd10579
; 
32'd125657: dataIn1 = 32'd504
; 
32'd125658: dataIn1 = 32'd1143
; 
32'd125659: dataIn1 = 32'd1144
; 
32'd125660: dataIn1 = 32'd1147
; 
32'd125661: dataIn1 = 32'd1148
; 
32'd125662: dataIn1 = 32'd10577
; 
32'd125663: dataIn1 = 32'd10578
; 
32'd125664: dataIn1 = 32'd251
; 
32'd125665: dataIn1 = 32'd1143
; 
32'd125666: dataIn1 = 32'd1145
; 
32'd125667: dataIn1 = 32'd1146
; 
32'd125668: dataIn1 = 32'd1151
; 
32'd125669: dataIn1 = 32'd10579
; 
32'd125670: dataIn1 = 32'd10580
; 
32'd125671: dataIn1 = 32'd251
; 
32'd125672: dataIn1 = 32'd504
; 
32'd125673: dataIn1 = 32'd1143
; 
32'd125674: dataIn1 = 32'd1145
; 
32'd125675: dataIn1 = 32'd1146
; 
32'd125676: dataIn1 = 32'd3556
; 
32'd125677: dataIn1 = 32'd3558
; 
32'd125678: dataIn1 = 32'd252
; 
32'd125679: dataIn1 = 32'd1144
; 
32'd125680: dataIn1 = 32'd1147
; 
32'd125681: dataIn1 = 32'd1148
; 
32'd125682: dataIn1 = 32'd1150
; 
32'd125683: dataIn1 = 32'd10576
; 
32'd125684: dataIn1 = 32'd10577
; 
32'd125685: dataIn1 = 32'd252
; 
32'd125686: dataIn1 = 32'd504
; 
32'd125687: dataIn1 = 32'd1144
; 
32'd125688: dataIn1 = 32'd1147
; 
32'd125689: dataIn1 = 32'd1148
; 
32'd125690: dataIn1 = 32'd3560
; 
32'd125691: dataIn1 = 32'd3562
; 
32'd125692: dataIn1 = 32'd505
; 
32'd125693: dataIn1 = 32'd506
; 
32'd125694: dataIn1 = 32'd1149
; 
32'd125695: dataIn1 = 32'd3558
; 
32'd125696: dataIn1 = 32'd3560
; 
32'd125697: dataIn1 = 32'd11687
; 
32'd125698: dataIn1 = 32'd11688
; 
32'd125699: dataIn1 = 32'd252
; 
32'd125700: dataIn1 = 32'd1147
; 
32'd125701: dataIn1 = 32'd1150
; 
32'd125702: dataIn1 = 32'd1164
; 
32'd125703: dataIn1 = 32'd1166
; 
32'd125704: dataIn1 = 32'd10575
; 
32'd125705: dataIn1 = 32'd10576
; 
32'd125706: dataIn1 = 32'd251
; 
32'd125707: dataIn1 = 32'd1145
; 
32'd125708: dataIn1 = 32'd1151
; 
32'd125709: dataIn1 = 32'd1189
; 
32'd125710: dataIn1 = 32'd1191
; 
32'd125711: dataIn1 = 32'd10580
; 
32'd125712: dataIn1 = 32'd10581
; 
32'd125713: dataIn1 = 32'd507
; 
32'd125714: dataIn1 = 32'd1152
; 
32'd125715: dataIn1 = 32'd1153
; 
32'd125716: dataIn1 = 32'd1154
; 
32'd125717: dataIn1 = 32'd1155
; 
32'd125718: dataIn1 = 32'd10570
; 
32'd125719: dataIn1 = 32'd10571
; 
32'd125720: dataIn1 = 32'd507
; 
32'd125721: dataIn1 = 32'd1152
; 
32'd125722: dataIn1 = 32'd1153
; 
32'd125723: dataIn1 = 32'd1156
; 
32'd125724: dataIn1 = 32'd1157
; 
32'd125725: dataIn1 = 32'd10569
; 
32'd125726: dataIn1 = 32'd10570
; 
32'd125727: dataIn1 = 32'd253
; 
32'd125728: dataIn1 = 32'd507
; 
32'd125729: dataIn1 = 32'd1152
; 
32'd125730: dataIn1 = 32'd1154
; 
32'd125731: dataIn1 = 32'd1155
; 
32'd125732: dataIn1 = 32'd3572
; 
32'd125733: dataIn1 = 32'd3574
; 
32'd125734: dataIn1 = 32'd253
; 
32'd125735: dataIn1 = 32'd1152
; 
32'd125736: dataIn1 = 32'd1154
; 
32'd125737: dataIn1 = 32'd1155
; 
32'd125738: dataIn1 = 32'd1159
; 
32'd125739: dataIn1 = 32'd10571
; 
32'd125740: dataIn1 = 32'd10572
; 
32'd125741: dataIn1 = 32'd254
; 
32'd125742: dataIn1 = 32'd507
; 
32'd125743: dataIn1 = 32'd1153
; 
32'd125744: dataIn1 = 32'd1156
; 
32'd125745: dataIn1 = 32'd1157
; 
32'd125746: dataIn1 = 32'd3576
; 
32'd125747: dataIn1 = 32'd3577
; 
32'd125748: dataIn1 = 32'd254
; 
32'd125749: dataIn1 = 32'd1153
; 
32'd125750: dataIn1 = 32'd1156
; 
32'd125751: dataIn1 = 32'd1157
; 
32'd125752: dataIn1 = 32'd1158
; 
32'd125753: dataIn1 = 32'd10567
; 
32'd125754: dataIn1 = 32'd10568
; 
32'd125755: dataIn1 = 32'd10569
; 
32'd125756: dataIn1 = 32'd254
; 
32'd125757: dataIn1 = 32'd1157
; 
32'd125758: dataIn1 = 32'd1158
; 
32'd125759: dataIn1 = 32'd1169
; 
32'd125760: dataIn1 = 32'd1171
; 
32'd125761: dataIn1 = 32'd10566
; 
32'd125762: dataIn1 = 32'd10567
; 
32'd125763: dataIn1 = 32'd253
; 
32'd125764: dataIn1 = 32'd1155
; 
32'd125765: dataIn1 = 32'd1159
; 
32'd125766: dataIn1 = 32'd1163
; 
32'd125767: dataIn1 = 32'd1165
; 
32'd125768: dataIn1 = 32'd10572
; 
32'd125769: dataIn1 = 32'd10573
; 
32'd125770: dataIn1 = 32'd508
; 
32'd125771: dataIn1 = 32'd509
; 
32'd125772: dataIn1 = 32'd1160
; 
32'd125773: dataIn1 = 32'd3574
; 
32'd125774: dataIn1 = 32'd3576
; 
32'd125775: dataIn1 = 32'd11679
; 
32'd125776: dataIn1 = 32'd11680
; 
32'd125777: dataIn1 = 32'd510
; 
32'd125778: dataIn1 = 32'd512
; 
32'd125779: dataIn1 = 32'd1161
; 
32'd125780: dataIn1 = 32'd3566
; 
32'd125781: dataIn1 = 32'd3568
; 
32'd125782: dataIn1 = 32'd11683
; 
32'd125783: dataIn1 = 32'd11684
; 
32'd125784: dataIn1 = 32'd505
; 
32'd125785: dataIn1 = 32'd510
; 
32'd125786: dataIn1 = 32'd1162
; 
32'd125787: dataIn1 = 32'd3562
; 
32'd125788: dataIn1 = 32'd3564
; 
32'd125789: dataIn1 = 32'd11685
; 
32'd125790: dataIn1 = 32'd11686
; 
32'd125791: dataIn1 = 32'd511
; 
32'd125792: dataIn1 = 32'd1159
; 
32'd125793: dataIn1 = 32'd1163
; 
32'd125794: dataIn1 = 32'd1164
; 
32'd125795: dataIn1 = 32'd1165
; 
32'd125796: dataIn1 = 32'd10573
; 
32'd125797: dataIn1 = 32'd10574
; 
32'd125798: dataIn1 = 32'd511
; 
32'd125799: dataIn1 = 32'd1150
; 
32'd125800: dataIn1 = 32'd1163
; 
32'd125801: dataIn1 = 32'd1164
; 
32'd125802: dataIn1 = 32'd1166
; 
32'd125803: dataIn1 = 32'd10574
; 
32'd125804: dataIn1 = 32'd10575
; 
32'd125805: dataIn1 = 32'd253
; 
32'd125806: dataIn1 = 32'd511
; 
32'd125807: dataIn1 = 32'd1159
; 
32'd125808: dataIn1 = 32'd1163
; 
32'd125809: dataIn1 = 32'd1165
; 
32'd125810: dataIn1 = 32'd3568
; 
32'd125811: dataIn1 = 32'd3570
; 
32'd125812: dataIn1 = 32'd252
; 
32'd125813: dataIn1 = 32'd511
; 
32'd125814: dataIn1 = 32'd1150
; 
32'd125815: dataIn1 = 32'd1164
; 
32'd125816: dataIn1 = 32'd1166
; 
32'd125817: dataIn1 = 32'd3564
; 
32'd125818: dataIn1 = 32'd3566
; 
32'd125819: dataIn1 = 32'd509
; 
32'd125820: dataIn1 = 32'd512
; 
32'd125821: dataIn1 = 32'd1167
; 
32'd125822: dataIn1 = 32'd3570
; 
32'd125823: dataIn1 = 32'd3572
; 
32'd125824: dataIn1 = 32'd11681
; 
32'd125825: dataIn1 = 32'd11682
; 
32'd125826: dataIn1 = 32'd514
; 
32'd125827: dataIn1 = 32'd515
; 
32'd125828: dataIn1 = 32'd1168
; 
32'd125829: dataIn1 = 32'd3579
; 
32'd125830: dataIn1 = 32'd3580
; 
32'd125831: dataIn1 = 32'd11676
; 
32'd125832: dataIn1 = 32'd11677
; 
32'd125833: dataIn1 = 32'd513
; 
32'd125834: dataIn1 = 32'd1158
; 
32'd125835: dataIn1 = 32'd1169
; 
32'd125836: dataIn1 = 32'd1170
; 
32'd125837: dataIn1 = 32'd1171
; 
32'd125838: dataIn1 = 32'd10565
; 
32'd125839: dataIn1 = 32'd10566
; 
32'd125840: dataIn1 = 32'd513
; 
32'd125841: dataIn1 = 32'd1169
; 
32'd125842: dataIn1 = 32'd1170
; 
32'd125843: dataIn1 = 32'd1172
; 
32'd125844: dataIn1 = 32'd1173
; 
32'd125845: dataIn1 = 32'd10565
; 
32'd125846: dataIn1 = 32'd11673
; 
32'd125847: dataIn1 = 32'd254
; 
32'd125848: dataIn1 = 32'd513
; 
32'd125849: dataIn1 = 32'd1158
; 
32'd125850: dataIn1 = 32'd1169
; 
32'd125851: dataIn1 = 32'd1171
; 
32'd125852: dataIn1 = 32'd3578
; 
32'd125853: dataIn1 = 32'd3579
; 
32'd125854: dataIn1 = 32'd255
; 
32'd125855: dataIn1 = 32'd1170
; 
32'd125856: dataIn1 = 32'd1172
; 
32'd125857: dataIn1 = 32'd1173
; 
32'd125858: dataIn1 = 32'd11673
; 
32'd125859: dataIn1 = 32'd255
; 
32'd125860: dataIn1 = 32'd513
; 
32'd125861: dataIn1 = 32'd1170
; 
32'd125862: dataIn1 = 32'd1172
; 
32'd125863: dataIn1 = 32'd1173
; 
32'd125864: dataIn1 = 32'd3580
; 
32'd125865: dataIn1 = 32'd3581
; 
32'd125866: dataIn1 = 32'd514
; 
32'd125867: dataIn1 = 32'd516
; 
32'd125868: dataIn1 = 32'd1174
; 
32'd125869: dataIn1 = 32'd3581
; 
32'd125870: dataIn1 = 32'd3582
; 
32'd125871: dataIn1 = 32'd11674
; 
32'd125872: dataIn1 = 32'd11675
; 
32'd125873: dataIn1 = 32'd508
; 
32'd125874: dataIn1 = 32'd515
; 
32'd125875: dataIn1 = 32'd1175
; 
32'd125876: dataIn1 = 32'd3577
; 
32'd125877: dataIn1 = 32'd3578
; 
32'd125878: dataIn1 = 32'd11677
; 
32'd125879: dataIn1 = 32'd11678
; 
32'd125880: dataIn1 = 32'd517
; 
32'd125881: dataIn1 = 32'd1176
; 
32'd125882: dataIn1 = 32'd1177
; 
32'd125883: dataIn1 = 32'd1178
; 
32'd125884: dataIn1 = 32'd1179
; 
32'd125885: dataIn1 = 32'd10584
; 
32'd125886: dataIn1 = 32'd10585
; 
32'd125887: dataIn1 = 32'd517
; 
32'd125888: dataIn1 = 32'd1176
; 
32'd125889: dataIn1 = 32'd1177
; 
32'd125890: dataIn1 = 32'd1180
; 
32'd125891: dataIn1 = 32'd1181
; 
32'd125892: dataIn1 = 32'd10585
; 
32'd125893: dataIn1 = 32'd10586
; 
32'd125894: dataIn1 = 32'd256
; 
32'd125895: dataIn1 = 32'd1176
; 
32'd125896: dataIn1 = 32'd1178
; 
32'd125897: dataIn1 = 32'd1179
; 
32'd125898: dataIn1 = 32'd1184
; 
32'd125899: dataIn1 = 32'd10583
; 
32'd125900: dataIn1 = 32'd10584
; 
32'd125901: dataIn1 = 32'd256
; 
32'd125902: dataIn1 = 32'd517
; 
32'd125903: dataIn1 = 32'd1176
; 
32'd125904: dataIn1 = 32'd1178
; 
32'd125905: dataIn1 = 32'd1179
; 
32'd125906: dataIn1 = 32'd3544
; 
32'd125907: dataIn1 = 32'd3546
; 
32'd125908: dataIn1 = 32'd257
; 
32'd125909: dataIn1 = 32'd517
; 
32'd125910: dataIn1 = 32'd1177
; 
32'd125911: dataIn1 = 32'd1180
; 
32'd125912: dataIn1 = 32'd1181
; 
32'd125913: dataIn1 = 32'd3540
; 
32'd125914: dataIn1 = 32'd3542
; 
32'd125915: dataIn1 = 32'd257
; 
32'd125916: dataIn1 = 32'd1177
; 
32'd125917: dataIn1 = 32'd1180
; 
32'd125918: dataIn1 = 32'd1181
; 
32'd125919: dataIn1 = 32'd1182
; 
32'd125920: dataIn1 = 32'd10586
; 
32'd125921: dataIn1 = 32'd10587
; 
32'd125922: dataIn1 = 32'd257
; 
32'd125923: dataIn1 = 32'd1181
; 
32'd125924: dataIn1 = 32'd1182
; 
32'd125925: dataIn1 = 32'd1194
; 
32'd125926: dataIn1 = 32'd1197
; 
32'd125927: dataIn1 = 32'd10587
; 
32'd125928: dataIn1 = 32'd10588
; 
32'd125929: dataIn1 = 32'd518
; 
32'd125930: dataIn1 = 32'd519
; 
32'd125931: dataIn1 = 32'd1183
; 
32'd125932: dataIn1 = 32'd3542
; 
32'd125933: dataIn1 = 32'd3544
; 
32'd125934: dataIn1 = 32'd11696
; 
32'd125935: dataIn1 = 32'd11697
; 
32'd125936: dataIn1 = 32'd256
; 
32'd125937: dataIn1 = 32'd1178
; 
32'd125938: dataIn1 = 32'd1184
; 
32'd125939: dataIn1 = 32'd1188
; 
32'd125940: dataIn1 = 32'd1190
; 
32'd125941: dataIn1 = 32'd10582
; 
32'd125942: dataIn1 = 32'd10583
; 
32'd125943: dataIn1 = 32'd520
; 
32'd125944: dataIn1 = 32'd521
; 
32'd125945: dataIn1 = 32'd1185
; 
32'd125946: dataIn1 = 32'd3550
; 
32'd125947: dataIn1 = 32'd3552
; 
32'd125948: dataIn1 = 32'd11691
; 
32'd125949: dataIn1 = 32'd11692
; 
32'd125950: dataIn1 = 32'd506
; 
32'd125951: dataIn1 = 32'd520
; 
32'd125952: dataIn1 = 32'd1186
; 
32'd125953: dataIn1 = 32'd3554
; 
32'd125954: dataIn1 = 32'd3556
; 
32'd125955: dataIn1 = 32'd11689
; 
32'd125956: dataIn1 = 32'd11690
; 
32'd125957: dataIn1 = 32'd519
; 
32'd125958: dataIn1 = 32'd521
; 
32'd125959: dataIn1 = 32'd1187
; 
32'd125960: dataIn1 = 32'd3546
; 
32'd125961: dataIn1 = 32'd3548
; 
32'd125962: dataIn1 = 32'd11693
; 
32'd125963: dataIn1 = 32'd11694
; 
32'd125964: dataIn1 = 32'd522
; 
32'd125965: dataIn1 = 32'd1184
; 
32'd125966: dataIn1 = 32'd1188
; 
32'd125967: dataIn1 = 32'd1189
; 
32'd125968: dataIn1 = 32'd1190
; 
32'd125969: dataIn1 = 32'd10581
; 
32'd125970: dataIn1 = 32'd10582
; 
32'd125971: dataIn1 = 32'd522
; 
32'd125972: dataIn1 = 32'd1151
; 
32'd125973: dataIn1 = 32'd1188
; 
32'd125974: dataIn1 = 32'd1189
; 
32'd125975: dataIn1 = 32'd1191
; 
32'd125976: dataIn1 = 32'd10581
; 
32'd125977: dataIn1 = 32'd256
; 
32'd125978: dataIn1 = 32'd522
; 
32'd125979: dataIn1 = 32'd1184
; 
32'd125980: dataIn1 = 32'd1188
; 
32'd125981: dataIn1 = 32'd1190
; 
32'd125982: dataIn1 = 32'd3548
; 
32'd125983: dataIn1 = 32'd3550
; 
32'd125984: dataIn1 = 32'd251
; 
32'd125985: dataIn1 = 32'd522
; 
32'd125986: dataIn1 = 32'd1151
; 
32'd125987: dataIn1 = 32'd1189
; 
32'd125988: dataIn1 = 32'd1191
; 
32'd125989: dataIn1 = 32'd3552
; 
32'd125990: dataIn1 = 32'd3554
; 
32'd125991: dataIn1 = 32'd524
; 
32'd125992: dataIn1 = 32'd525
; 
32'd125993: dataIn1 = 32'd1192
; 
32'd125994: dataIn1 = 32'd3534
; 
32'd125995: dataIn1 = 32'd3536
; 
32'd125996: dataIn1 = 32'd11700
; 
32'd125997: dataIn1 = 32'd11701
; 
32'd125998: dataIn1 = 32'd523
; 
32'd125999: dataIn1 = 32'd1193
; 
32'd126000: dataIn1 = 32'd1194
; 
32'd126001: dataIn1 = 32'd1195
; 
32'd126002: dataIn1 = 32'd1196
; 
32'd126003: dataIn1 = 32'd10589
; 
32'd126004: dataIn1 = 32'd10590
; 
32'd126005: dataIn1 = 32'd523
; 
32'd126006: dataIn1 = 32'd1182
; 
32'd126007: dataIn1 = 32'd1193
; 
32'd126008: dataIn1 = 32'd1194
; 
32'd126009: dataIn1 = 32'd1197
; 
32'd126010: dataIn1 = 32'd10588
; 
32'd126011: dataIn1 = 32'd10589
; 
32'd126012: dataIn1 = 32'd258
; 
32'd126013: dataIn1 = 32'd1193
; 
32'd126014: dataIn1 = 32'd1195
; 
32'd126015: dataIn1 = 32'd1196
; 
32'd126016: dataIn1 = 32'd1205
; 
32'd126017: dataIn1 = 32'd10590
; 
32'd126018: dataIn1 = 32'd10591
; 
32'd126019: dataIn1 = 32'd258
; 
32'd126020: dataIn1 = 32'd523
; 
32'd126021: dataIn1 = 32'd1193
; 
32'd126022: dataIn1 = 32'd1195
; 
32'd126023: dataIn1 = 32'd1196
; 
32'd126024: dataIn1 = 32'd3532
; 
32'd126025: dataIn1 = 32'd3534
; 
32'd126026: dataIn1 = 32'd257
; 
32'd126027: dataIn1 = 32'd523
; 
32'd126028: dataIn1 = 32'd1182
; 
32'd126029: dataIn1 = 32'd1194
; 
32'd126030: dataIn1 = 32'd1197
; 
32'd126031: dataIn1 = 32'd3536
; 
32'd126032: dataIn1 = 32'd3538
; 
32'd126033: dataIn1 = 32'd518
; 
32'd126034: dataIn1 = 32'd524
; 
32'd126035: dataIn1 = 32'd1198
; 
32'd126036: dataIn1 = 32'd3538
; 
32'd126037: dataIn1 = 32'd3540
; 
32'd126038: dataIn1 = 32'd11698
; 
32'd126039: dataIn1 = 32'd11699
; 
32'd126040: dataIn1 = 32'd525
; 
32'd126041: dataIn1 = 32'd526
; 
32'd126042: dataIn1 = 32'd1199
; 
32'd126043: dataIn1 = 32'd3530
; 
32'd126044: dataIn1 = 32'd3532
; 
32'd126045: dataIn1 = 32'd11702
; 
32'd126046: dataIn1 = 32'd11703
; 
32'd126047: dataIn1 = 32'd527
; 
32'd126048: dataIn1 = 32'd1200
; 
32'd126049: dataIn1 = 32'd1201
; 
32'd126050: dataIn1 = 32'd1202
; 
32'd126051: dataIn1 = 32'd1203
; 
32'd126052: dataIn1 = 32'd10595
; 
32'd126053: dataIn1 = 32'd10596
; 
32'd126054: dataIn1 = 32'd10597
; 
32'd126055: dataIn1 = 32'd527
; 
32'd126056: dataIn1 = 32'd1200
; 
32'd126057: dataIn1 = 32'd1201
; 
32'd126058: dataIn1 = 32'd1204
; 
32'd126059: dataIn1 = 32'd1205
; 
32'd126060: dataIn1 = 32'd10593
; 
32'd126061: dataIn1 = 32'd10594
; 
32'd126062: dataIn1 = 32'd10595
; 
32'd126063: dataIn1 = 32'd259
; 
32'd126064: dataIn1 = 32'd1200
; 
32'd126065: dataIn1 = 32'd1202
; 
32'd126066: dataIn1 = 32'd1203
; 
32'd126067: dataIn1 = 32'd1207
; 
32'd126068: dataIn1 = 32'd10597
; 
32'd126069: dataIn1 = 32'd10598
; 
32'd126070: dataIn1 = 32'd10599
; 
32'd126071: dataIn1 = 32'd259
; 
32'd126072: dataIn1 = 32'd527
; 
32'd126073: dataIn1 = 32'd1200
; 
32'd126074: dataIn1 = 32'd1202
; 
32'd126075: dataIn1 = 32'd1203
; 
32'd126076: dataIn1 = 32'd3524
; 
32'd126077: dataIn1 = 32'd3526
; 
32'd126078: dataIn1 = 32'd258
; 
32'd126079: dataIn1 = 32'd527
; 
32'd126080: dataIn1 = 32'd1201
; 
32'd126081: dataIn1 = 32'd1204
; 
32'd126082: dataIn1 = 32'd1205
; 
32'd126083: dataIn1 = 32'd3528
; 
32'd126084: dataIn1 = 32'd3530
; 
32'd126085: dataIn1 = 32'd258
; 
32'd126086: dataIn1 = 32'd1195
; 
32'd126087: dataIn1 = 32'd1201
; 
32'd126088: dataIn1 = 32'd1204
; 
32'd126089: dataIn1 = 32'd1205
; 
32'd126090: dataIn1 = 32'd10591
; 
32'd126091: dataIn1 = 32'd10592
; 
32'd126092: dataIn1 = 32'd10593
; 
32'd126093: dataIn1 = 32'd526
; 
32'd126094: dataIn1 = 32'd528
; 
32'd126095: dataIn1 = 32'd1206
; 
32'd126096: dataIn1 = 32'd3526
; 
32'd126097: dataIn1 = 32'd3528
; 
32'd126098: dataIn1 = 32'd11704
; 
32'd126099: dataIn1 = 32'd11705
; 
32'd126100: dataIn1 = 32'd259
; 
32'd126101: dataIn1 = 32'd1202
; 
32'd126102: dataIn1 = 32'd1207
; 
32'd126103: dataIn1 = 32'd1235
; 
32'd126104: dataIn1 = 32'd1237
; 
32'd126105: dataIn1 = 32'd10599
; 
32'd126106: dataIn1 = 32'd10600
; 
32'd126107: dataIn1 = 32'd10601
; 
32'd126108: dataIn1 = 32'd529
; 
32'd126109: dataIn1 = 32'd1208
; 
32'd126110: dataIn1 = 32'd1209
; 
32'd126111: dataIn1 = 32'd1210
; 
32'd126112: dataIn1 = 32'd1211
; 
32'd126113: dataIn1 = 32'd10627
; 
32'd126114: dataIn1 = 32'd10628
; 
32'd126115: dataIn1 = 32'd10629
; 
32'd126116: dataIn1 = 32'd529
; 
32'd126117: dataIn1 = 32'd1208
; 
32'd126118: dataIn1 = 32'd1209
; 
32'd126119: dataIn1 = 32'd1212
; 
32'd126120: dataIn1 = 32'd1213
; 
32'd126121: dataIn1 = 32'd10625
; 
32'd126122: dataIn1 = 32'd10626
; 
32'd126123: dataIn1 = 32'd10627
; 
32'd126124: dataIn1 = 32'd260
; 
32'd126125: dataIn1 = 32'd1208
; 
32'd126126: dataIn1 = 32'd1210
; 
32'd126127: dataIn1 = 32'd1211
; 
32'd126128: dataIn1 = 32'd1216
; 
32'd126129: dataIn1 = 32'd10629
; 
32'd126130: dataIn1 = 32'd10630
; 
32'd126131: dataIn1 = 32'd10631
; 
32'd126132: dataIn1 = 32'd260
; 
32'd126133: dataIn1 = 32'd529
; 
32'd126134: dataIn1 = 32'd1208
; 
32'd126135: dataIn1 = 32'd1210
; 
32'd126136: dataIn1 = 32'd1211
; 
32'd126137: dataIn1 = 32'd3482
; 
32'd126138: dataIn1 = 32'd3486
; 
32'd126139: dataIn1 = 32'd261
; 
32'd126140: dataIn1 = 32'd1209
; 
32'd126141: dataIn1 = 32'd1212
; 
32'd126142: dataIn1 = 32'd1213
; 
32'd126143: dataIn1 = 32'd1215
; 
32'd126144: dataIn1 = 32'd10623
; 
32'd126145: dataIn1 = 32'd10624
; 
32'd126146: dataIn1 = 32'd10625
; 
32'd126147: dataIn1 = 32'd261
; 
32'd126148: dataIn1 = 32'd529
; 
32'd126149: dataIn1 = 32'd1209
; 
32'd126150: dataIn1 = 32'd1212
; 
32'd126151: dataIn1 = 32'd1213
; 
32'd126152: dataIn1 = 32'd3490
; 
32'd126153: dataIn1 = 32'd3494
; 
32'd126154: dataIn1 = 32'd530
; 
32'd126155: dataIn1 = 32'd531
; 
32'd126156: dataIn1 = 32'd1214
; 
32'd126157: dataIn1 = 32'd3486
; 
32'd126158: dataIn1 = 32'd3490
; 
32'd126159: dataIn1 = 32'd11720
; 
32'd126160: dataIn1 = 32'd11721
; 
32'd126161: dataIn1 = 32'd261
; 
32'd126162: dataIn1 = 32'd1212
; 
32'd126163: dataIn1 = 32'd1215
; 
32'd126164: dataIn1 = 32'd1229
; 
32'd126165: dataIn1 = 32'd1231
; 
32'd126166: dataIn1 = 32'd10621
; 
32'd126167: dataIn1 = 32'd10622
; 
32'd126168: dataIn1 = 32'd10623
; 
32'd126169: dataIn1 = 32'd260
; 
32'd126170: dataIn1 = 32'd1210
; 
32'd126171: dataIn1 = 32'd1216
; 
32'd126172: dataIn1 = 32'd1255
; 
32'd126173: dataIn1 = 32'd1257
; 
32'd126174: dataIn1 = 32'd10631
; 
32'd126175: dataIn1 = 32'd10632
; 
32'd126176: dataIn1 = 32'd10633
; 
32'd126177: dataIn1 = 32'd532
; 
32'd126178: dataIn1 = 32'd1217
; 
32'd126179: dataIn1 = 32'd1218
; 
32'd126180: dataIn1 = 32'd1219
; 
32'd126181: dataIn1 = 32'd1220
; 
32'd126182: dataIn1 = 32'd10612
; 
32'd126183: dataIn1 = 32'd10613
; 
32'd126184: dataIn1 = 32'd10614
; 
32'd126185: dataIn1 = 32'd532
; 
32'd126186: dataIn1 = 32'd1217
; 
32'd126187: dataIn1 = 32'd1218
; 
32'd126188: dataIn1 = 32'd1221
; 
32'd126189: dataIn1 = 32'd1222
; 
32'd126190: dataIn1 = 32'd10610
; 
32'd126191: dataIn1 = 32'd10611
; 
32'd126192: dataIn1 = 32'd10612
; 
32'd126193: dataIn1 = 32'd262
; 
32'd126194: dataIn1 = 32'd532
; 
32'd126195: dataIn1 = 32'd1217
; 
32'd126196: dataIn1 = 32'd1219
; 
32'd126197: dataIn1 = 32'd1220
; 
32'd126198: dataIn1 = 32'd3508
; 
32'd126199: dataIn1 = 32'd3510
; 
32'd126200: dataIn1 = 32'd262
; 
32'd126201: dataIn1 = 32'd1217
; 
32'd126202: dataIn1 = 32'd1219
; 
32'd126203: dataIn1 = 32'd1220
; 
32'd126204: dataIn1 = 32'd1224
; 
32'd126205: dataIn1 = 32'd10614
; 
32'd126206: dataIn1 = 32'd10615
; 
32'd126207: dataIn1 = 32'd10616
; 
32'd126208: dataIn1 = 32'd263
; 
32'd126209: dataIn1 = 32'd532
; 
32'd126210: dataIn1 = 32'd1218
; 
32'd126211: dataIn1 = 32'd1221
; 
32'd126212: dataIn1 = 32'd1222
; 
32'd126213: dataIn1 = 32'd3512
; 
32'd126214: dataIn1 = 32'd3514
; 
32'd126215: dataIn1 = 32'd263
; 
32'd126216: dataIn1 = 32'd1218
; 
32'd126217: dataIn1 = 32'd1221
; 
32'd126218: dataIn1 = 32'd1222
; 
32'd126219: dataIn1 = 32'd1223
; 
32'd126220: dataIn1 = 32'd10607
; 
32'd126221: dataIn1 = 32'd10608
; 
32'd126222: dataIn1 = 32'd10609
; 
32'd126223: dataIn1 = 32'd10610
; 
32'd126224: dataIn1 = 32'd263
; 
32'd126225: dataIn1 = 32'd1222
; 
32'd126226: dataIn1 = 32'd1223
; 
32'd126227: dataIn1 = 32'd1234
; 
32'd126228: dataIn1 = 32'd1236
; 
32'd126229: dataIn1 = 32'd10605
; 
32'd126230: dataIn1 = 32'd10606
; 
32'd126231: dataIn1 = 32'd10607
; 
32'd126232: dataIn1 = 32'd262
; 
32'd126233: dataIn1 = 32'd1220
; 
32'd126234: dataIn1 = 32'd1224
; 
32'd126235: dataIn1 = 32'd1228
; 
32'd126236: dataIn1 = 32'd1230
; 
32'd126237: dataIn1 = 32'd10616
; 
32'd126238: dataIn1 = 32'd10617
; 
32'd126239: dataIn1 = 32'd10618
; 
32'd126240: dataIn1 = 32'd533
; 
32'd126241: dataIn1 = 32'd534
; 
32'd126242: dataIn1 = 32'd1225
; 
32'd126243: dataIn1 = 32'd3510
; 
32'd126244: dataIn1 = 32'd3512
; 
32'd126245: dataIn1 = 32'd11712
; 
32'd126246: dataIn1 = 32'd11713
; 
32'd126247: dataIn1 = 32'd535
; 
32'd126248: dataIn1 = 32'd537
; 
32'd126249: dataIn1 = 32'd1226
; 
32'd126250: dataIn1 = 32'd3501
; 
32'd126251: dataIn1 = 32'd3504
; 
32'd126252: dataIn1 = 32'd11716
; 
32'd126253: dataIn1 = 32'd11717
; 
32'd126254: dataIn1 = 32'd530
; 
32'd126255: dataIn1 = 32'd535
; 
32'd126256: dataIn1 = 32'd1227
; 
32'd126257: dataIn1 = 32'd3494
; 
32'd126258: dataIn1 = 32'd3498
; 
32'd126259: dataIn1 = 32'd11718
; 
32'd126260: dataIn1 = 32'd11719
; 
32'd126261: dataIn1 = 32'd536
; 
32'd126262: dataIn1 = 32'd1224
; 
32'd126263: dataIn1 = 32'd1228
; 
32'd126264: dataIn1 = 32'd1229
; 
32'd126265: dataIn1 = 32'd1230
; 
32'd126266: dataIn1 = 32'd10618
; 
32'd126267: dataIn1 = 32'd10619
; 
32'd126268: dataIn1 = 32'd10620
; 
32'd126269: dataIn1 = 32'd536
; 
32'd126270: dataIn1 = 32'd1215
; 
32'd126271: dataIn1 = 32'd1228
; 
32'd126272: dataIn1 = 32'd1229
; 
32'd126273: dataIn1 = 32'd1231
; 
32'd126274: dataIn1 = 32'd10620
; 
32'd126275: dataIn1 = 32'd10621
; 
32'd126276: dataIn1 = 32'd262
; 
32'd126277: dataIn1 = 32'd536
; 
32'd126278: dataIn1 = 32'd1224
; 
32'd126279: dataIn1 = 32'd1228
; 
32'd126280: dataIn1 = 32'd1230
; 
32'd126281: dataIn1 = 32'd3504
; 
32'd126282: dataIn1 = 32'd3506
; 
32'd126283: dataIn1 = 32'd261
; 
32'd126284: dataIn1 = 32'd536
; 
32'd126285: dataIn1 = 32'd1215
; 
32'd126286: dataIn1 = 32'd1229
; 
32'd126287: dataIn1 = 32'd1231
; 
32'd126288: dataIn1 = 32'd3498
; 
32'd126289: dataIn1 = 32'd3501
; 
32'd126290: dataIn1 = 32'd534
; 
32'd126291: dataIn1 = 32'd537
; 
32'd126292: dataIn1 = 32'd1232
; 
32'd126293: dataIn1 = 32'd3506
; 
32'd126294: dataIn1 = 32'd3508
; 
32'd126295: dataIn1 = 32'd11714
; 
32'd126296: dataIn1 = 32'd11715
; 
32'd126297: dataIn1 = 32'd539
; 
32'd126298: dataIn1 = 32'd540
; 
32'd126299: dataIn1 = 32'd1233
; 
32'd126300: dataIn1 = 32'd3518
; 
32'd126301: dataIn1 = 32'd3520
; 
32'd126302: dataIn1 = 32'd11708
; 
32'd126303: dataIn1 = 32'd11709
; 
32'd126304: dataIn1 = 32'd538
; 
32'd126305: dataIn1 = 32'd1223
; 
32'd126306: dataIn1 = 32'd1234
; 
32'd126307: dataIn1 = 32'd1235
; 
32'd126308: dataIn1 = 32'd1236
; 
32'd126309: dataIn1 = 32'd10603
; 
32'd126310: dataIn1 = 32'd10604
; 
32'd126311: dataIn1 = 32'd10605
; 
32'd126312: dataIn1 = 32'd538
; 
32'd126313: dataIn1 = 32'd1207
; 
32'd126314: dataIn1 = 32'd1234
; 
32'd126315: dataIn1 = 32'd1235
; 
32'd126316: dataIn1 = 32'd1237
; 
32'd126317: dataIn1 = 32'd10601
; 
32'd126318: dataIn1 = 32'd10602
; 
32'd126319: dataIn1 = 32'd10603
; 
32'd126320: dataIn1 = 32'd263
; 
32'd126321: dataIn1 = 32'd538
; 
32'd126322: dataIn1 = 32'd1223
; 
32'd126323: dataIn1 = 32'd1234
; 
32'd126324: dataIn1 = 32'd1236
; 
32'd126325: dataIn1 = 32'd3516
; 
32'd126326: dataIn1 = 32'd3518
; 
32'd126327: dataIn1 = 32'd259
; 
32'd126328: dataIn1 = 32'd538
; 
32'd126329: dataIn1 = 32'd1207
; 
32'd126330: dataIn1 = 32'd1235
; 
32'd126331: dataIn1 = 32'd1237
; 
32'd126332: dataIn1 = 32'd3520
; 
32'd126333: dataIn1 = 32'd3522
; 
32'd126334: dataIn1 = 32'd528
; 
32'd126335: dataIn1 = 32'd539
; 
32'd126336: dataIn1 = 32'd1238
; 
32'd126337: dataIn1 = 32'd3522
; 
32'd126338: dataIn1 = 32'd3524
; 
32'd126339: dataIn1 = 32'd11706
; 
32'd126340: dataIn1 = 32'd11707
; 
32'd126341: dataIn1 = 32'd533
; 
32'd126342: dataIn1 = 32'd540
; 
32'd126343: dataIn1 = 32'd1239
; 
32'd126344: dataIn1 = 32'd3514
; 
32'd126345: dataIn1 = 32'd3516
; 
32'd126346: dataIn1 = 32'd11710
; 
32'd126347: dataIn1 = 32'd11711
; 
32'd126348: dataIn1 = 32'd541
; 
32'd126349: dataIn1 = 32'd1240
; 
32'd126350: dataIn1 = 32'd1241
; 
32'd126351: dataIn1 = 32'd1242
; 
32'd126352: dataIn1 = 32'd1243
; 
32'd126353: dataIn1 = 32'd10641
; 
32'd126354: dataIn1 = 32'd10642
; 
32'd126355: dataIn1 = 32'd10643
; 
32'd126356: dataIn1 = 32'd541
; 
32'd126357: dataIn1 = 32'd1240
; 
32'd126358: dataIn1 = 32'd1241
; 
32'd126359: dataIn1 = 32'd1244
; 
32'd126360: dataIn1 = 32'd1245
; 
32'd126361: dataIn1 = 32'd10643
; 
32'd126362: dataIn1 = 32'd10644
; 
32'd126363: dataIn1 = 32'd10645
; 
32'd126364: dataIn1 = 32'd264
; 
32'd126365: dataIn1 = 32'd1240
; 
32'd126366: dataIn1 = 32'd1242
; 
32'd126367: dataIn1 = 32'd1243
; 
32'd126368: dataIn1 = 32'd1250
; 
32'd126369: dataIn1 = 32'd10639
; 
32'd126370: dataIn1 = 32'd10640
; 
32'd126371: dataIn1 = 32'd10641
; 
32'd126372: dataIn1 = 32'd264
; 
32'd126373: dataIn1 = 32'd541
; 
32'd126374: dataIn1 = 32'd1240
; 
32'd126375: dataIn1 = 32'd1242
; 
32'd126376: dataIn1 = 32'd1243
; 
32'd126377: dataIn1 = 32'd2754
; 
32'd126378: dataIn1 = 32'd3438
; 
32'd126379: dataIn1 = 32'd265
; 
32'd126380: dataIn1 = 32'd541
; 
32'd126381: dataIn1 = 32'd1241
; 
32'd126382: dataIn1 = 32'd1244
; 
32'd126383: dataIn1 = 32'd1245
; 
32'd126384: dataIn1 = 32'd2481
; 
32'd126385: dataIn1 = 32'd2753
; 
32'd126386: dataIn1 = 32'd265
; 
32'd126387: dataIn1 = 32'd1241
; 
32'd126388: dataIn1 = 32'd1244
; 
32'd126389: dataIn1 = 32'd1245
; 
32'd126390: dataIn1 = 32'd1246
; 
32'd126391: dataIn1 = 32'd10645
; 
32'd126392: dataIn1 = 32'd10646
; 
32'd126393: dataIn1 = 32'd10647
; 
32'd126394: dataIn1 = 32'd265
; 
32'd126395: dataIn1 = 32'd1245
; 
32'd126396: dataIn1 = 32'd1246
; 
32'd126397: dataIn1 = 32'd1258
; 
32'd126398: dataIn1 = 32'd1260
; 
32'd126399: dataIn1 = 32'd10647
; 
32'd126400: dataIn1 = 32'd10648
; 
32'd126401: dataIn1 = 32'd10649
; 
32'd126402: dataIn1 = 32'd10650
; 
32'd126403: dataIn1 = 32'd543
; 
32'd126404: dataIn1 = 32'd1247
; 
32'd126405: dataIn1 = 32'd1248
; 
32'd126406: dataIn1 = 32'd1249
; 
32'd126407: dataIn1 = 32'd11727
; 
32'd126408: dataIn1 = 32'd11728
; 
32'd126409: dataIn1 = 32'd11729
; 
32'd126410: dataIn1 = 32'd542
; 
32'd126411: dataIn1 = 32'd543
; 
32'd126412: dataIn1 = 32'd1247
; 
32'd126413: dataIn1 = 32'd1248
; 
32'd126414: dataIn1 = 32'd1249
; 
32'd126415: dataIn1 = 32'd2753
; 
32'd126416: dataIn1 = 32'd2754
; 
32'd126417: dataIn1 = 32'd542
; 
32'd126418: dataIn1 = 32'd1247
; 
32'd126419: dataIn1 = 32'd1248
; 
32'd126420: dataIn1 = 32'd1249
; 
32'd126421: dataIn1 = 32'd1261
; 
32'd126422: dataIn1 = 32'd1262
; 
32'd126423: dataIn1 = 32'd11729
; 
32'd126424: dataIn1 = 32'd11730
; 
32'd126425: dataIn1 = 32'd264
; 
32'd126426: dataIn1 = 32'd1242
; 
32'd126427: dataIn1 = 32'd1250
; 
32'd126428: dataIn1 = 32'd1254
; 
32'd126429: dataIn1 = 32'd1256
; 
32'd126430: dataIn1 = 32'd10637
; 
32'd126431: dataIn1 = 32'd10638
; 
32'd126432: dataIn1 = 32'd10639
; 
32'd126433: dataIn1 = 32'd544
; 
32'd126434: dataIn1 = 32'd545
; 
32'd126435: dataIn1 = 32'd1251
; 
32'd126436: dataIn1 = 32'd3468
; 
32'd126437: dataIn1 = 32'd3474
; 
32'd126438: dataIn1 = 32'd11724
; 
32'd126439: dataIn1 = 32'd11725
; 
32'd126440: dataIn1 = 32'd531
; 
32'd126441: dataIn1 = 32'd544
; 
32'd126442: dataIn1 = 32'd1252
; 
32'd126443: dataIn1 = 32'd3478
; 
32'd126444: dataIn1 = 32'd3482
; 
32'd126445: dataIn1 = 32'd11722
; 
32'd126446: dataIn1 = 32'd11723
; 
32'd126447: dataIn1 = 32'd543
; 
32'd126448: dataIn1 = 32'd545
; 
32'd126449: dataIn1 = 32'd1253
; 
32'd126450: dataIn1 = 32'd3438
; 
32'd126451: dataIn1 = 32'd3458
; 
32'd126452: dataIn1 = 32'd11726
; 
32'd126453: dataIn1 = 32'd11727
; 
32'd126454: dataIn1 = 32'd546
; 
32'd126455: dataIn1 = 32'd1250
; 
32'd126456: dataIn1 = 32'd1254
; 
32'd126457: dataIn1 = 32'd1255
; 
32'd126458: dataIn1 = 32'd1256
; 
32'd126459: dataIn1 = 32'd10635
; 
32'd126460: dataIn1 = 32'd10636
; 
32'd126461: dataIn1 = 32'd10637
; 
32'd126462: dataIn1 = 32'd546
; 
32'd126463: dataIn1 = 32'd1216
; 
32'd126464: dataIn1 = 32'd1254
; 
32'd126465: dataIn1 = 32'd1255
; 
32'd126466: dataIn1 = 32'd1257
; 
32'd126467: dataIn1 = 32'd10633
; 
32'd126468: dataIn1 = 32'd10634
; 
32'd126469: dataIn1 = 32'd10635
; 
32'd126470: dataIn1 = 32'd264
; 
32'd126471: dataIn1 = 32'd546
; 
32'd126472: dataIn1 = 32'd1250
; 
32'd126473: dataIn1 = 32'd1254
; 
32'd126474: dataIn1 = 32'd1256
; 
32'd126475: dataIn1 = 32'd3458
; 
32'd126476: dataIn1 = 32'd3468
; 
32'd126477: dataIn1 = 32'd260
; 
32'd126478: dataIn1 = 32'd546
; 
32'd126479: dataIn1 = 32'd1216
; 
32'd126480: dataIn1 = 32'd1255
; 
32'd126481: dataIn1 = 32'd1257
; 
32'd126482: dataIn1 = 32'd3474
; 
32'd126483: dataIn1 = 32'd3478
; 
32'd126484: dataIn1 = 32'd547
; 
32'd126485: dataIn1 = 32'd1246
; 
32'd126486: dataIn1 = 32'd1258
; 
32'd126487: dataIn1 = 32'd1260
; 
32'd126488: dataIn1 = 32'd10650
; 
32'd126489: dataIn1 = 32'd10651
; 
32'd126490: dataIn1 = 32'd10652
; 
32'd126491: dataIn1 = 32'd267
; 
32'd126492: dataIn1 = 32'd547
; 
32'd126493: dataIn1 = 32'd1259
; 
32'd126494: dataIn1 = 32'd10249
; 
32'd126495: dataIn1 = 32'd10250
; 
32'd126496: dataIn1 = 32'd10652
; 
32'd126497: dataIn1 = 32'd10653
; 
32'd126498: dataIn1 = 32'd10654
; 
32'd126499: dataIn1 = 32'd265
; 
32'd126500: dataIn1 = 32'd547
; 
32'd126501: dataIn1 = 32'd1246
; 
32'd126502: dataIn1 = 32'd1258
; 
32'd126503: dataIn1 = 32'd1260
; 
32'd126504: dataIn1 = 32'd2480
; 
32'd126505: dataIn1 = 32'd2755
; 
32'd126506: dataIn1 = 32'd549
; 
32'd126507: dataIn1 = 32'd1249
; 
32'd126508: dataIn1 = 32'd1261
; 
32'd126509: dataIn1 = 32'd1262
; 
32'd126510: dataIn1 = 32'd1432
; 
32'd126511: dataIn1 = 32'd11730
; 
32'd126512: dataIn1 = 32'd11731
; 
32'd126513: dataIn1 = 32'd11732
; 
32'd126514: dataIn1 = 32'd542
; 
32'd126515: dataIn1 = 32'd549
; 
32'd126516: dataIn1 = 32'd1249
; 
32'd126517: dataIn1 = 32'd1261
; 
32'd126518: dataIn1 = 32'd1262
; 
32'd126519: dataIn1 = 32'd2482
; 
32'd126520: dataIn1 = 32'd2756
; 
32'd126521: dataIn1 = 32'd550
; 
32'd126522: dataIn1 = 32'd1263
; 
32'd126523: dataIn1 = 32'd1264
; 
32'd126524: dataIn1 = 32'd1265
; 
32'd126525: dataIn1 = 32'd10658
; 
32'd126526: dataIn1 = 32'd10659
; 
32'd126527: dataIn1 = 32'd10660
; 
32'd126528: dataIn1 = 32'd1
; 
32'd126529: dataIn1 = 32'd1263
; 
32'd126530: dataIn1 = 32'd1264
; 
32'd126531: dataIn1 = 32'd1265
; 
32'd126532: dataIn1 = 32'd1267
; 
32'd126533: dataIn1 = 32'd10660
; 
32'd126534: dataIn1 = 32'd10661
; 
32'd126535: dataIn1 = 32'd10662
; 
32'd126536: dataIn1 = 32'd1
; 
32'd126537: dataIn1 = 32'd550
; 
32'd126538: dataIn1 = 32'd959
; 
32'd126539: dataIn1 = 32'd1263
; 
32'd126540: dataIn1 = 32'd1264
; 
32'd126541: dataIn1 = 32'd1265
; 
32'd126542: dataIn1 = 32'd267
; 
32'd126543: dataIn1 = 32'd550
; 
32'd126544: dataIn1 = 32'd1266
; 
32'd126545: dataIn1 = 32'd10249
; 
32'd126546: dataIn1 = 32'd10253
; 
32'd126547: dataIn1 = 32'd10656
; 
32'd126548: dataIn1 = 32'd10657
; 
32'd126549: dataIn1 = 32'd10658
; 
32'd126550: dataIn1 = 32'd1
; 
32'd126551: dataIn1 = 32'd1264
; 
32'd126552: dataIn1 = 32'd1267
; 
32'd126553: dataIn1 = 32'd1467
; 
32'd126554: dataIn1 = 32'd1469
; 
32'd126555: dataIn1 = 32'd10662
; 
32'd126556: dataIn1 = 32'd10663
; 
32'd126557: dataIn1 = 32'd10664
; 
32'd126558: dataIn1 = 32'd10665
; 
32'd126559: dataIn1 = 32'd551
; 
32'd126560: dataIn1 = 32'd552
; 
32'd126561: dataIn1 = 32'd553
; 
32'd126562: dataIn1 = 32'd1268
; 
32'd126563: dataIn1 = 32'd11640
; 
32'd126564: dataIn1 = 32'd11641
; 
32'd126565: dataIn1 = 32'd11642
; 
32'd126566: dataIn1 = 32'd269
; 
32'd126567: dataIn1 = 32'd551
; 
32'd126568: dataIn1 = 32'd554
; 
32'd126569: dataIn1 = 32'd1269
; 
32'd126570: dataIn1 = 32'd11635
; 
32'd126571: dataIn1 = 32'd11636
; 
32'd126572: dataIn1 = 32'd11637
; 
32'd126573: dataIn1 = 32'd11638
; 
32'd126574: dataIn1 = 32'd268
; 
32'd126575: dataIn1 = 32'd553
; 
32'd126576: dataIn1 = 32'd555
; 
32'd126577: dataIn1 = 32'd1270
; 
32'd126578: dataIn1 = 32'd11644
; 
32'd126579: dataIn1 = 32'd11645
; 
32'd126580: dataIn1 = 32'd270
; 
32'd126581: dataIn1 = 32'd556
; 
32'd126582: dataIn1 = 32'd1271
; 
32'd126583: dataIn1 = 32'd10564
; 
32'd126584: dataIn1 = 32'd11660
; 
32'd126585: dataIn1 = 32'd11661
; 
32'd126586: dataIn1 = 32'd11662
; 
32'd126587: dataIn1 = 32'd556
; 
32'd126588: dataIn1 = 32'd1272
; 
32'd126589: dataIn1 = 32'd10247
; 
32'd126590: dataIn1 = 32'd10254
; 
32'd126591: dataIn1 = 32'd11657
; 
32'd126592: dataIn1 = 32'd11658
; 
32'd126593: dataIn1 = 32'd11659
; 
32'd126594: dataIn1 = 32'd555
; 
32'd126595: dataIn1 = 32'd557
; 
32'd126596: dataIn1 = 32'd1273
; 
32'd126597: dataIn1 = 32'd10248
; 
32'd126598: dataIn1 = 32'd10255
; 
32'd126599: dataIn1 = 32'd11647
; 
32'd126600: dataIn1 = 32'd11648
; 
32'd126601: dataIn1 = 32'd11649
; 
32'd126602: dataIn1 = 32'd11650
; 
32'd126603: dataIn1 = 32'd554
; 
32'd126604: dataIn1 = 32'd559
; 
32'd126605: dataIn1 = 32'd560
; 
32'd126606: dataIn1 = 32'd1274
; 
32'd126607: dataIn1 = 32'd11631
; 
32'd126608: dataIn1 = 32'd11632
; 
32'd126609: dataIn1 = 32'd11633
; 
32'd126610: dataIn1 = 32'd561
; 
32'd126611: dataIn1 = 32'd1275
; 
32'd126612: dataIn1 = 32'd1276
; 
32'd126613: dataIn1 = 32'd1277
; 
32'd126614: dataIn1 = 32'd1278
; 
32'd126615: dataIn1 = 32'd11602
; 
32'd126616: dataIn1 = 32'd11603
; 
32'd126617: dataIn1 = 32'd11604
; 
32'd126618: dataIn1 = 32'd11605
; 
32'd126619: dataIn1 = 32'd274
; 
32'd126620: dataIn1 = 32'd561
; 
32'd126621: dataIn1 = 32'd562
; 
32'd126622: dataIn1 = 32'd1275
; 
32'd126623: dataIn1 = 32'd1276
; 
32'd126624: dataIn1 = 32'd11605
; 
32'd126625: dataIn1 = 32'd273
; 
32'd126626: dataIn1 = 32'd1275
; 
32'd126627: dataIn1 = 32'd1277
; 
32'd126628: dataIn1 = 32'd1278
; 
32'd126629: dataIn1 = 32'd11600
; 
32'd126630: dataIn1 = 32'd11601
; 
32'd126631: dataIn1 = 32'd11602
; 
32'd126632: dataIn1 = 32'd273
; 
32'd126633: dataIn1 = 32'd561
; 
32'd126634: dataIn1 = 32'd1275
; 
32'd126635: dataIn1 = 32'd1277
; 
32'd126636: dataIn1 = 32'd1278
; 
32'd126637: dataIn1 = 32'd1721
; 
32'd126638: dataIn1 = 32'd274
; 
32'd126639: dataIn1 = 32'd562
; 
32'd126640: dataIn1 = 32'd563
; 
32'd126641: dataIn1 = 32'd1279
; 
32'd126642: dataIn1 = 32'd11607
; 
32'd126643: dataIn1 = 32'd11608
; 
32'd126644: dataIn1 = 32'd11609
; 
32'd126645: dataIn1 = 32'd11610
; 
32'd126646: dataIn1 = 32'd275
; 
32'd126647: dataIn1 = 32'd564
; 
32'd126648: dataIn1 = 32'd566
; 
32'd126649: dataIn1 = 32'd1280
; 
32'd126650: dataIn1 = 32'd1281
; 
32'd126651: dataIn1 = 32'd11618
; 
32'd126652: dataIn1 = 32'd11619
; 
32'd126653: dataIn1 = 32'd275
; 
32'd126654: dataIn1 = 32'd1280
; 
32'd126655: dataIn1 = 32'd1281
; 
32'd126656: dataIn1 = 32'd1282
; 
32'd126657: dataIn1 = 32'd11616
; 
32'd126658: dataIn1 = 32'd11617
; 
32'd126659: dataIn1 = 32'd11618
; 
32'd126660: dataIn1 = 32'd275
; 
32'd126661: dataIn1 = 32'd567
; 
32'd126662: dataIn1 = 32'd1281
; 
32'd126663: dataIn1 = 32'd1282
; 
32'd126664: dataIn1 = 32'd1285
; 
32'd126665: dataIn1 = 32'd11614
; 
32'd126666: dataIn1 = 32'd11615
; 
32'd126667: dataIn1 = 32'd11616
; 
32'd126668: dataIn1 = 32'd564
; 
32'd126669: dataIn1 = 32'd565
; 
32'd126670: dataIn1 = 32'd566
; 
32'd126671: dataIn1 = 32'd1283
; 
32'd126672: dataIn1 = 32'd1284
; 
32'd126673: dataIn1 = 32'd11621
; 
32'd126674: dataIn1 = 32'd565
; 
32'd126675: dataIn1 = 32'd1283
; 
32'd126676: dataIn1 = 32'd1284
; 
32'd126677: dataIn1 = 32'd1288
; 
32'd126678: dataIn1 = 32'd11621
; 
32'd126679: dataIn1 = 32'd11622
; 
32'd126680: dataIn1 = 32'd11623
; 
32'd126681: dataIn1 = 32'd563
; 
32'd126682: dataIn1 = 32'd567
; 
32'd126683: dataIn1 = 32'd1282
; 
32'd126684: dataIn1 = 32'd1285
; 
32'd126685: dataIn1 = 32'd11612
; 
32'd126686: dataIn1 = 32'd11613
; 
32'd126687: dataIn1 = 32'd11614
; 
32'd126688: dataIn1 = 32'd568
; 
32'd126689: dataIn1 = 32'd569
; 
32'd126690: dataIn1 = 32'd570
; 
32'd126691: dataIn1 = 32'd1286
; 
32'd126692: dataIn1 = 32'd11624
; 
32'd126693: dataIn1 = 32'd11625
; 
32'd126694: dataIn1 = 32'd272
; 
32'd126695: dataIn1 = 32'd560
; 
32'd126696: dataIn1 = 32'd568
; 
32'd126697: dataIn1 = 32'd1287
; 
32'd126698: dataIn1 = 32'd11627
; 
32'd126699: dataIn1 = 32'd11628
; 
32'd126700: dataIn1 = 32'd11629
; 
32'd126701: dataIn1 = 32'd565
; 
32'd126702: dataIn1 = 32'd570
; 
32'd126703: dataIn1 = 32'd571
; 
32'd126704: dataIn1 = 32'd1284
; 
32'd126705: dataIn1 = 32'd1288
; 
32'd126706: dataIn1 = 32'd11623
; 
32'd126707: dataIn1 = 32'd11624
; 
32'd126708: dataIn1 = 32'd572
; 
32'd126709: dataIn1 = 32'd1289
; 
32'd126710: dataIn1 = 32'd1290
; 
32'd126711: dataIn1 = 32'd1291
; 
32'd126712: dataIn1 = 32'd1292
; 
32'd126713: dataIn1 = 32'd11596
; 
32'd126714: dataIn1 = 32'd11597
; 
32'd126715: dataIn1 = 32'd11598
; 
32'd126716: dataIn1 = 32'd278
; 
32'd126717: dataIn1 = 32'd572
; 
32'd126718: dataIn1 = 32'd573
; 
32'd126719: dataIn1 = 32'd1289
; 
32'd126720: dataIn1 = 32'd1290
; 
32'd126721: dataIn1 = 32'd11596
; 
32'd126722: dataIn1 = 32'd273
; 
32'd126723: dataIn1 = 32'd1289
; 
32'd126724: dataIn1 = 32'd1291
; 
32'd126725: dataIn1 = 32'd1292
; 
32'd126726: dataIn1 = 32'd11598
; 
32'd126727: dataIn1 = 32'd11599
; 
32'd126728: dataIn1 = 32'd11600
; 
32'd126729: dataIn1 = 32'd273
; 
32'd126730: dataIn1 = 32'd572
; 
32'd126731: dataIn1 = 32'd1289
; 
32'd126732: dataIn1 = 32'd1291
; 
32'd126733: dataIn1 = 32'd1292
; 
32'd126734: dataIn1 = 32'd1721
; 
32'd126735: dataIn1 = 32'd278
; 
32'd126736: dataIn1 = 32'd573
; 
32'd126737: dataIn1 = 32'd574
; 
32'd126738: dataIn1 = 32'd1293
; 
32'd126739: dataIn1 = 32'd11591
; 
32'd126740: dataIn1 = 32'd11592
; 
32'd126741: dataIn1 = 32'd11593
; 
32'd126742: dataIn1 = 32'd11594
; 
32'd126743: dataIn1 = 32'd575
; 
32'd126744: dataIn1 = 32'd576
; 
32'd126745: dataIn1 = 32'd577
; 
32'd126746: dataIn1 = 32'd1294
; 
32'd126747: dataIn1 = 32'd11579
; 
32'd126748: dataIn1 = 32'd11580
; 
32'd126749: dataIn1 = 32'd11581
; 
32'd126750: dataIn1 = 32'd281
; 
32'd126751: dataIn1 = 32'd576
; 
32'd126752: dataIn1 = 32'd578
; 
32'd126753: dataIn1 = 32'd1295
; 
32'd126754: dataIn1 = 32'd11583
; 
32'd126755: dataIn1 = 32'd11584
; 
32'd126756: dataIn1 = 32'd11585
; 
32'd126757: dataIn1 = 32'd280
; 
32'd126758: dataIn1 = 32'd577
; 
32'd126759: dataIn1 = 32'd579
; 
32'd126760: dataIn1 = 32'd1296
; 
32'd126761: dataIn1 = 32'd11575
; 
32'd126762: dataIn1 = 32'd11576
; 
32'd126763: dataIn1 = 32'd11577
; 
32'd126764: dataIn1 = 32'd579
; 
32'd126765: dataIn1 = 32'd580
; 
32'd126766: dataIn1 = 32'd581
; 
32'd126767: dataIn1 = 32'd1297
; 
32'd126768: dataIn1 = 32'd11571
; 
32'd126769: dataIn1 = 32'd11572
; 
32'd126770: dataIn1 = 32'd11573
; 
32'd126771: dataIn1 = 32'd574
; 
32'd126772: dataIn1 = 32'd578
; 
32'd126773: dataIn1 = 32'd582
; 
32'd126774: dataIn1 = 32'd1298
; 
32'd126775: dataIn1 = 32'd11587
; 
32'd126776: dataIn1 = 32'd11588
; 
32'd126777: dataIn1 = 32'd11589
; 
32'd126778: dataIn1 = 32'd583
; 
32'd126779: dataIn1 = 32'd1299
; 
32'd126780: dataIn1 = 32'd2768
; 
32'd126781: dataIn1 = 32'd3054
; 
32'd126782: dataIn1 = 32'd10987
; 
32'd126783: dataIn1 = 32'd10988
; 
32'd126784: dataIn1 = 32'd10989
; 
32'd126785: dataIn1 = 32'd584
; 
32'd126786: dataIn1 = 32'd585
; 
32'd126787: dataIn1 = 32'd1300
; 
32'd126788: dataIn1 = 32'd2483
; 
32'd126789: dataIn1 = 32'd2488
; 
32'd126790: dataIn1 = 32'd10979
; 
32'd126791: dataIn1 = 32'd10980
; 
32'd126792: dataIn1 = 32'd10981
; 
32'd126793: dataIn1 = 32'd587
; 
32'd126794: dataIn1 = 32'd588
; 
32'd126795: dataIn1 = 32'd589
; 
32'd126796: dataIn1 = 32'd1301
; 
32'd126797: dataIn1 = 32'd11548
; 
32'd126798: dataIn1 = 32'd11549
; 
32'd126799: dataIn1 = 32'd288
; 
32'd126800: dataIn1 = 32'd587
; 
32'd126801: dataIn1 = 32'd590
; 
32'd126802: dataIn1 = 32'd1302
; 
32'd126803: dataIn1 = 32'd11551
; 
32'd126804: dataIn1 = 32'd11552
; 
32'd126805: dataIn1 = 32'd11553
; 
32'd126806: dataIn1 = 32'd287
; 
32'd126807: dataIn1 = 32'd589
; 
32'd126808: dataIn1 = 32'd591
; 
32'd126809: dataIn1 = 32'd1303
; 
32'd126810: dataIn1 = 32'd11544
; 
32'd126811: dataIn1 = 32'd11545
; 
32'd126812: dataIn1 = 32'd11546
; 
32'd126813: dataIn1 = 32'd591
; 
32'd126814: dataIn1 = 32'd592
; 
32'd126815: dataIn1 = 32'd593
; 
32'd126816: dataIn1 = 32'd1304
; 
32'd126817: dataIn1 = 32'd11539
; 
32'd126818: dataIn1 = 32'd11540
; 
32'd126819: dataIn1 = 32'd11541
; 
32'd126820: dataIn1 = 32'd11542
; 
32'd126821: dataIn1 = 32'd590
; 
32'd126822: dataIn1 = 32'd594
; 
32'd126823: dataIn1 = 32'd595
; 
32'd126824: dataIn1 = 32'd1305
; 
32'd126825: dataIn1 = 32'd11556
; 
32'd126826: dataIn1 = 32'd11557
; 
32'd126827: dataIn1 = 32'd11558
; 
32'd126828: dataIn1 = 32'd596
; 
32'd126829: dataIn1 = 32'd597
; 
32'd126830: dataIn1 = 32'd598
; 
32'd126831: dataIn1 = 32'd1306
; 
32'd126832: dataIn1 = 32'd11564
; 
32'd126833: dataIn1 = 32'd11565
; 
32'd126834: dataIn1 = 32'd11566
; 
32'd126835: dataIn1 = 32'd292
; 
32'd126836: dataIn1 = 32'd595
; 
32'd126837: dataIn1 = 32'd596
; 
32'd126838: dataIn1 = 32'd1307
; 
32'd126839: dataIn1 = 32'd11560
; 
32'd126840: dataIn1 = 32'd11561
; 
32'd126841: dataIn1 = 32'd11562
; 
32'd126842: dataIn1 = 32'd282
; 
32'd126843: dataIn1 = 32'd580
; 
32'd126844: dataIn1 = 32'd597
; 
32'd126845: dataIn1 = 32'd1308
; 
32'd126846: dataIn1 = 32'd11567
; 
32'd126847: dataIn1 = 32'd11568
; 
32'd126848: dataIn1 = 32'd11569
; 
32'd126849: dataIn1 = 32'd599
; 
32'd126850: dataIn1 = 32'd600
; 
32'd126851: dataIn1 = 32'd601
; 
32'd126852: dataIn1 = 32'd1309
; 
32'd126853: dataIn1 = 32'd11532
; 
32'd126854: dataIn1 = 32'd11533
; 
32'd126855: dataIn1 = 32'd11534
; 
32'd126856: dataIn1 = 32'd294
; 
32'd126857: dataIn1 = 32'd600
; 
32'd126858: dataIn1 = 32'd602
; 
32'd126859: dataIn1 = 32'd1310
; 
32'd126860: dataIn1 = 32'd11528
; 
32'd126861: dataIn1 = 32'd11529
; 
32'd126862: dataIn1 = 32'd11530
; 
32'd126863: dataIn1 = 32'd289
; 
32'd126864: dataIn1 = 32'd592
; 
32'd126865: dataIn1 = 32'd601
; 
32'd126866: dataIn1 = 32'd1311
; 
32'd126867: dataIn1 = 32'd11536
; 
32'd126868: dataIn1 = 32'd11537
; 
32'd126869: dataIn1 = 32'd603
; 
32'd126870: dataIn1 = 32'd604
; 
32'd126871: dataIn1 = 32'd605
; 
32'd126872: dataIn1 = 32'd1312
; 
32'd126873: dataIn1 = 32'd11515
; 
32'd126874: dataIn1 = 32'd11516
; 
32'd126875: dataIn1 = 32'd11517
; 
32'd126876: dataIn1 = 32'd297
; 
32'd126877: dataIn1 = 32'd604
; 
32'd126878: dataIn1 = 32'd606
; 
32'd126879: dataIn1 = 32'd1313
; 
32'd126880: dataIn1 = 32'd11519
; 
32'd126881: dataIn1 = 32'd11520
; 
32'd126882: dataIn1 = 32'd11521
; 
32'd126883: dataIn1 = 32'd296
; 
32'd126884: dataIn1 = 32'd605
; 
32'd126885: dataIn1 = 32'd607
; 
32'd126886: dataIn1 = 32'd1314
; 
32'd126887: dataIn1 = 32'd11511
; 
32'd126888: dataIn1 = 32'd11512
; 
32'd126889: dataIn1 = 32'd11513
; 
32'd126890: dataIn1 = 32'd607
; 
32'd126891: dataIn1 = 32'd608
; 
32'd126892: dataIn1 = 32'd609
; 
32'd126893: dataIn1 = 32'd1315
; 
32'd126894: dataIn1 = 32'd11507
; 
32'd126895: dataIn1 = 32'd11508
; 
32'd126896: dataIn1 = 32'd11509
; 
32'd126897: dataIn1 = 32'd602
; 
32'd126898: dataIn1 = 32'd606
; 
32'd126899: dataIn1 = 32'd610
; 
32'd126900: dataIn1 = 32'd1316
; 
32'd126901: dataIn1 = 32'd11524
; 
32'd126902: dataIn1 = 32'd11525
; 
32'd126903: dataIn1 = 32'd11526
; 
32'd126904: dataIn1 = 32'd611
; 
32'd126905: dataIn1 = 32'd612
; 
32'd126906: dataIn1 = 32'd613
; 
32'd126907: dataIn1 = 32'd1317
; 
32'd126908: dataIn1 = 32'd11484
; 
32'd126909: dataIn1 = 32'd11485
; 
32'd126910: dataIn1 = 32'd11486
; 
32'd126911: dataIn1 = 32'd304
; 
32'd126912: dataIn1 = 32'd611
; 
32'd126913: dataIn1 = 32'd614
; 
32'd126914: dataIn1 = 32'd1318
; 
32'd126915: dataIn1 = 32'd11488
; 
32'd126916: dataIn1 = 32'd11489
; 
32'd126917: dataIn1 = 32'd11490
; 
32'd126918: dataIn1 = 32'd303
; 
32'd126919: dataIn1 = 32'd613
; 
32'd126920: dataIn1 = 32'd615
; 
32'd126921: dataIn1 = 32'd1319
; 
32'd126922: dataIn1 = 32'd11480
; 
32'd126923: dataIn1 = 32'd11481
; 
32'd126924: dataIn1 = 32'd11482
; 
32'd126925: dataIn1 = 32'd615
; 
32'd126926: dataIn1 = 32'd616
; 
32'd126927: dataIn1 = 32'd617
; 
32'd126928: dataIn1 = 32'd1320
; 
32'd126929: dataIn1 = 32'd11476
; 
32'd126930: dataIn1 = 32'd11477
; 
32'd126931: dataIn1 = 32'd11478
; 
32'd126932: dataIn1 = 32'd614
; 
32'd126933: dataIn1 = 32'd618
; 
32'd126934: dataIn1 = 32'd619
; 
32'd126935: dataIn1 = 32'd1321
; 
32'd126936: dataIn1 = 32'd11492
; 
32'd126937: dataIn1 = 32'd11493
; 
32'd126938: dataIn1 = 32'd11494
; 
32'd126939: dataIn1 = 32'd620
; 
32'd126940: dataIn1 = 32'd621
; 
32'd126941: dataIn1 = 32'd622
; 
32'd126942: dataIn1 = 32'd1322
; 
32'd126943: dataIn1 = 32'd11499
; 
32'd126944: dataIn1 = 32'd11500
; 
32'd126945: dataIn1 = 32'd11501
; 
32'd126946: dataIn1 = 32'd308
; 
32'd126947: dataIn1 = 32'd619
; 
32'd126948: dataIn1 = 32'd620
; 
32'd126949: dataIn1 = 32'd1323
; 
32'd126950: dataIn1 = 32'd11496
; 
32'd126951: dataIn1 = 32'd11497
; 
32'd126952: dataIn1 = 32'd11498
; 
32'd126953: dataIn1 = 32'd298
; 
32'd126954: dataIn1 = 32'd608
; 
32'd126955: dataIn1 = 32'd621
; 
32'd126956: dataIn1 = 32'd1324
; 
32'd126957: dataIn1 = 32'd11503
; 
32'd126958: dataIn1 = 32'd11504
; 
32'd126959: dataIn1 = 32'd11505
; 
32'd126960: dataIn1 = 32'd623
; 
32'd126961: dataIn1 = 32'd624
; 
32'd126962: dataIn1 = 32'd625
; 
32'd126963: dataIn1 = 32'd1325
; 
32'd126964: dataIn1 = 32'd11468
; 
32'd126965: dataIn1 = 32'd11469
; 
32'd126966: dataIn1 = 32'd11470
; 
32'd126967: dataIn1 = 32'd310
; 
32'd126968: dataIn1 = 32'd624
; 
32'd126969: dataIn1 = 32'd626
; 
32'd126970: dataIn1 = 32'd1326
; 
32'd126971: dataIn1 = 32'd11463
; 
32'd126972: dataIn1 = 32'd11464
; 
32'd126973: dataIn1 = 32'd11465
; 
32'd126974: dataIn1 = 32'd11466
; 
32'd126975: dataIn1 = 32'd305
; 
32'd126976: dataIn1 = 32'd616
; 
32'd126977: dataIn1 = 32'd625
; 
32'd126978: dataIn1 = 32'd1327
; 
32'd126979: dataIn1 = 32'd11472
; 
32'd126980: dataIn1 = 32'd11473
; 
32'd126981: dataIn1 = 32'd11474
; 
32'd126982: dataIn1 = 32'd627
; 
32'd126983: dataIn1 = 32'd628
; 
32'd126984: dataIn1 = 32'd629
; 
32'd126985: dataIn1 = 32'd1328
; 
32'd126986: dataIn1 = 32'd11451
; 
32'd126987: dataIn1 = 32'd11452
; 
32'd126988: dataIn1 = 32'd11453
; 
32'd126989: dataIn1 = 32'd313
; 
32'd126990: dataIn1 = 32'd628
; 
32'd126991: dataIn1 = 32'd630
; 
32'd126992: dataIn1 = 32'd1329
; 
32'd126993: dataIn1 = 32'd11455
; 
32'd126994: dataIn1 = 32'd11456
; 
32'd126995: dataIn1 = 32'd11457
; 
32'd126996: dataIn1 = 32'd312
; 
32'd126997: dataIn1 = 32'd629
; 
32'd126998: dataIn1 = 32'd631
; 
32'd126999: dataIn1 = 32'd1330
; 
32'd127000: dataIn1 = 32'd11447
; 
32'd127001: dataIn1 = 32'd11448
; 
32'd127002: dataIn1 = 32'd11449
; 
32'd127003: dataIn1 = 32'd631
; 
32'd127004: dataIn1 = 32'd632
; 
32'd127005: dataIn1 = 32'd633
; 
32'd127006: dataIn1 = 32'd1331
; 
32'd127007: dataIn1 = 32'd11443
; 
32'd127008: dataIn1 = 32'd11444
; 
32'd127009: dataIn1 = 32'd11445
; 
32'd127010: dataIn1 = 32'd626
; 
32'd127011: dataIn1 = 32'd630
; 
32'd127012: dataIn1 = 32'd634
; 
32'd127013: dataIn1 = 32'd1332
; 
32'd127014: dataIn1 = 32'd11459
; 
32'd127015: dataIn1 = 32'd11460
; 
32'd127016: dataIn1 = 32'd11461
; 
32'd127017: dataIn1 = 32'd635
; 
32'd127018: dataIn1 = 32'd636
; 
32'd127019: dataIn1 = 32'd637
; 
32'd127020: dataIn1 = 32'd1333
; 
32'd127021: dataIn1 = 32'd11419
; 
32'd127022: dataIn1 = 32'd11420
; 
32'd127023: dataIn1 = 32'd11421
; 
32'd127024: dataIn1 = 32'd320
; 
32'd127025: dataIn1 = 32'd635
; 
32'd127026: dataIn1 = 32'd638
; 
32'd127027: dataIn1 = 32'd1334
; 
32'd127028: dataIn1 = 32'd11423
; 
32'd127029: dataIn1 = 32'd11424
; 
32'd127030: dataIn1 = 32'd11425
; 
32'd127031: dataIn1 = 32'd11426
; 
32'd127032: dataIn1 = 32'd319
; 
32'd127033: dataIn1 = 32'd637
; 
32'd127034: dataIn1 = 32'd639
; 
32'd127035: dataIn1 = 32'd1335
; 
32'd127036: dataIn1 = 32'd11415
; 
32'd127037: dataIn1 = 32'd11416
; 
32'd127038: dataIn1 = 32'd11417
; 
32'd127039: dataIn1 = 32'd639
; 
32'd127040: dataIn1 = 32'd640
; 
32'd127041: dataIn1 = 32'd641
; 
32'd127042: dataIn1 = 32'd1336
; 
32'd127043: dataIn1 = 32'd11411
; 
32'd127044: dataIn1 = 32'd11412
; 
32'd127045: dataIn1 = 32'd11413
; 
32'd127046: dataIn1 = 32'd11414
; 
32'd127047: dataIn1 = 32'd638
; 
32'd127048: dataIn1 = 32'd642
; 
32'd127049: dataIn1 = 32'd643
; 
32'd127050: dataIn1 = 32'd1337
; 
32'd127051: dataIn1 = 32'd11428
; 
32'd127052: dataIn1 = 32'd11429
; 
32'd127053: dataIn1 = 32'd11430
; 
32'd127054: dataIn1 = 32'd644
; 
32'd127055: dataIn1 = 32'd645
; 
32'd127056: dataIn1 = 32'd646
; 
32'd127057: dataIn1 = 32'd1338
; 
32'd127058: dataIn1 = 32'd11436
; 
32'd127059: dataIn1 = 32'd11437
; 
32'd127060: dataIn1 = 32'd11438
; 
32'd127061: dataIn1 = 32'd324
; 
32'd127062: dataIn1 = 32'd643
; 
32'd127063: dataIn1 = 32'd644
; 
32'd127064: dataIn1 = 32'd1339
; 
32'd127065: dataIn1 = 32'd11431
; 
32'd127066: dataIn1 = 32'd11432
; 
32'd127067: dataIn1 = 32'd11433
; 
32'd127068: dataIn1 = 32'd11434
; 
32'd127069: dataIn1 = 32'd314
; 
32'd127070: dataIn1 = 32'd632
; 
32'd127071: dataIn1 = 32'd645
; 
32'd127072: dataIn1 = 32'd1340
; 
32'd127073: dataIn1 = 32'd11439
; 
32'd127074: dataIn1 = 32'd11440
; 
32'd127075: dataIn1 = 32'd11441
; 
32'd127076: dataIn1 = 32'd647
; 
32'd127077: dataIn1 = 32'd648
; 
32'd127078: dataIn1 = 32'd649
; 
32'd127079: dataIn1 = 32'd1341
; 
32'd127080: dataIn1 = 32'd11403
; 
32'd127081: dataIn1 = 32'd11404
; 
32'd127082: dataIn1 = 32'd11405
; 
32'd127083: dataIn1 = 32'd326
; 
32'd127084: dataIn1 = 32'd648
; 
32'd127085: dataIn1 = 32'd650
; 
32'd127086: dataIn1 = 32'd1342
; 
32'd127087: dataIn1 = 32'd11400
; 
32'd127088: dataIn1 = 32'd11401
; 
32'd127089: dataIn1 = 32'd11402
; 
32'd127090: dataIn1 = 32'd321
; 
32'd127091: dataIn1 = 32'd640
; 
32'd127092: dataIn1 = 32'd649
; 
32'd127093: dataIn1 = 32'd1343
; 
32'd127094: dataIn1 = 32'd11407
; 
32'd127095: dataIn1 = 32'd11408
; 
32'd127096: dataIn1 = 32'd11409
; 
32'd127097: dataIn1 = 32'd651
; 
32'd127098: dataIn1 = 32'd652
; 
32'd127099: dataIn1 = 32'd653
; 
32'd127100: dataIn1 = 32'd1344
; 
32'd127101: dataIn1 = 32'd11387
; 
32'd127102: dataIn1 = 32'd11388
; 
32'd127103: dataIn1 = 32'd11389
; 
32'd127104: dataIn1 = 32'd329
; 
32'd127105: dataIn1 = 32'd652
; 
32'd127106: dataIn1 = 32'd654
; 
32'd127107: dataIn1 = 32'd1345
; 
32'd127108: dataIn1 = 32'd11391
; 
32'd127109: dataIn1 = 32'd11392
; 
32'd127110: dataIn1 = 32'd11393
; 
32'd127111: dataIn1 = 32'd11394
; 
32'd127112: dataIn1 = 32'd328
; 
32'd127113: dataIn1 = 32'd653
; 
32'd127114: dataIn1 = 32'd655
; 
32'd127115: dataIn1 = 32'd1346
; 
32'd127116: dataIn1 = 32'd11384
; 
32'd127117: dataIn1 = 32'd11385
; 
32'd127118: dataIn1 = 32'd655
; 
32'd127119: dataIn1 = 32'd656
; 
32'd127120: dataIn1 = 32'd657
; 
32'd127121: dataIn1 = 32'd1347
; 
32'd127122: dataIn1 = 32'd11380
; 
32'd127123: dataIn1 = 32'd11381
; 
32'd127124: dataIn1 = 32'd650
; 
32'd127125: dataIn1 = 32'd654
; 
32'd127126: dataIn1 = 32'd658
; 
32'd127127: dataIn1 = 32'd1348
; 
32'd127128: dataIn1 = 32'd11395
; 
32'd127129: dataIn1 = 32'd11396
; 
32'd127130: dataIn1 = 32'd11397
; 
32'd127131: dataIn1 = 32'd659
; 
32'd127132: dataIn1 = 32'd660
; 
32'd127133: dataIn1 = 32'd661
; 
32'd127134: dataIn1 = 32'd1349
; 
32'd127135: dataIn1 = 32'd11355
; 
32'd127136: dataIn1 = 32'd11356
; 
32'd127137: dataIn1 = 32'd11357
; 
32'd127138: dataIn1 = 32'd336
; 
32'd127139: dataIn1 = 32'd659
; 
32'd127140: dataIn1 = 32'd662
; 
32'd127141: dataIn1 = 32'd1350
; 
32'd127142: dataIn1 = 32'd11360
; 
32'd127143: dataIn1 = 32'd11361
; 
32'd127144: dataIn1 = 32'd11362
; 
32'd127145: dataIn1 = 32'd335
; 
32'd127146: dataIn1 = 32'd661
; 
32'd127147: dataIn1 = 32'd663
; 
32'd127148: dataIn1 = 32'd1351
; 
32'd127149: dataIn1 = 32'd11351
; 
32'd127150: dataIn1 = 32'd11352
; 
32'd127151: dataIn1 = 32'd11353
; 
32'd127152: dataIn1 = 32'd11354
; 
32'd127153: dataIn1 = 32'd663
; 
32'd127154: dataIn1 = 32'd664
; 
32'd127155: dataIn1 = 32'd665
; 
32'd127156: dataIn1 = 32'd1352
; 
32'd127157: dataIn1 = 32'd11347
; 
32'd127158: dataIn1 = 32'd11348
; 
32'd127159: dataIn1 = 32'd11349
; 
32'd127160: dataIn1 = 32'd11350
; 
32'd127161: dataIn1 = 32'd662
; 
32'd127162: dataIn1 = 32'd666
; 
32'd127163: dataIn1 = 32'd667
; 
32'd127164: dataIn1 = 32'd1353
; 
32'd127165: dataIn1 = 32'd11364
; 
32'd127166: dataIn1 = 32'd11365
; 
32'd127167: dataIn1 = 32'd668
; 
32'd127168: dataIn1 = 32'd669
; 
32'd127169: dataIn1 = 32'd670
; 
32'd127170: dataIn1 = 32'd1354
; 
32'd127171: dataIn1 = 32'd11371
; 
32'd127172: dataIn1 = 32'd11372
; 
32'd127173: dataIn1 = 32'd11373
; 
32'd127174: dataIn1 = 32'd11374
; 
32'd127175: dataIn1 = 32'd340
; 
32'd127176: dataIn1 = 32'd667
; 
32'd127177: dataIn1 = 32'd668
; 
32'd127178: dataIn1 = 32'd1355
; 
32'd127179: dataIn1 = 32'd11367
; 
32'd127180: dataIn1 = 32'd11368
; 
32'd127181: dataIn1 = 32'd11369
; 
32'd127182: dataIn1 = 32'd11370
; 
32'd127183: dataIn1 = 32'd330
; 
32'd127184: dataIn1 = 32'd656
; 
32'd127185: dataIn1 = 32'd669
; 
32'd127186: dataIn1 = 32'd1356
; 
32'd127187: dataIn1 = 32'd11375
; 
32'd127188: dataIn1 = 32'd11376
; 
32'd127189: dataIn1 = 32'd11377
; 
32'd127190: dataIn1 = 32'd11378
; 
32'd127191: dataIn1 = 32'd671
; 
32'd127192: dataIn1 = 32'd672
; 
32'd127193: dataIn1 = 32'd673
; 
32'd127194: dataIn1 = 32'd1357
; 
32'd127195: dataIn1 = 32'd11340
; 
32'd127196: dataIn1 = 32'd11341
; 
32'd127197: dataIn1 = 32'd11342
; 
32'd127198: dataIn1 = 32'd342
; 
32'd127199: dataIn1 = 32'd672
; 
32'd127200: dataIn1 = 32'd674
; 
32'd127201: dataIn1 = 32'd1358
; 
32'd127202: dataIn1 = 32'd11335
; 
32'd127203: dataIn1 = 32'd11336
; 
32'd127204: dataIn1 = 32'd11337
; 
32'd127205: dataIn1 = 32'd337
; 
32'd127206: dataIn1 = 32'd664
; 
32'd127207: dataIn1 = 32'd673
; 
32'd127208: dataIn1 = 32'd1359
; 
32'd127209: dataIn1 = 32'd11344
; 
32'd127210: dataIn1 = 32'd11345
; 
32'd127211: dataIn1 = 32'd11346
; 
32'd127212: dataIn1 = 32'd675
; 
32'd127213: dataIn1 = 32'd676
; 
32'd127214: dataIn1 = 32'd677
; 
32'd127215: dataIn1 = 32'd1360
; 
32'd127216: dataIn1 = 32'd11323
; 
32'd127217: dataIn1 = 32'd11324
; 
32'd127218: dataIn1 = 32'd11325
; 
32'd127219: dataIn1 = 32'd11326
; 
32'd127220: dataIn1 = 32'd345
; 
32'd127221: dataIn1 = 32'd676
; 
32'd127222: dataIn1 = 32'd678
; 
32'd127223: dataIn1 = 32'd1361
; 
32'd127224: dataIn1 = 32'd11327
; 
32'd127225: dataIn1 = 32'd11328
; 
32'd127226: dataIn1 = 32'd11329
; 
32'd127227: dataIn1 = 32'd11330
; 
32'd127228: dataIn1 = 32'd344
; 
32'd127229: dataIn1 = 32'd677
; 
32'd127230: dataIn1 = 32'd679
; 
32'd127231: dataIn1 = 32'd1362
; 
32'd127232: dataIn1 = 32'd11319
; 
32'd127233: dataIn1 = 32'd11320
; 
32'd127234: dataIn1 = 32'd11321
; 
32'd127235: dataIn1 = 32'd11322
; 
32'd127236: dataIn1 = 32'd679
; 
32'd127237: dataIn1 = 32'd680
; 
32'd127238: dataIn1 = 32'd681
; 
32'd127239: dataIn1 = 32'd1363
; 
32'd127240: dataIn1 = 32'd11315
; 
32'd127241: dataIn1 = 32'd11316
; 
32'd127242: dataIn1 = 32'd11317
; 
32'd127243: dataIn1 = 32'd674
; 
32'd127244: dataIn1 = 32'd678
; 
32'd127245: dataIn1 = 32'd682
; 
32'd127246: dataIn1 = 32'd1364
; 
32'd127247: dataIn1 = 32'd11332
; 
32'd127248: dataIn1 = 32'd11333
; 
32'd127249: dataIn1 = 32'd11334
; 
32'd127250: dataIn1 = 32'd683
; 
32'd127251: dataIn1 = 32'd684
; 
32'd127252: dataIn1 = 32'd685
; 
32'd127253: dataIn1 = 32'd1365
; 
32'd127254: dataIn1 = 32'd11291
; 
32'd127255: dataIn1 = 32'd11292
; 
32'd127256: dataIn1 = 32'd11293
; 
32'd127257: dataIn1 = 32'd352
; 
32'd127258: dataIn1 = 32'd683
; 
32'd127259: dataIn1 = 32'd686
; 
32'd127260: dataIn1 = 32'd1366
; 
32'd127261: dataIn1 = 32'd11295
; 
32'd127262: dataIn1 = 32'd11296
; 
32'd127263: dataIn1 = 32'd11297
; 
32'd127264: dataIn1 = 32'd11298
; 
32'd127265: dataIn1 = 32'd351
; 
32'd127266: dataIn1 = 32'd685
; 
32'd127267: dataIn1 = 32'd687
; 
32'd127268: dataIn1 = 32'd1367
; 
32'd127269: dataIn1 = 32'd11288
; 
32'd127270: dataIn1 = 32'd11289
; 
32'd127271: dataIn1 = 32'd11290
; 
32'd127272: dataIn1 = 32'd687
; 
32'd127273: dataIn1 = 32'd688
; 
32'd127274: dataIn1 = 32'd689
; 
32'd127275: dataIn1 = 32'd1368
; 
32'd127276: dataIn1 = 32'd11283
; 
32'd127277: dataIn1 = 32'd11284
; 
32'd127278: dataIn1 = 32'd11285
; 
32'd127279: dataIn1 = 32'd686
; 
32'd127280: dataIn1 = 32'd690
; 
32'd127281: dataIn1 = 32'd691
; 
32'd127282: dataIn1 = 32'd1369
; 
32'd127283: dataIn1 = 32'd11299
; 
32'd127284: dataIn1 = 32'd11300
; 
32'd127285: dataIn1 = 32'd11301
; 
32'd127286: dataIn1 = 32'd11302
; 
32'd127287: dataIn1 = 32'd692
; 
32'd127288: dataIn1 = 32'd693
; 
32'd127289: dataIn1 = 32'd694
; 
32'd127290: dataIn1 = 32'd1370
; 
32'd127291: dataIn1 = 32'd11307
; 
32'd127292: dataIn1 = 32'd11308
; 
32'd127293: dataIn1 = 32'd11309
; 
32'd127294: dataIn1 = 32'd356
; 
32'd127295: dataIn1 = 32'd691
; 
32'd127296: dataIn1 = 32'd692
; 
32'd127297: dataIn1 = 32'd1371
; 
32'd127298: dataIn1 = 32'd11303
; 
32'd127299: dataIn1 = 32'd11304
; 
32'd127300: dataIn1 = 32'd11305
; 
32'd127301: dataIn1 = 32'd11306
; 
32'd127302: dataIn1 = 32'd346
; 
32'd127303: dataIn1 = 32'd680
; 
32'd127304: dataIn1 = 32'd693
; 
32'd127305: dataIn1 = 32'd1372
; 
32'd127306: dataIn1 = 32'd11311
; 
32'd127307: dataIn1 = 32'd11312
; 
32'd127308: dataIn1 = 32'd11313
; 
32'd127309: dataIn1 = 32'd695
; 
32'd127310: dataIn1 = 32'd696
; 
32'd127311: dataIn1 = 32'd697
; 
32'd127312: dataIn1 = 32'd1373
; 
32'd127313: dataIn1 = 32'd11275
; 
32'd127314: dataIn1 = 32'd11276
; 
32'd127315: dataIn1 = 32'd11277
; 
32'd127316: dataIn1 = 32'd11278
; 
32'd127317: dataIn1 = 32'd358
; 
32'd127318: dataIn1 = 32'd696
; 
32'd127319: dataIn1 = 32'd698
; 
32'd127320: dataIn1 = 32'd1374
; 
32'd127321: dataIn1 = 32'd11271
; 
32'd127322: dataIn1 = 32'd11272
; 
32'd127323: dataIn1 = 32'd11273
; 
32'd127324: dataIn1 = 32'd11274
; 
32'd127325: dataIn1 = 32'd353
; 
32'd127326: dataIn1 = 32'd688
; 
32'd127327: dataIn1 = 32'd697
; 
32'd127328: dataIn1 = 32'd1375
; 
32'd127329: dataIn1 = 32'd11279
; 
32'd127330: dataIn1 = 32'd11280
; 
32'd127331: dataIn1 = 32'd11281
; 
32'd127332: dataIn1 = 32'd11282
; 
32'd127333: dataIn1 = 32'd699
; 
32'd127334: dataIn1 = 32'd700
; 
32'd127335: dataIn1 = 32'd701
; 
32'd127336: dataIn1 = 32'd1376
; 
32'd127337: dataIn1 = 32'd11259
; 
32'd127338: dataIn1 = 32'd11260
; 
32'd127339: dataIn1 = 32'd11261
; 
32'd127340: dataIn1 = 32'd11262
; 
32'd127341: dataIn1 = 32'd361
; 
32'd127342: dataIn1 = 32'd700
; 
32'd127343: dataIn1 = 32'd702
; 
32'd127344: dataIn1 = 32'd1377
; 
32'd127345: dataIn1 = 32'd11264
; 
32'd127346: dataIn1 = 32'd11265
; 
32'd127347: dataIn1 = 32'd360
; 
32'd127348: dataIn1 = 32'd701
; 
32'd127349: dataIn1 = 32'd703
; 
32'd127350: dataIn1 = 32'd1378
; 
32'd127351: dataIn1 = 32'd11256
; 
32'd127352: dataIn1 = 32'd11257
; 
32'd127353: dataIn1 = 32'd11258
; 
32'd127354: dataIn1 = 32'd703
; 
32'd127355: dataIn1 = 32'd704
; 
32'd127356: dataIn1 = 32'd705
; 
32'd127357: dataIn1 = 32'd1379
; 
32'd127358: dataIn1 = 32'd11251
; 
32'd127359: dataIn1 = 32'd11252
; 
32'd127360: dataIn1 = 32'd11253
; 
32'd127361: dataIn1 = 32'd11254
; 
32'd127362: dataIn1 = 32'd698
; 
32'd127363: dataIn1 = 32'd702
; 
32'd127364: dataIn1 = 32'd706
; 
32'd127365: dataIn1 = 32'd1380
; 
32'd127366: dataIn1 = 32'd11268
; 
32'd127367: dataIn1 = 32'd11269
; 
32'd127368: dataIn1 = 32'd11270
; 
32'd127369: dataIn1 = 32'd707
; 
32'd127370: dataIn1 = 32'd708
; 
32'd127371: dataIn1 = 32'd709
; 
32'd127372: dataIn1 = 32'd1381
; 
32'd127373: dataIn1 = 32'd11227
; 
32'd127374: dataIn1 = 32'd11228
; 
32'd127375: dataIn1 = 32'd11229
; 
32'd127376: dataIn1 = 32'd368
; 
32'd127377: dataIn1 = 32'd707
; 
32'd127378: dataIn1 = 32'd710
; 
32'd127379: dataIn1 = 32'd1382
; 
32'd127380: dataIn1 = 32'd11231
; 
32'd127381: dataIn1 = 32'd11232
; 
32'd127382: dataIn1 = 32'd11233
; 
32'd127383: dataIn1 = 32'd11234
; 
32'd127384: dataIn1 = 32'd367
; 
32'd127385: dataIn1 = 32'd709
; 
32'd127386: dataIn1 = 32'd711
; 
32'd127387: dataIn1 = 32'd1383
; 
32'd127388: dataIn1 = 32'd11223
; 
32'd127389: dataIn1 = 32'd11224
; 
32'd127390: dataIn1 = 32'd11225
; 
32'd127391: dataIn1 = 32'd711
; 
32'd127392: dataIn1 = 32'd712
; 
32'd127393: dataIn1 = 32'd713
; 
32'd127394: dataIn1 = 32'd1384
; 
32'd127395: dataIn1 = 32'd11220
; 
32'd127396: dataIn1 = 32'd11221
; 
32'd127397: dataIn1 = 32'd11222
; 
32'd127398: dataIn1 = 32'd710
; 
32'd127399: dataIn1 = 32'd714
; 
32'd127400: dataIn1 = 32'd715
; 
32'd127401: dataIn1 = 32'd1385
; 
32'd127402: dataIn1 = 32'd11236
; 
32'd127403: dataIn1 = 32'd11237
; 
32'd127404: dataIn1 = 32'd716
; 
32'd127405: dataIn1 = 32'd717
; 
32'd127406: dataIn1 = 32'd718
; 
32'd127407: dataIn1 = 32'd1386
; 
32'd127408: dataIn1 = 32'd11243
; 
32'd127409: dataIn1 = 32'd11244
; 
32'd127410: dataIn1 = 32'd11245
; 
32'd127411: dataIn1 = 32'd372
; 
32'd127412: dataIn1 = 32'd715
; 
32'd127413: dataIn1 = 32'd716
; 
32'd127414: dataIn1 = 32'd1387
; 
32'd127415: dataIn1 = 32'd11239
; 
32'd127416: dataIn1 = 32'd11240
; 
32'd127417: dataIn1 = 32'd11241
; 
32'd127418: dataIn1 = 32'd362
; 
32'd127419: dataIn1 = 32'd704
; 
32'd127420: dataIn1 = 32'd717
; 
32'd127421: dataIn1 = 32'd1388
; 
32'd127422: dataIn1 = 32'd11247
; 
32'd127423: dataIn1 = 32'd11248
; 
32'd127424: dataIn1 = 32'd11249
; 
32'd127425: dataIn1 = 32'd11250
; 
32'd127426: dataIn1 = 32'd719
; 
32'd127427: dataIn1 = 32'd720
; 
32'd127428: dataIn1 = 32'd721
; 
32'd127429: dataIn1 = 32'd1389
; 
32'd127430: dataIn1 = 32'd11212
; 
32'd127431: dataIn1 = 32'd11213
; 
32'd127432: dataIn1 = 32'd374
; 
32'd127433: dataIn1 = 32'd720
; 
32'd127434: dataIn1 = 32'd722
; 
32'd127435: dataIn1 = 32'd1390
; 
32'd127436: dataIn1 = 32'd11208
; 
32'd127437: dataIn1 = 32'd11209
; 
32'd127438: dataIn1 = 32'd11210
; 
32'd127439: dataIn1 = 32'd369
; 
32'd127440: dataIn1 = 32'd712
; 
32'd127441: dataIn1 = 32'd721
; 
32'd127442: dataIn1 = 32'd1391
; 
32'd127443: dataIn1 = 32'd11216
; 
32'd127444: dataIn1 = 32'd11217
; 
32'd127445: dataIn1 = 32'd376
; 
32'd127446: dataIn1 = 32'd723
; 
32'd127447: dataIn1 = 32'd724
; 
32'd127448: dataIn1 = 32'd725
; 
32'd127449: dataIn1 = 32'd1392
; 
32'd127450: dataIn1 = 32'd11202
; 
32'd127451: dataIn1 = 32'd11203
; 
32'd127452: dataIn1 = 32'd377
; 
32'd127453: dataIn1 = 32'd723
; 
32'd127454: dataIn1 = 32'd724
; 
32'd127455: dataIn1 = 32'd726
; 
32'd127456: dataIn1 = 32'd1393
; 
32'd127457: dataIn1 = 32'd11204
; 
32'd127458: dataIn1 = 32'd11205
; 
32'd127459: dataIn1 = 32'd376
; 
32'd127460: dataIn1 = 32'd725
; 
32'd127461: dataIn1 = 32'd727
; 
32'd127462: dataIn1 = 32'd729
; 
32'd127463: dataIn1 = 32'd1394
; 
32'd127464: dataIn1 = 32'd11199
; 
32'd127465: dataIn1 = 32'd11200
; 
32'd127466: dataIn1 = 32'd11201
; 
32'd127467: dataIn1 = 32'd378
; 
32'd127468: dataIn1 = 32'd727
; 
32'd127469: dataIn1 = 32'd728
; 
32'd127470: dataIn1 = 32'd729
; 
32'd127471: dataIn1 = 32'd1395
; 
32'd127472: dataIn1 = 32'd10563
; 
32'd127473: dataIn1 = 32'd11198
; 
32'd127474: dataIn1 = 32'd377
; 
32'd127475: dataIn1 = 32'd722
; 
32'd127476: dataIn1 = 32'd726
; 
32'd127477: dataIn1 = 32'd730
; 
32'd127478: dataIn1 = 32'd1396
; 
32'd127479: dataIn1 = 32'd11206
; 
32'd127480: dataIn1 = 32'd194
; 
32'd127481: dataIn1 = 32'd731
; 
32'd127482: dataIn1 = 32'd1397
; 
32'd127483: dataIn1 = 32'd1829
; 
32'd127484: dataIn1 = 32'd1830
; 
32'd127485: dataIn1 = 32'd10751
; 
32'd127486: dataIn1 = 32'd10752
; 
32'd127487: dataIn1 = 32'd10753
; 
32'd127488: dataIn1 = 32'd383
; 
32'd127489: dataIn1 = 32'd731
; 
32'd127490: dataIn1 = 32'd1398
; 
32'd127491: dataIn1 = 32'd1829
; 
32'd127492: dataIn1 = 32'd1832
; 
32'd127493: dataIn1 = 32'd10749
; 
32'd127494: dataIn1 = 32'd10750
; 
32'd127495: dataIn1 = 32'd383
; 
32'd127496: dataIn1 = 32'd732
; 
32'd127497: dataIn1 = 32'd1399
; 
32'd127498: dataIn1 = 32'd1831
; 
32'd127499: dataIn1 = 32'd1832
; 
32'd127500: dataIn1 = 32'd10747
; 
32'd127501: dataIn1 = 32'd10748
; 
32'd127502: dataIn1 = 32'd196
; 
32'd127503: dataIn1 = 32'd732
; 
32'd127504: dataIn1 = 32'd1400
; 
32'd127505: dataIn1 = 32'd1831
; 
32'd127506: dataIn1 = 32'd1839
; 
32'd127507: dataIn1 = 32'd10745
; 
32'd127508: dataIn1 = 32'd10746
; 
32'd127509: dataIn1 = 32'd194
; 
32'd127510: dataIn1 = 32'd733
; 
32'd127511: dataIn1 = 32'd1401
; 
32'd127512: dataIn1 = 32'd1830
; 
32'd127513: dataIn1 = 32'd1834
; 
32'd127514: dataIn1 = 32'd10754
; 
32'd127515: dataIn1 = 32'd384
; 
32'd127516: dataIn1 = 32'd733
; 
32'd127517: dataIn1 = 32'd1402
; 
32'd127518: dataIn1 = 32'd1833
; 
32'd127519: dataIn1 = 32'd1834
; 
32'd127520: dataIn1 = 32'd10755
; 
32'd127521: dataIn1 = 32'd10756
; 
32'd127522: dataIn1 = 32'd10757
; 
32'd127523: dataIn1 = 32'd197
; 
32'd127524: dataIn1 = 32'd734
; 
32'd127525: dataIn1 = 32'd1403
; 
32'd127526: dataIn1 = 32'd1835
; 
32'd127527: dataIn1 = 32'd1836
; 
32'd127528: dataIn1 = 32'd10760
; 
32'd127529: dataIn1 = 32'd384
; 
32'd127530: dataIn1 = 32'd734
; 
32'd127531: dataIn1 = 32'd1404
; 
32'd127532: dataIn1 = 32'd1833
; 
32'd127533: dataIn1 = 32'd1835
; 
32'd127534: dataIn1 = 32'd10758
; 
32'd127535: dataIn1 = 32'd10759
; 
32'd127536: dataIn1 = 32'd385
; 
32'd127537: dataIn1 = 32'd735
; 
32'd127538: dataIn1 = 32'd1405
; 
32'd127539: dataIn1 = 32'd1837
; 
32'd127540: dataIn1 = 32'd1838
; 
32'd127541: dataIn1 = 32'd10739
; 
32'd127542: dataIn1 = 32'd10740
; 
32'd127543: dataIn1 = 32'd198
; 
32'd127544: dataIn1 = 32'd735
; 
32'd127545: dataIn1 = 32'd1406
; 
32'd127546: dataIn1 = 32'd1837
; 
32'd127547: dataIn1 = 32'd10737
; 
32'd127548: dataIn1 = 32'd10738
; 
32'd127549: dataIn1 = 32'd385
; 
32'd127550: dataIn1 = 32'd736
; 
32'd127551: dataIn1 = 32'd1407
; 
32'd127552: dataIn1 = 32'd1838
; 
32'd127553: dataIn1 = 32'd1840
; 
32'd127554: dataIn1 = 32'd10741
; 
32'd127555: dataIn1 = 32'd10742
; 
32'd127556: dataIn1 = 32'd196
; 
32'd127557: dataIn1 = 32'd736
; 
32'd127558: dataIn1 = 32'd1408
; 
32'd127559: dataIn1 = 32'd1839
; 
32'd127560: dataIn1 = 32'd1840
; 
32'd127561: dataIn1 = 32'd10743
; 
32'd127562: dataIn1 = 32'd10744
; 
32'd127563: dataIn1 = 32'd386
; 
32'd127564: dataIn1 = 32'd737
; 
32'd127565: dataIn1 = 32'd1409
; 
32'd127566: dataIn1 = 32'd1842
; 
32'd127567: dataIn1 = 32'd10733
; 
32'd127568: dataIn1 = 32'd10734
; 
32'd127569: dataIn1 = 32'd198
; 
32'd127570: dataIn1 = 32'd737
; 
32'd127571: dataIn1 = 32'd1410
; 
32'd127572: dataIn1 = 32'd1841
; 
32'd127573: dataIn1 = 32'd10735
; 
32'd127574: dataIn1 = 32'd10736
; 
32'd127575: dataIn1 = 32'd386
; 
32'd127576: dataIn1 = 32'd738
; 
32'd127577: dataIn1 = 32'd1411
; 
32'd127578: dataIn1 = 32'd1844
; 
32'd127579: dataIn1 = 32'd10731
; 
32'd127580: dataIn1 = 32'd10732
; 
32'd127581: dataIn1 = 32'd200
; 
32'd127582: dataIn1 = 32'd738
; 
32'd127583: dataIn1 = 32'd1412
; 
32'd127584: dataIn1 = 32'd1843
; 
32'd127585: dataIn1 = 32'd10729
; 
32'd127586: dataIn1 = 32'd10730
; 
32'd127587: dataIn1 = 32'd201
; 
32'd127588: dataIn1 = 32'd739
; 
32'd127589: dataIn1 = 32'd1413
; 
32'd127590: dataIn1 = 32'd1846
; 
32'd127591: dataIn1 = 32'd10719
; 
32'd127592: dataIn1 = 32'd10720
; 
32'd127593: dataIn1 = 32'd387
; 
32'd127594: dataIn1 = 32'd739
; 
32'd127595: dataIn1 = 32'd1414
; 
32'd127596: dataIn1 = 32'd1845
; 
32'd127597: dataIn1 = 32'd10717
; 
32'd127598: dataIn1 = 32'd10718
; 
32'd127599: dataIn1 = 32'd387
; 
32'd127600: dataIn1 = 32'd740
; 
32'd127601: dataIn1 = 32'd1415
; 
32'd127602: dataIn1 = 32'd1848
; 
32'd127603: dataIn1 = 32'd10715
; 
32'd127604: dataIn1 = 32'd10716
; 
32'd127605: dataIn1 = 32'd203
; 
32'd127606: dataIn1 = 32'd740
; 
32'd127607: dataIn1 = 32'd1416
; 
32'd127608: dataIn1 = 32'd3409
; 
32'd127609: dataIn1 = 32'd3446
; 
32'd127610: dataIn1 = 32'd10713
; 
32'd127611: dataIn1 = 32'd10714
; 
32'd127612: dataIn1 = 32'd201
; 
32'd127613: dataIn1 = 32'd741
; 
32'd127614: dataIn1 = 32'd1417
; 
32'd127615: dataIn1 = 32'd1850
; 
32'd127616: dataIn1 = 32'd10721
; 
32'd127617: dataIn1 = 32'd10722
; 
32'd127618: dataIn1 = 32'd388
; 
32'd127619: dataIn1 = 32'd741
; 
32'd127620: dataIn1 = 32'd1418
; 
32'd127621: dataIn1 = 32'd1849
; 
32'd127622: dataIn1 = 32'd10723
; 
32'd127623: dataIn1 = 32'd10724
; 
32'd127624: dataIn1 = 32'd200
; 
32'd127625: dataIn1 = 32'd742
; 
32'd127626: dataIn1 = 32'd1419
; 
32'd127627: dataIn1 = 32'd1852
; 
32'd127628: dataIn1 = 32'd10727
; 
32'd127629: dataIn1 = 32'd10728
; 
32'd127630: dataIn1 = 32'd388
; 
32'd127631: dataIn1 = 32'd742
; 
32'd127632: dataIn1 = 32'd1420
; 
32'd127633: dataIn1 = 32'd1851
; 
32'd127634: dataIn1 = 32'd10725
; 
32'd127635: dataIn1 = 32'd10726
; 
32'd127636: dataIn1 = 32'd390
; 
32'd127637: dataIn1 = 32'd743
; 
32'd127638: dataIn1 = 32'd1421
; 
32'd127639: dataIn1 = 32'd1422
; 
32'd127640: dataIn1 = 32'd3462
; 
32'd127641: dataIn1 = 32'd3470
; 
32'd127642: dataIn1 = 32'd11736
; 
32'd127643: dataIn1 = 32'd11737
; 
32'd127644: dataIn1 = 32'd390
; 
32'd127645: dataIn1 = 32'd1421
; 
32'd127646: dataIn1 = 32'd1422
; 
32'd127647: dataIn1 = 32'd1423
; 
32'd127648: dataIn1 = 32'd11734
; 
32'd127649: dataIn1 = 32'd11735
; 
32'd127650: dataIn1 = 32'd11736
; 
32'd127651: dataIn1 = 32'd390
; 
32'd127652: dataIn1 = 32'd744
; 
32'd127653: dataIn1 = 32'd750
; 
32'd127654: dataIn1 = 32'd1422
; 
32'd127655: dataIn1 = 32'd1423
; 
32'd127656: dataIn1 = 32'd11734
; 
32'd127657: dataIn1 = 32'd743
; 
32'd127658: dataIn1 = 32'd746
; 
32'd127659: dataIn1 = 32'd1424
; 
32'd127660: dataIn1 = 32'd3448
; 
32'd127661: dataIn1 = 32'd3462
; 
32'd127662: dataIn1 = 32'd10560
; 
32'd127663: dataIn1 = 32'd10561
; 
32'd127664: dataIn1 = 32'd10707
; 
32'd127665: dataIn1 = 32'd389
; 
32'd127666: dataIn1 = 32'd747
; 
32'd127667: dataIn1 = 32'd1425
; 
32'd127668: dataIn1 = 32'd3027
; 
32'd127669: dataIn1 = 32'd3442
; 
32'd127670: dataIn1 = 32'd10709
; 
32'd127671: dataIn1 = 32'd10710
; 
32'd127672: dataIn1 = 32'd203
; 
32'd127673: dataIn1 = 32'd747
; 
32'd127674: dataIn1 = 32'd1426
; 
32'd127675: dataIn1 = 32'd3029
; 
32'd127676: dataIn1 = 32'd3410
; 
32'd127677: dataIn1 = 32'd10711
; 
32'd127678: dataIn1 = 32'd10712
; 
32'd127679: dataIn1 = 32'd748
; 
32'd127680: dataIn1 = 32'd1427
; 
32'd127681: dataIn1 = 32'd1428
; 
32'd127682: dataIn1 = 32'd1431
; 
32'd127683: dataIn1 = 32'd10555
; 
32'd127684: dataIn1 = 32'd10556
; 
32'd127685: dataIn1 = 32'd10557
; 
32'd127686: dataIn1 = 32'd392
; 
32'd127687: dataIn1 = 32'd748
; 
32'd127688: dataIn1 = 32'd749
; 
32'd127689: dataIn1 = 32'd1427
; 
32'd127690: dataIn1 = 32'd1428
; 
32'd127691: dataIn1 = 32'd10557
; 
32'd127692: dataIn1 = 32'd10558
; 
32'd127693: dataIn1 = 32'd389
; 
32'd127694: dataIn1 = 32'd749
; 
32'd127695: dataIn1 = 32'd1429
; 
32'd127696: dataIn1 = 32'd3442
; 
32'd127697: dataIn1 = 32'd3460
; 
32'd127698: dataIn1 = 32'd10558
; 
32'd127699: dataIn1 = 32'd10559
; 
32'd127700: dataIn1 = 32'd204
; 
32'd127701: dataIn1 = 32'd746
; 
32'd127702: dataIn1 = 32'd1430
; 
32'd127703: dataIn1 = 32'd3416
; 
32'd127704: dataIn1 = 32'd3448
; 
32'd127705: dataIn1 = 32'd10553
; 
32'd127706: dataIn1 = 32'd10554
; 
32'd127707: dataIn1 = 32'd10555
; 
32'd127708: dataIn1 = 32'd748
; 
32'd127709: dataIn1 = 32'd1427
; 
32'd127710: dataIn1 = 32'd1431
; 
32'd127711: dataIn1 = 32'd1441
; 
32'd127712: dataIn1 = 32'd1450
; 
32'd127713: dataIn1 = 32'd10553
; 
32'd127714: dataIn1 = 32'd10554
; 
32'd127715: dataIn1 = 32'd10555
; 
32'd127716: dataIn1 = 32'd549
; 
32'd127717: dataIn1 = 32'd744
; 
32'd127718: dataIn1 = 32'd750
; 
32'd127719: dataIn1 = 32'd1261
; 
32'd127720: dataIn1 = 32'd1432
; 
32'd127721: dataIn1 = 32'd11732
; 
32'd127722: dataIn1 = 32'd751
; 
32'd127723: dataIn1 = 32'd752
; 
32'd127724: dataIn1 = 32'd753
; 
32'd127725: dataIn1 = 32'd1433
; 
32'd127726: dataIn1 = 32'd1434
; 
32'd127727: dataIn1 = 32'd1435
; 
32'd127728: dataIn1 = 32'd753
; 
32'd127729: dataIn1 = 32'd1433
; 
32'd127730: dataIn1 = 32'd1434
; 
32'd127731: dataIn1 = 32'd1435
; 
32'd127732: dataIn1 = 32'd1442
; 
32'd127733: dataIn1 = 32'd10542
; 
32'd127734: dataIn1 = 32'd10543
; 
32'd127735: dataIn1 = 32'd10544
; 
32'd127736: dataIn1 = 32'd752
; 
32'd127737: dataIn1 = 32'd1433
; 
32'd127738: dataIn1 = 32'd1434
; 
32'd127739: dataIn1 = 32'd1435
; 
32'd127740: dataIn1 = 32'd1436
; 
32'd127741: dataIn1 = 32'd10544
; 
32'd127742: dataIn1 = 32'd10545
; 
32'd127743: dataIn1 = 32'd10546
; 
32'd127744: dataIn1 = 32'd752
; 
32'd127745: dataIn1 = 32'd1435
; 
32'd127746: dataIn1 = 32'd1436
; 
32'd127747: dataIn1 = 32'd1437
; 
32'd127748: dataIn1 = 32'd1438
; 
32'd127749: dataIn1 = 32'd10546
; 
32'd127750: dataIn1 = 32'd10547
; 
32'd127751: dataIn1 = 32'd10548
; 
32'd127752: dataIn1 = 32'd754
; 
32'd127753: dataIn1 = 32'd1436
; 
32'd127754: dataIn1 = 32'd1437
; 
32'd127755: dataIn1 = 32'd1438
; 
32'd127756: dataIn1 = 32'd1441
; 
32'd127757: dataIn1 = 32'd10548
; 
32'd127758: dataIn1 = 32'd10549
; 
32'd127759: dataIn1 = 32'd10550
; 
32'd127760: dataIn1 = 32'd10551
; 
32'd127761: dataIn1 = 32'd396
; 
32'd127762: dataIn1 = 32'd752
; 
32'd127763: dataIn1 = 32'd754
; 
32'd127764: dataIn1 = 32'd1436
; 
32'd127765: dataIn1 = 32'd1437
; 
32'd127766: dataIn1 = 32'd1438
; 
32'd127767: dataIn1 = 32'd394
; 
32'd127768: dataIn1 = 32'd755
; 
32'd127769: dataIn1 = 32'd1439
; 
32'd127770: dataIn1 = 32'd3032
; 
32'd127771: dataIn1 = 32'd3413
; 
32'd127772: dataIn1 = 32'd10546
; 
32'd127773: dataIn1 = 32'd10547
; 
32'd127774: dataIn1 = 32'd10548
; 
32'd127775: dataIn1 = 32'd204
; 
32'd127776: dataIn1 = 32'd755
; 
32'd127777: dataIn1 = 32'd1440
; 
32'd127778: dataIn1 = 32'd3033
; 
32'd127779: dataIn1 = 32'd3414
; 
32'd127780: dataIn1 = 32'd10550
; 
32'd127781: dataIn1 = 32'd10551
; 
32'd127782: dataIn1 = 32'd754
; 
32'd127783: dataIn1 = 32'd1431
; 
32'd127784: dataIn1 = 32'd1437
; 
32'd127785: dataIn1 = 32'd1441
; 
32'd127786: dataIn1 = 32'd1450
; 
32'd127787: dataIn1 = 32'd10551
; 
32'd127788: dataIn1 = 32'd10552
; 
32'd127789: dataIn1 = 32'd10553
; 
32'd127790: dataIn1 = 32'd753
; 
32'd127791: dataIn1 = 32'd1434
; 
32'd127792: dataIn1 = 32'd1442
; 
32'd127793: dataIn1 = 32'd1443
; 
32'd127794: dataIn1 = 32'd1444
; 
32'd127795: dataIn1 = 32'd10540
; 
32'd127796: dataIn1 = 32'd10541
; 
32'd127797: dataIn1 = 32'd10542
; 
32'd127798: dataIn1 = 32'd395
; 
32'd127799: dataIn1 = 32'd753
; 
32'd127800: dataIn1 = 32'd756
; 
32'd127801: dataIn1 = 32'd1442
; 
32'd127802: dataIn1 = 32'd1443
; 
32'd127803: dataIn1 = 32'd1444
; 
32'd127804: dataIn1 = 32'd756
; 
32'd127805: dataIn1 = 32'd1442
; 
32'd127806: dataIn1 = 32'd1443
; 
32'd127807: dataIn1 = 32'd1444
; 
32'd127808: dataIn1 = 32'd1446
; 
32'd127809: dataIn1 = 32'd10538
; 
32'd127810: dataIn1 = 32'd10539
; 
32'd127811: dataIn1 = 32'd10540
; 
32'd127812: dataIn1 = 32'd394
; 
32'd127813: dataIn1 = 32'd757
; 
32'd127814: dataIn1 = 32'd1445
; 
32'd127815: dataIn1 = 32'd3412
; 
32'd127816: dataIn1 = 32'd3447
; 
32'd127817: dataIn1 = 32'd10542
; 
32'd127818: dataIn1 = 32'd10543
; 
32'd127819: dataIn1 = 32'd10544
; 
32'd127820: dataIn1 = 32'd756
; 
32'd127821: dataIn1 = 32'd1444
; 
32'd127822: dataIn1 = 32'd1446
; 
32'd127823: dataIn1 = 32'd1448
; 
32'd127824: dataIn1 = 32'd1449
; 
32'd127825: dataIn1 = 32'd10538
; 
32'd127826: dataIn1 = 32'd10704
; 
32'd127827: dataIn1 = 32'd10705
; 
32'd127828: dataIn1 = 32'd10706
; 
32'd127829: dataIn1 = 32'd757
; 
32'd127830: dataIn1 = 32'd1447
; 
32'd127831: dataIn1 = 32'd3447
; 
32'd127832: dataIn1 = 32'd3461
; 
32'd127833: dataIn1 = 32'd10673
; 
32'd127834: dataIn1 = 32'd10674
; 
32'd127835: dataIn1 = 32'd10675
; 
32'd127836: dataIn1 = 32'd759
; 
32'd127837: dataIn1 = 32'd1446
; 
32'd127838: dataIn1 = 32'd1448
; 
32'd127839: dataIn1 = 32'd1449
; 
32'd127840: dataIn1 = 32'd1479
; 
32'd127841: dataIn1 = 32'd10703
; 
32'd127842: dataIn1 = 32'd10704
; 
32'd127843: dataIn1 = 32'd756
; 
32'd127844: dataIn1 = 32'd759
; 
32'd127845: dataIn1 = 32'd760
; 
32'd127846: dataIn1 = 32'd1446
; 
32'd127847: dataIn1 = 32'd1448
; 
32'd127848: dataIn1 = 32'd1449
; 
32'd127849: dataIn1 = 32'd748
; 
32'd127850: dataIn1 = 32'd754
; 
32'd127851: dataIn1 = 32'd761
; 
32'd127852: dataIn1 = 32'd1431
; 
32'd127853: dataIn1 = 32'd1441
; 
32'd127854: dataIn1 = 32'd1450
; 
32'd127855: dataIn1 = 32'd764
; 
32'd127856: dataIn1 = 32'd1451
; 
32'd127857: dataIn1 = 32'd1452
; 
32'd127858: dataIn1 = 32'd1453
; 
32'd127859: dataIn1 = 32'd1459
; 
32'd127860: dataIn1 = 32'd10530
; 
32'd127861: dataIn1 = 32'd10531
; 
32'd127862: dataIn1 = 32'd10532
; 
32'd127863: dataIn1 = 32'd762
; 
32'd127864: dataIn1 = 32'd763
; 
32'd127865: dataIn1 = 32'd764
; 
32'd127866: dataIn1 = 32'd1451
; 
32'd127867: dataIn1 = 32'd1452
; 
32'd127868: dataIn1 = 32'd1453
; 
32'd127869: dataIn1 = 32'd762
; 
32'd127870: dataIn1 = 32'd1451
; 
32'd127871: dataIn1 = 32'd1452
; 
32'd127872: dataIn1 = 32'd1453
; 
32'd127873: dataIn1 = 32'd1455
; 
32'd127874: dataIn1 = 32'd10532
; 
32'd127875: dataIn1 = 32'd10533
; 
32'd127876: dataIn1 = 32'd10534
; 
32'd127877: dataIn1 = 32'd765
; 
32'd127878: dataIn1 = 32'd1454
; 
32'd127879: dataIn1 = 32'd1455
; 
32'd127880: dataIn1 = 32'd1456
; 
32'd127881: dataIn1 = 32'd1457
; 
32'd127882: dataIn1 = 32'd10536
; 
32'd127883: dataIn1 = 32'd10537
; 
32'd127884: dataIn1 = 32'd10686
; 
32'd127885: dataIn1 = 32'd762
; 
32'd127886: dataIn1 = 32'd1453
; 
32'd127887: dataIn1 = 32'd1454
; 
32'd127888: dataIn1 = 32'd1455
; 
32'd127889: dataIn1 = 32'd1456
; 
32'd127890: dataIn1 = 32'd10534
; 
32'd127891: dataIn1 = 32'd10535
; 
32'd127892: dataIn1 = 32'd10536
; 
32'd127893: dataIn1 = 32'd403
; 
32'd127894: dataIn1 = 32'd762
; 
32'd127895: dataIn1 = 32'd765
; 
32'd127896: dataIn1 = 32'd1454
; 
32'd127897: dataIn1 = 32'd1455
; 
32'd127898: dataIn1 = 32'd1456
; 
32'd127899: dataIn1 = 32'd765
; 
32'd127900: dataIn1 = 32'd1454
; 
32'd127901: dataIn1 = 32'd1457
; 
32'd127902: dataIn1 = 32'd1464
; 
32'd127903: dataIn1 = 32'd1465
; 
32'd127904: dataIn1 = 32'd10686
; 
32'd127905: dataIn1 = 32'd10687
; 
32'd127906: dataIn1 = 32'd10688
; 
32'd127907: dataIn1 = 32'd402
; 
32'd127908: dataIn1 = 32'd1458
; 
32'd127909: dataIn1 = 32'd10532
; 
32'd127910: dataIn1 = 32'd10533
; 
32'd127911: dataIn1 = 32'd10534
; 
32'd127912: dataIn1 = 32'd10678
; 
32'd127913: dataIn1 = 32'd10679
; 
32'd127914: dataIn1 = 32'd764
; 
32'd127915: dataIn1 = 32'd766
; 
32'd127916: dataIn1 = 32'd767
; 
32'd127917: dataIn1 = 32'd1451
; 
32'd127918: dataIn1 = 32'd1459
; 
32'd127919: dataIn1 = 32'd10529
; 
32'd127920: dataIn1 = 32'd10530
; 
32'd127921: dataIn1 = 32'd402
; 
32'd127922: dataIn1 = 32'd1460
; 
32'd127923: dataIn1 = 32'd10527
; 
32'd127924: dataIn1 = 32'd10528
; 
32'd127925: dataIn1 = 32'd10529
; 
32'd127926: dataIn1 = 32'd10530
; 
32'd127927: dataIn1 = 32'd10681
; 
32'd127928: dataIn1 = 32'd10682
; 
32'd127929: dataIn1 = 32'd768
; 
32'd127930: dataIn1 = 32'd1461
; 
32'd127931: dataIn1 = 32'd1462
; 
32'd127932: dataIn1 = 32'd10526
; 
32'd127933: dataIn1 = 32'd10684
; 
32'd127934: dataIn1 = 32'd11671
; 
32'd127935: dataIn1 = 32'd11672
; 
32'd127936: dataIn1 = 32'd768
; 
32'd127937: dataIn1 = 32'd1461
; 
32'd127938: dataIn1 = 32'd1462
; 
32'd127939: dataIn1 = 32'd2758
; 
32'd127940: dataIn1 = 32'd3439
; 
32'd127941: dataIn1 = 32'd11669
; 
32'd127942: dataIn1 = 32'd11670
; 
32'd127943: dataIn1 = 32'd11671
; 
32'd127944: dataIn1 = 32'd207
; 
32'd127945: dataIn1 = 32'd766
; 
32'd127946: dataIn1 = 32'd767
; 
32'd127947: dataIn1 = 32'd1463
; 
32'd127948: dataIn1 = 32'd10525
; 
32'd127949: dataIn1 = 32'd10526
; 
32'd127950: dataIn1 = 32'd765
; 
32'd127951: dataIn1 = 32'd769
; 
32'd127952: dataIn1 = 32'd770
; 
32'd127953: dataIn1 = 32'd1457
; 
32'd127954: dataIn1 = 32'd1464
; 
32'd127955: dataIn1 = 32'd1465
; 
32'd127956: dataIn1 = 32'd770
; 
32'd127957: dataIn1 = 32'd1457
; 
32'd127958: dataIn1 = 32'd1464
; 
32'd127959: dataIn1 = 32'd1465
; 
32'd127960: dataIn1 = 32'd1475
; 
32'd127961: dataIn1 = 32'd10688
; 
32'd127962: dataIn1 = 32'd10689
; 
32'd127963: dataIn1 = 32'd10690
; 
32'd127964: dataIn1 = 32'd10691
; 
32'd127965: dataIn1 = 32'd397
; 
32'd127966: dataIn1 = 32'd1466
; 
32'd127967: dataIn1 = 32'd1468
; 
32'd127968: dataIn1 = 32'd1470
; 
32'd127969: dataIn1 = 32'd10669
; 
32'd127970: dataIn1 = 32'd10670
; 
32'd127971: dataIn1 = 32'd10671
; 
32'd127972: dataIn1 = 32'd771
; 
32'd127973: dataIn1 = 32'd1267
; 
32'd127974: dataIn1 = 32'd1467
; 
32'd127975: dataIn1 = 32'd1468
; 
32'd127976: dataIn1 = 32'd1469
; 
32'd127977: dataIn1 = 32'd10665
; 
32'd127978: dataIn1 = 32'd10666
; 
32'd127979: dataIn1 = 32'd10667
; 
32'd127980: dataIn1 = 32'd771
; 
32'd127981: dataIn1 = 32'd1466
; 
32'd127982: dataIn1 = 32'd1467
; 
32'd127983: dataIn1 = 32'd1468
; 
32'd127984: dataIn1 = 32'd1470
; 
32'd127985: dataIn1 = 32'd10667
; 
32'd127986: dataIn1 = 32'd10668
; 
32'd127987: dataIn1 = 32'd10669
; 
32'd127988: dataIn1 = 32'd1
; 
32'd127989: dataIn1 = 32'd771
; 
32'd127990: dataIn1 = 32'd1267
; 
32'd127991: dataIn1 = 32'd1467
; 
32'd127992: dataIn1 = 32'd1469
; 
32'd127993: dataIn1 = 32'd1859
; 
32'd127994: dataIn1 = 32'd397
; 
32'd127995: dataIn1 = 32'd771
; 
32'd127996: dataIn1 = 32'd1466
; 
32'd127997: dataIn1 = 32'd1468
; 
32'd127998: dataIn1 = 32'd1470
; 
32'd127999: dataIn1 = 32'd10259
; 
32'd128000: dataIn1 = 32'd10284
; 
32'd128001: dataIn1 = 32'd397
; 
32'd128002: dataIn1 = 32'd1471
; 
32'd128003: dataIn1 = 32'd3461
; 
32'd128004: dataIn1 = 32'd3469
; 
32'd128005: dataIn1 = 32'd10671
; 
32'd128006: dataIn1 = 32'd10672
; 
32'd128007: dataIn1 = 32'd10673
; 
32'd128008: dataIn1 = 32'd773
; 
32'd128009: dataIn1 = 32'd1472
; 
32'd128010: dataIn1 = 32'd1473
; 
32'd128011: dataIn1 = 32'd1474
; 
32'd128012: dataIn1 = 32'd1480
; 
32'd128013: dataIn1 = 32'd10697
; 
32'd128014: dataIn1 = 32'd10698
; 
32'd128015: dataIn1 = 32'd772
; 
32'd128016: dataIn1 = 32'd1472
; 
32'd128017: dataIn1 = 32'd1473
; 
32'd128018: dataIn1 = 32'd1474
; 
32'd128019: dataIn1 = 32'd1477
; 
32'd128020: dataIn1 = 32'd10695
; 
32'd128021: dataIn1 = 32'd10696
; 
32'd128022: dataIn1 = 32'd10697
; 
32'd128023: dataIn1 = 32'd772
; 
32'd128024: dataIn1 = 32'd773
; 
32'd128025: dataIn1 = 32'd774
; 
32'd128026: dataIn1 = 32'd1472
; 
32'd128027: dataIn1 = 32'd1473
; 
32'd128028: dataIn1 = 32'd1474
; 
32'd128029: dataIn1 = 32'd770
; 
32'd128030: dataIn1 = 32'd1465
; 
32'd128031: dataIn1 = 32'd1475
; 
32'd128032: dataIn1 = 32'd1476
; 
32'd128033: dataIn1 = 32'd1477
; 
32'd128034: dataIn1 = 32'd10691
; 
32'd128035: dataIn1 = 32'd10692
; 
32'd128036: dataIn1 = 32'd10693
; 
32'd128037: dataIn1 = 32'd405
; 
32'd128038: dataIn1 = 32'd770
; 
32'd128039: dataIn1 = 32'd772
; 
32'd128040: dataIn1 = 32'd1475
; 
32'd128041: dataIn1 = 32'd1476
; 
32'd128042: dataIn1 = 32'd1477
; 
32'd128043: dataIn1 = 32'd772
; 
32'd128044: dataIn1 = 32'd1473
; 
32'd128045: dataIn1 = 32'd1475
; 
32'd128046: dataIn1 = 32'd1476
; 
32'd128047: dataIn1 = 32'd1477
; 
32'd128048: dataIn1 = 32'd10693
; 
32'd128049: dataIn1 = 32'd10694
; 
32'd128050: dataIn1 = 32'd10695
; 
32'd128051: dataIn1 = 32'd398
; 
32'd128052: dataIn1 = 32'd759
; 
32'd128053: dataIn1 = 32'd773
; 
32'd128054: dataIn1 = 32'd1478
; 
32'd128055: dataIn1 = 32'd1479
; 
32'd128056: dataIn1 = 32'd1480
; 
32'd128057: dataIn1 = 32'd759
; 
32'd128058: dataIn1 = 32'd1448
; 
32'd128059: dataIn1 = 32'd1478
; 
32'd128060: dataIn1 = 32'd1479
; 
32'd128061: dataIn1 = 32'd1480
; 
32'd128062: dataIn1 = 32'd10701
; 
32'd128063: dataIn1 = 32'd10702
; 
32'd128064: dataIn1 = 32'd10703
; 
32'd128065: dataIn1 = 32'd773
; 
32'd128066: dataIn1 = 32'd1472
; 
32'd128067: dataIn1 = 32'd1478
; 
32'd128068: dataIn1 = 32'd1479
; 
32'd128069: dataIn1 = 32'd1480
; 
32'd128070: dataIn1 = 32'd10698
; 
32'd128071: dataIn1 = 32'd10699
; 
32'd128072: dataIn1 = 32'd10700
; 
32'd128073: dataIn1 = 32'd10701
; 
32'd128074: dataIn1 = 32'd776
; 
32'd128075: dataIn1 = 32'd777
; 
32'd128076: dataIn1 = 32'd1481
; 
32'd128077: dataIn1 = 32'd2492
; 
32'd128078: dataIn1 = 32'd2496
; 
32'd128079: dataIn1 = 32'd10520
; 
32'd128080: dataIn1 = 32'd10521
; 
32'd128081: dataIn1 = 32'd776
; 
32'd128082: dataIn1 = 32'd778
; 
32'd128083: dataIn1 = 32'd1482
; 
32'd128084: dataIn1 = 32'd2494
; 
32'd128085: dataIn1 = 32'd2504
; 
32'd128086: dataIn1 = 32'd10518
; 
32'd128087: dataIn1 = 32'd10519
; 
32'd128088: dataIn1 = 32'd406
; 
32'd128089: dataIn1 = 32'd779
; 
32'd128090: dataIn1 = 32'd1483
; 
32'd128091: dataIn1 = 32'd1861
; 
32'd128092: dataIn1 = 32'd10519
; 
32'd128093: dataIn1 = 32'd10520
; 
32'd128094: dataIn1 = 32'd208
; 
32'd128095: dataIn1 = 32'd779
; 
32'd128096: dataIn1 = 32'd1484
; 
32'd128097: dataIn1 = 32'd1860
; 
32'd128098: dataIn1 = 32'd10517
; 
32'd128099: dataIn1 = 32'd10518
; 
32'd128100: dataIn1 = 32'd777
; 
32'd128101: dataIn1 = 32'd780
; 
32'd128102: dataIn1 = 32'd1485
; 
32'd128103: dataIn1 = 32'd2491
; 
32'd128104: dataIn1 = 32'd2499
; 
32'd128105: dataIn1 = 32'd10522
; 
32'd128106: dataIn1 = 32'd10523
; 
32'd128107: dataIn1 = 32'd406
; 
32'd128108: dataIn1 = 32'd781
; 
32'd128109: dataIn1 = 32'd1486
; 
32'd128110: dataIn1 = 32'd1863
; 
32'd128111: dataIn1 = 32'd10521
; 
32'd128112: dataIn1 = 32'd10522
; 
32'd128113: dataIn1 = 32'd207
; 
32'd128114: dataIn1 = 32'd781
; 
32'd128115: dataIn1 = 32'd1487
; 
32'd128116: dataIn1 = 32'd1862
; 
32'd128117: dataIn1 = 32'd10523
; 
32'd128118: dataIn1 = 32'd10524
; 
32'd128119: dataIn1 = 32'd270
; 
32'd128120: dataIn1 = 32'd782
; 
32'd128121: dataIn1 = 32'd1488
; 
32'd128122: dataIn1 = 32'd10564
; 
32'd128123: dataIn1 = 32'd11663
; 
32'd128124: dataIn1 = 32'd11664
; 
32'd128125: dataIn1 = 32'd11665
; 
32'd128126: dataIn1 = 32'd782
; 
32'd128127: dataIn1 = 32'd1489
; 
32'd128128: dataIn1 = 32'd3439
; 
32'd128129: dataIn1 = 32'd3459
; 
32'd128130: dataIn1 = 32'd11666
; 
32'd128131: dataIn1 = 32'd11667
; 
32'd128132: dataIn1 = 32'd11668
; 
32'd128133: dataIn1 = 32'd768
; 
32'd128134: dataIn1 = 32'd780
; 
32'd128135: dataIn1 = 32'd1490
; 
32'd128136: dataIn1 = 32'd2498
; 
32'd128137: dataIn1 = 32'd2758
; 
32'd128138: dataIn1 = 32'd10524
; 
32'd128139: dataIn1 = 32'd10525
; 
32'd128140: dataIn1 = 32'd778
; 
32'd128141: dataIn1 = 32'd785
; 
32'd128142: dataIn1 = 32'd1491
; 
32'd128143: dataIn1 = 32'd2500
; 
32'd128144: dataIn1 = 32'd2505
; 
32'd128145: dataIn1 = 32'd10516
; 
32'd128146: dataIn1 = 32'd10517
; 
32'd128147: dataIn1 = 32'd787
; 
32'd128148: dataIn1 = 32'd788
; 
32'd128149: dataIn1 = 32'd1492
; 
32'd128150: dataIn1 = 32'd2507
; 
32'd128151: dataIn1 = 32'd2511
; 
32'd128152: dataIn1 = 32'd10512
; 
32'd128153: dataIn1 = 32'd10513
; 
32'd128154: dataIn1 = 32'd785
; 
32'd128155: dataIn1 = 32'd787
; 
32'd128156: dataIn1 = 32'd1493
; 
32'd128157: dataIn1 = 32'd2501
; 
32'd128158: dataIn1 = 32'd2509
; 
32'd128159: dataIn1 = 32'd10514
; 
32'd128160: dataIn1 = 32'd10515
; 
32'd128161: dataIn1 = 32'd410
; 
32'd128162: dataIn1 = 32'd789
; 
32'd128163: dataIn1 = 32'd1494
; 
32'd128164: dataIn1 = 32'd1865
; 
32'd128165: dataIn1 = 32'd10513
; 
32'd128166: dataIn1 = 32'd10514
; 
32'd128167: dataIn1 = 32'd208
; 
32'd128168: dataIn1 = 32'd789
; 
32'd128169: dataIn1 = 32'd1495
; 
32'd128170: dataIn1 = 32'd1864
; 
32'd128171: dataIn1 = 32'd10515
; 
32'd128172: dataIn1 = 32'd10516
; 
32'd128173: dataIn1 = 32'd788
; 
32'd128174: dataIn1 = 32'd790
; 
32'd128175: dataIn1 = 32'd1496
; 
32'd128176: dataIn1 = 32'd2506
; 
32'd128177: dataIn1 = 32'd2519
; 
32'd128178: dataIn1 = 32'd10510
; 
32'd128179: dataIn1 = 32'd10511
; 
32'd128180: dataIn1 = 32'd410
; 
32'd128181: dataIn1 = 32'd791
; 
32'd128182: dataIn1 = 32'd1497
; 
32'd128183: dataIn1 = 32'd1867
; 
32'd128184: dataIn1 = 32'd10511
; 
32'd128185: dataIn1 = 32'd10512
; 
32'd128186: dataIn1 = 32'd210
; 
32'd128187: dataIn1 = 32'd791
; 
32'd128188: dataIn1 = 32'd1498
; 
32'd128189: dataIn1 = 32'd1866
; 
32'd128190: dataIn1 = 32'd10509
; 
32'd128191: dataIn1 = 32'd10510
; 
32'd128192: dataIn1 = 32'd792
; 
32'd128193: dataIn1 = 32'd793
; 
32'd128194: dataIn1 = 32'd1499
; 
32'd128195: dataIn1 = 32'd10496
; 
32'd128196: dataIn1 = 32'd10497
; 
32'd128197: dataIn1 = 32'd10966
; 
32'd128198: dataIn1 = 32'd10967
; 
32'd128199: dataIn1 = 32'd792
; 
32'd128200: dataIn1 = 32'd794
; 
32'd128201: dataIn1 = 32'd1500
; 
32'd128202: dataIn1 = 32'd10498
; 
32'd128203: dataIn1 = 32'd10499
; 
32'd128204: dataIn1 = 32'd10968
; 
32'd128205: dataIn1 = 32'd10969
; 
32'd128206: dataIn1 = 32'd211
; 
32'd128207: dataIn1 = 32'd795
; 
32'd128208: dataIn1 = 32'd1501
; 
32'd128209: dataIn1 = 32'd3035
; 
32'd128210: dataIn1 = 32'd3444
; 
32'd128211: dataIn1 = 32'd10499
; 
32'd128212: dataIn1 = 32'd10500
; 
32'd128213: dataIn1 = 32'd412
; 
32'd128214: dataIn1 = 32'd795
; 
32'd128215: dataIn1 = 32'd1502
; 
32'd128216: dataIn1 = 32'd3036
; 
32'd128217: dataIn1 = 32'd3443
; 
32'd128218: dataIn1 = 32'd10497
; 
32'd128219: dataIn1 = 32'd10498
; 
32'd128220: dataIn1 = 32'd793
; 
32'd128221: dataIn1 = 32'd797
; 
32'd128222: dataIn1 = 32'd1503
; 
32'd128223: dataIn1 = 32'd10494
; 
32'd128224: dataIn1 = 32'd10495
; 
32'd128225: dataIn1 = 32'd10964
; 
32'd128226: dataIn1 = 32'd10965
; 
32'd128227: dataIn1 = 32'd412
; 
32'd128228: dataIn1 = 32'd796
; 
32'd128229: dataIn1 = 32'd1504
; 
32'd128230: dataIn1 = 32'd1871
; 
32'd128231: dataIn1 = 32'd10495
; 
32'd128232: dataIn1 = 32'd10496
; 
32'd128233: dataIn1 = 32'd213
; 
32'd128234: dataIn1 = 32'd796
; 
32'd128235: dataIn1 = 32'd1505
; 
32'd128236: dataIn1 = 32'd1870
; 
32'd128237: dataIn1 = 32'd10493
; 
32'd128238: dataIn1 = 32'd10494
; 
32'd128239: dataIn1 = 32'd798
; 
32'd128240: dataIn1 = 32'd799
; 
32'd128241: dataIn1 = 32'd1506
; 
32'd128242: dataIn1 = 32'd2512
; 
32'd128243: dataIn1 = 32'd2759
; 
32'd128244: dataIn1 = 32'd10504
; 
32'd128245: dataIn1 = 32'd10505
; 
32'd128246: dataIn1 = 32'd798
; 
32'd128247: dataIn1 = 32'd802
; 
32'd128248: dataIn1 = 32'd1507
; 
32'd128249: dataIn1 = 32'd1517
; 
32'd128250: dataIn1 = 32'd1872
; 
32'd128251: dataIn1 = 32'd10502
; 
32'd128252: dataIn1 = 32'd10503
; 
32'd128253: dataIn1 = 32'd211
; 
32'd128254: dataIn1 = 32'd801
; 
32'd128255: dataIn1 = 32'd1508
; 
32'd128256: dataIn1 = 32'd10262
; 
32'd128257: dataIn1 = 32'd10285
; 
32'd128258: dataIn1 = 32'd10501
; 
32'd128259: dataIn1 = 32'd10502
; 
32'd128260: dataIn1 = 32'd415
; 
32'd128261: dataIn1 = 32'd801
; 
32'd128262: dataIn1 = 32'd1509
; 
32'd128263: dataIn1 = 32'd1873
; 
32'd128264: dataIn1 = 32'd10503
; 
32'd128265: dataIn1 = 32'd10504
; 
32'd128266: dataIn1 = 32'd799
; 
32'd128267: dataIn1 = 32'd804
; 
32'd128268: dataIn1 = 32'd1510
; 
32'd128269: dataIn1 = 32'd2514
; 
32'd128270: dataIn1 = 32'd2516
; 
32'd128271: dataIn1 = 32'd10506
; 
32'd128272: dataIn1 = 32'd10507
; 
32'd128273: dataIn1 = 32'd210
; 
32'd128274: dataIn1 = 32'd803
; 
32'd128275: dataIn1 = 32'd1511
; 
32'd128276: dataIn1 = 32'd1876
; 
32'd128277: dataIn1 = 32'd10507
; 
32'd128278: dataIn1 = 32'd10508
; 
32'd128279: dataIn1 = 32'd415
; 
32'd128280: dataIn1 = 32'd803
; 
32'd128281: dataIn1 = 32'd1512
; 
32'd128282: dataIn1 = 32'd1875
; 
32'd128283: dataIn1 = 32'd10505
; 
32'd128284: dataIn1 = 32'd10506
; 
32'd128285: dataIn1 = 32'd790
; 
32'd128286: dataIn1 = 32'd804
; 
32'd128287: dataIn1 = 32'd1513
; 
32'd128288: dataIn1 = 32'd2515
; 
32'd128289: dataIn1 = 32'd2520
; 
32'd128290: dataIn1 = 32'd10508
; 
32'd128291: dataIn1 = 32'd10509
; 
32'd128292: dataIn1 = 32'd414
; 
32'd128293: dataIn1 = 32'd1514
; 
32'd128294: dataIn1 = 32'd2760
; 
32'd128295: dataIn1 = 32'd3440
; 
32'd128296: dataIn1 = 32'd10974
; 
32'd128297: dataIn1 = 32'd10975
; 
32'd128298: dataIn1 = 32'd10976
; 
32'd128299: dataIn1 = 32'd794
; 
32'd128300: dataIn1 = 32'd802
; 
32'd128301: dataIn1 = 32'd1515
; 
32'd128302: dataIn1 = 32'd1516
; 
32'd128303: dataIn1 = 32'd10500
; 
32'd128304: dataIn1 = 32'd10501
; 
32'd128305: dataIn1 = 32'd10970
; 
32'd128306: dataIn1 = 32'd802
; 
32'd128307: dataIn1 = 32'd1515
; 
32'd128308: dataIn1 = 32'd1516
; 
32'd128309: dataIn1 = 32'd1517
; 
32'd128310: dataIn1 = 32'd10970
; 
32'd128311: dataIn1 = 32'd10971
; 
32'd128312: dataIn1 = 32'd10972
; 
32'd128313: dataIn1 = 32'd10973
; 
32'd128314: dataIn1 = 32'd414
; 
32'd128315: dataIn1 = 32'd802
; 
32'd128316: dataIn1 = 32'd1507
; 
32'd128317: dataIn1 = 32'd1516
; 
32'd128318: dataIn1 = 32'd1517
; 
32'd128319: dataIn1 = 32'd1872
; 
32'd128320: dataIn1 = 32'd10973
; 
32'd128321: dataIn1 = 32'd585
; 
32'd128322: dataIn1 = 32'd1518
; 
32'd128323: dataIn1 = 32'd2522
; 
32'd128324: dataIn1 = 32'd2760
; 
32'd128325: dataIn1 = 32'd10976
; 
32'd128326: dataIn1 = 32'd10977
; 
32'd128327: dataIn1 = 32'd10978
; 
32'd128328: dataIn1 = 32'd807
; 
32'd128329: dataIn1 = 32'd808
; 
32'd128330: dataIn1 = 32'd1519
; 
32'd128331: dataIn1 = 32'd10488
; 
32'd128332: dataIn1 = 32'd10489
; 
32'd128333: dataIn1 = 32'd10958
; 
32'd128334: dataIn1 = 32'd10959
; 
32'd128335: dataIn1 = 32'd807
; 
32'd128336: dataIn1 = 32'd809
; 
32'd128337: dataIn1 = 32'd1520
; 
32'd128338: dataIn1 = 32'd10486
; 
32'd128339: dataIn1 = 32'd10487
; 
32'd128340: dataIn1 = 32'd10956
; 
32'd128341: dataIn1 = 32'd10957
; 
32'd128342: dataIn1 = 32'd417
; 
32'd128343: dataIn1 = 32'd810
; 
32'd128344: dataIn1 = 32'd1521
; 
32'd128345: dataIn1 = 32'd1878
; 
32'd128346: dataIn1 = 32'd10487
; 
32'd128347: dataIn1 = 32'd10488
; 
32'd128348: dataIn1 = 32'd214
; 
32'd128349: dataIn1 = 32'd810
; 
32'd128350: dataIn1 = 32'd1522
; 
32'd128351: dataIn1 = 32'd1877
; 
32'd128352: dataIn1 = 32'd10485
; 
32'd128353: dataIn1 = 32'd10486
; 
32'd128354: dataIn1 = 32'd808
; 
32'd128355: dataIn1 = 32'd811
; 
32'd128356: dataIn1 = 32'd1523
; 
32'd128357: dataIn1 = 32'd10490
; 
32'd128358: dataIn1 = 32'd10491
; 
32'd128359: dataIn1 = 32'd10960
; 
32'd128360: dataIn1 = 32'd10961
; 
32'd128361: dataIn1 = 32'd417
; 
32'd128362: dataIn1 = 32'd812
; 
32'd128363: dataIn1 = 32'd1524
; 
32'd128364: dataIn1 = 32'd1880
; 
32'd128365: dataIn1 = 32'd10489
; 
32'd128366: dataIn1 = 32'd10490
; 
32'd128367: dataIn1 = 32'd213
; 
32'd128368: dataIn1 = 32'd812
; 
32'd128369: dataIn1 = 32'd1525
; 
32'd128370: dataIn1 = 32'd1879
; 
32'd128371: dataIn1 = 32'd10491
; 
32'd128372: dataIn1 = 32'd10492
; 
32'd128373: dataIn1 = 32'd797
; 
32'd128374: dataIn1 = 32'd811
; 
32'd128375: dataIn1 = 32'd1526
; 
32'd128376: dataIn1 = 32'd10492
; 
32'd128377: dataIn1 = 32'd10493
; 
32'd128378: dataIn1 = 32'd10962
; 
32'd128379: dataIn1 = 32'd10963
; 
32'd128380: dataIn1 = 32'd809
; 
32'd128381: dataIn1 = 32'd813
; 
32'd128382: dataIn1 = 32'd1527
; 
32'd128383: dataIn1 = 32'd10484
; 
32'd128384: dataIn1 = 32'd10485
; 
32'd128385: dataIn1 = 32'd10954
; 
32'd128386: dataIn1 = 32'd10955
; 
32'd128387: dataIn1 = 32'd814
; 
32'd128388: dataIn1 = 32'd815
; 
32'd128389: dataIn1 = 32'd1528
; 
32'd128390: dataIn1 = 32'd10480
; 
32'd128391: dataIn1 = 32'd10481
; 
32'd128392: dataIn1 = 32'd10950
; 
32'd128393: dataIn1 = 32'd10951
; 
32'd128394: dataIn1 = 32'd813
; 
32'd128395: dataIn1 = 32'd814
; 
32'd128396: dataIn1 = 32'd1529
; 
32'd128397: dataIn1 = 32'd10482
; 
32'd128398: dataIn1 = 32'd10483
; 
32'd128399: dataIn1 = 32'd10952
; 
32'd128400: dataIn1 = 32'd10953
; 
32'd128401: dataIn1 = 32'd418
; 
32'd128402: dataIn1 = 32'd816
; 
32'd128403: dataIn1 = 32'd1530
; 
32'd128404: dataIn1 = 32'd1882
; 
32'd128405: dataIn1 = 32'd10481
; 
32'd128406: dataIn1 = 32'd10482
; 
32'd128407: dataIn1 = 32'd214
; 
32'd128408: dataIn1 = 32'd816
; 
32'd128409: dataIn1 = 32'd1531
; 
32'd128410: dataIn1 = 32'd1881
; 
32'd128411: dataIn1 = 32'd10483
; 
32'd128412: dataIn1 = 32'd10484
; 
32'd128413: dataIn1 = 32'd815
; 
32'd128414: dataIn1 = 32'd817
; 
32'd128415: dataIn1 = 32'd1532
; 
32'd128416: dataIn1 = 32'd10478
; 
32'd128417: dataIn1 = 32'd10479
; 
32'd128418: dataIn1 = 32'd10948
; 
32'd128419: dataIn1 = 32'd10949
; 
32'd128420: dataIn1 = 32'd418
; 
32'd128421: dataIn1 = 32'd818
; 
32'd128422: dataIn1 = 32'd1533
; 
32'd128423: dataIn1 = 32'd1884
; 
32'd128424: dataIn1 = 32'd10479
; 
32'd128425: dataIn1 = 32'd10480
; 
32'd128426: dataIn1 = 32'd216
; 
32'd128427: dataIn1 = 32'd818
; 
32'd128428: dataIn1 = 32'd1534
; 
32'd128429: dataIn1 = 32'd1883
; 
32'd128430: dataIn1 = 32'd10477
; 
32'd128431: dataIn1 = 32'd10478
; 
32'd128432: dataIn1 = 32'd819
; 
32'd128433: dataIn1 = 32'd820
; 
32'd128434: dataIn1 = 32'd1535
; 
32'd128435: dataIn1 = 32'd10464
; 
32'd128436: dataIn1 = 32'd10465
; 
32'd128437: dataIn1 = 32'd10934
; 
32'd128438: dataIn1 = 32'd10935
; 
32'd128439: dataIn1 = 32'd819
; 
32'd128440: dataIn1 = 32'd821
; 
32'd128441: dataIn1 = 32'd1536
; 
32'd128442: dataIn1 = 32'd10466
; 
32'd128443: dataIn1 = 32'd10467
; 
32'd128444: dataIn1 = 32'd10936
; 
32'd128445: dataIn1 = 32'd10937
; 
32'd128446: dataIn1 = 32'd217
; 
32'd128447: dataIn1 = 32'd822
; 
32'd128448: dataIn1 = 32'd1537
; 
32'd128449: dataIn1 = 32'd1886
; 
32'd128450: dataIn1 = 32'd10467
; 
32'd128451: dataIn1 = 32'd10468
; 
32'd128452: dataIn1 = 32'd419
; 
32'd128453: dataIn1 = 32'd822
; 
32'd128454: dataIn1 = 32'd1538
; 
32'd128455: dataIn1 = 32'd1885
; 
32'd128456: dataIn1 = 32'd10465
; 
32'd128457: dataIn1 = 32'd10466
; 
32'd128458: dataIn1 = 32'd820
; 
32'd128459: dataIn1 = 32'd824
; 
32'd128460: dataIn1 = 32'd1539
; 
32'd128461: dataIn1 = 32'd10462
; 
32'd128462: dataIn1 = 32'd10463
; 
32'd128463: dataIn1 = 32'd10932
; 
32'd128464: dataIn1 = 32'd10933
; 
32'd128465: dataIn1 = 32'd419
; 
32'd128466: dataIn1 = 32'd823
; 
32'd128467: dataIn1 = 32'd1540
; 
32'd128468: dataIn1 = 32'd1888
; 
32'd128469: dataIn1 = 32'd10463
; 
32'd128470: dataIn1 = 32'd10464
; 
32'd128471: dataIn1 = 32'd219
; 
32'd128472: dataIn1 = 32'd823
; 
32'd128473: dataIn1 = 32'd1541
; 
32'd128474: dataIn1 = 32'd1887
; 
32'd128475: dataIn1 = 32'd10461
; 
32'd128476: dataIn1 = 32'd10462
; 
32'd128477: dataIn1 = 32'd825
; 
32'd128478: dataIn1 = 32'd826
; 
32'd128479: dataIn1 = 32'd1542
; 
32'd128480: dataIn1 = 32'd10472
; 
32'd128481: dataIn1 = 32'd10473
; 
32'd128482: dataIn1 = 32'd10942
; 
32'd128483: dataIn1 = 32'd10943
; 
32'd128484: dataIn1 = 32'd825
; 
32'd128485: dataIn1 = 32'd828
; 
32'd128486: dataIn1 = 32'd1543
; 
32'd128487: dataIn1 = 32'd10470
; 
32'd128488: dataIn1 = 32'd10471
; 
32'd128489: dataIn1 = 32'd10940
; 
32'd128490: dataIn1 = 32'd10941
; 
32'd128491: dataIn1 = 32'd217
; 
32'd128492: dataIn1 = 32'd827
; 
32'd128493: dataIn1 = 32'd1544
; 
32'd128494: dataIn1 = 32'd1890
; 
32'd128495: dataIn1 = 32'd10469
; 
32'd128496: dataIn1 = 32'd10470
; 
32'd128497: dataIn1 = 32'd420
; 
32'd128498: dataIn1 = 32'd827
; 
32'd128499: dataIn1 = 32'd1545
; 
32'd128500: dataIn1 = 32'd1889
; 
32'd128501: dataIn1 = 32'd10471
; 
32'd128502: dataIn1 = 32'd10472
; 
32'd128503: dataIn1 = 32'd826
; 
32'd128504: dataIn1 = 32'd830
; 
32'd128505: dataIn1 = 32'd1546
; 
32'd128506: dataIn1 = 32'd10474
; 
32'd128507: dataIn1 = 32'd10475
; 
32'd128508: dataIn1 = 32'd10944
; 
32'd128509: dataIn1 = 32'd10945
; 
32'd128510: dataIn1 = 32'd216
; 
32'd128511: dataIn1 = 32'd829
; 
32'd128512: dataIn1 = 32'd1547
; 
32'd128513: dataIn1 = 32'd1892
; 
32'd128514: dataIn1 = 32'd10475
; 
32'd128515: dataIn1 = 32'd10476
; 
32'd128516: dataIn1 = 32'd420
; 
32'd128517: dataIn1 = 32'd829
; 
32'd128518: dataIn1 = 32'd1548
; 
32'd128519: dataIn1 = 32'd1891
; 
32'd128520: dataIn1 = 32'd10473
; 
32'd128521: dataIn1 = 32'd10474
; 
32'd128522: dataIn1 = 32'd817
; 
32'd128523: dataIn1 = 32'd830
; 
32'd128524: dataIn1 = 32'd1549
; 
32'd128525: dataIn1 = 32'd10476
; 
32'd128526: dataIn1 = 32'd10477
; 
32'd128527: dataIn1 = 32'd10946
; 
32'd128528: dataIn1 = 32'd10947
; 
32'd128529: dataIn1 = 32'd821
; 
32'd128530: dataIn1 = 32'd828
; 
32'd128531: dataIn1 = 32'd1550
; 
32'd128532: dataIn1 = 32'd10468
; 
32'd128533: dataIn1 = 32'd10469
; 
32'd128534: dataIn1 = 32'd10938
; 
32'd128535: dataIn1 = 32'd10939
; 
32'd128536: dataIn1 = 32'd831
; 
32'd128537: dataIn1 = 32'd832
; 
32'd128538: dataIn1 = 32'd1551
; 
32'd128539: dataIn1 = 32'd10456
; 
32'd128540: dataIn1 = 32'd10457
; 
32'd128541: dataIn1 = 32'd10926
; 
32'd128542: dataIn1 = 32'd10927
; 
32'd128543: dataIn1 = 32'd831
; 
32'd128544: dataIn1 = 32'd833
; 
32'd128545: dataIn1 = 32'd1552
; 
32'd128546: dataIn1 = 32'd10454
; 
32'd128547: dataIn1 = 32'd10455
; 
32'd128548: dataIn1 = 32'd10924
; 
32'd128549: dataIn1 = 32'd10925
; 
32'd128550: dataIn1 = 32'd421
; 
32'd128551: dataIn1 = 32'd834
; 
32'd128552: dataIn1 = 32'd1553
; 
32'd128553: dataIn1 = 32'd1894
; 
32'd128554: dataIn1 = 32'd10455
; 
32'd128555: dataIn1 = 32'd10456
; 
32'd128556: dataIn1 = 32'd220
; 
32'd128557: dataIn1 = 32'd834
; 
32'd128558: dataIn1 = 32'd1554
; 
32'd128559: dataIn1 = 32'd1893
; 
32'd128560: dataIn1 = 32'd10453
; 
32'd128561: dataIn1 = 32'd10454
; 
32'd128562: dataIn1 = 32'd832
; 
32'd128563: dataIn1 = 32'd835
; 
32'd128564: dataIn1 = 32'd1555
; 
32'd128565: dataIn1 = 32'd10458
; 
32'd128566: dataIn1 = 32'd10459
; 
32'd128567: dataIn1 = 32'd10928
; 
32'd128568: dataIn1 = 32'd10929
; 
32'd128569: dataIn1 = 32'd421
; 
32'd128570: dataIn1 = 32'd836
; 
32'd128571: dataIn1 = 32'd1556
; 
32'd128572: dataIn1 = 32'd1896
; 
32'd128573: dataIn1 = 32'd10457
; 
32'd128574: dataIn1 = 32'd10458
; 
32'd128575: dataIn1 = 32'd219
; 
32'd128576: dataIn1 = 32'd836
; 
32'd128577: dataIn1 = 32'd1557
; 
32'd128578: dataIn1 = 32'd1895
; 
32'd128579: dataIn1 = 32'd10459
; 
32'd128580: dataIn1 = 32'd10460
; 
32'd128581: dataIn1 = 32'd824
; 
32'd128582: dataIn1 = 32'd835
; 
32'd128583: dataIn1 = 32'd1558
; 
32'd128584: dataIn1 = 32'd10460
; 
32'd128585: dataIn1 = 32'd10461
; 
32'd128586: dataIn1 = 32'd10930
; 
32'd128587: dataIn1 = 32'd10931
; 
32'd128588: dataIn1 = 32'd833
; 
32'd128589: dataIn1 = 32'd837
; 
32'd128590: dataIn1 = 32'd1559
; 
32'd128591: dataIn1 = 32'd10452
; 
32'd128592: dataIn1 = 32'd10453
; 
32'd128593: dataIn1 = 32'd10922
; 
32'd128594: dataIn1 = 32'd10923
; 
32'd128595: dataIn1 = 32'd838
; 
32'd128596: dataIn1 = 32'd839
; 
32'd128597: dataIn1 = 32'd1560
; 
32'd128598: dataIn1 = 32'd10448
; 
32'd128599: dataIn1 = 32'd10449
; 
32'd128600: dataIn1 = 32'd10918
; 
32'd128601: dataIn1 = 32'd10919
; 
32'd128602: dataIn1 = 32'd837
; 
32'd128603: dataIn1 = 32'd838
; 
32'd128604: dataIn1 = 32'd1561
; 
32'd128605: dataIn1 = 32'd10450
; 
32'd128606: dataIn1 = 32'd10451
; 
32'd128607: dataIn1 = 32'd10920
; 
32'd128608: dataIn1 = 32'd10921
; 
32'd128609: dataIn1 = 32'd422
; 
32'd128610: dataIn1 = 32'd840
; 
32'd128611: dataIn1 = 32'd1562
; 
32'd128612: dataIn1 = 32'd1898
; 
32'd128613: dataIn1 = 32'd10449
; 
32'd128614: dataIn1 = 32'd10450
; 
32'd128615: dataIn1 = 32'd220
; 
32'd128616: dataIn1 = 32'd840
; 
32'd128617: dataIn1 = 32'd1563
; 
32'd128618: dataIn1 = 32'd1897
; 
32'd128619: dataIn1 = 32'd10451
; 
32'd128620: dataIn1 = 32'd10452
; 
32'd128621: dataIn1 = 32'd839
; 
32'd128622: dataIn1 = 32'd841
; 
32'd128623: dataIn1 = 32'd1564
; 
32'd128624: dataIn1 = 32'd10446
; 
32'd128625: dataIn1 = 32'd10447
; 
32'd128626: dataIn1 = 32'd10916
; 
32'd128627: dataIn1 = 32'd10917
; 
32'd128628: dataIn1 = 32'd422
; 
32'd128629: dataIn1 = 32'd842
; 
32'd128630: dataIn1 = 32'd1565
; 
32'd128631: dataIn1 = 32'd1900
; 
32'd128632: dataIn1 = 32'd10447
; 
32'd128633: dataIn1 = 32'd10448
; 
32'd128634: dataIn1 = 32'd222
; 
32'd128635: dataIn1 = 32'd842
; 
32'd128636: dataIn1 = 32'd1566
; 
32'd128637: dataIn1 = 32'd1899
; 
32'd128638: dataIn1 = 32'd10445
; 
32'd128639: dataIn1 = 32'd10446
; 
32'd128640: dataIn1 = 32'd843
; 
32'd128641: dataIn1 = 32'd844
; 
32'd128642: dataIn1 = 32'd1567
; 
32'd128643: dataIn1 = 32'd10432
; 
32'd128644: dataIn1 = 32'd10433
; 
32'd128645: dataIn1 = 32'd10902
; 
32'd128646: dataIn1 = 32'd10903
; 
32'd128647: dataIn1 = 32'd843
; 
32'd128648: dataIn1 = 32'd845
; 
32'd128649: dataIn1 = 32'd1568
; 
32'd128650: dataIn1 = 32'd10434
; 
32'd128651: dataIn1 = 32'd10435
; 
32'd128652: dataIn1 = 32'd10904
; 
32'd128653: dataIn1 = 32'd10905
; 
32'd128654: dataIn1 = 32'd223
; 
32'd128655: dataIn1 = 32'd846
; 
32'd128656: dataIn1 = 32'd1569
; 
32'd128657: dataIn1 = 32'd1902
; 
32'd128658: dataIn1 = 32'd10435
; 
32'd128659: dataIn1 = 32'd10436
; 
32'd128660: dataIn1 = 32'd423
; 
32'd128661: dataIn1 = 32'd846
; 
32'd128662: dataIn1 = 32'd1570
; 
32'd128663: dataIn1 = 32'd1901
; 
32'd128664: dataIn1 = 32'd10433
; 
32'd128665: dataIn1 = 32'd10434
; 
32'd128666: dataIn1 = 32'd844
; 
32'd128667: dataIn1 = 32'd848
; 
32'd128668: dataIn1 = 32'd1571
; 
32'd128669: dataIn1 = 32'd10430
; 
32'd128670: dataIn1 = 32'd10431
; 
32'd128671: dataIn1 = 32'd10900
; 
32'd128672: dataIn1 = 32'd10901
; 
32'd128673: dataIn1 = 32'd423
; 
32'd128674: dataIn1 = 32'd847
; 
32'd128675: dataIn1 = 32'd1572
; 
32'd128676: dataIn1 = 32'd1904
; 
32'd128677: dataIn1 = 32'd10431
; 
32'd128678: dataIn1 = 32'd10432
; 
32'd128679: dataIn1 = 32'd225
; 
32'd128680: dataIn1 = 32'd847
; 
32'd128681: dataIn1 = 32'd1573
; 
32'd128682: dataIn1 = 32'd1903
; 
32'd128683: dataIn1 = 32'd10429
; 
32'd128684: dataIn1 = 32'd10430
; 
32'd128685: dataIn1 = 32'd849
; 
32'd128686: dataIn1 = 32'd850
; 
32'd128687: dataIn1 = 32'd1574
; 
32'd128688: dataIn1 = 32'd10440
; 
32'd128689: dataIn1 = 32'd10441
; 
32'd128690: dataIn1 = 32'd10910
; 
32'd128691: dataIn1 = 32'd10911
; 
32'd128692: dataIn1 = 32'd849
; 
32'd128693: dataIn1 = 32'd852
; 
32'd128694: dataIn1 = 32'd1575
; 
32'd128695: dataIn1 = 32'd10438
; 
32'd128696: dataIn1 = 32'd10439
; 
32'd128697: dataIn1 = 32'd10908
; 
32'd128698: dataIn1 = 32'd10909
; 
32'd128699: dataIn1 = 32'd223
; 
32'd128700: dataIn1 = 32'd851
; 
32'd128701: dataIn1 = 32'd1576
; 
32'd128702: dataIn1 = 32'd1906
; 
32'd128703: dataIn1 = 32'd10437
; 
32'd128704: dataIn1 = 32'd10438
; 
32'd128705: dataIn1 = 32'd424
; 
32'd128706: dataIn1 = 32'd851
; 
32'd128707: dataIn1 = 32'd1577
; 
32'd128708: dataIn1 = 32'd1905
; 
32'd128709: dataIn1 = 32'd10439
; 
32'd128710: dataIn1 = 32'd10440
; 
32'd128711: dataIn1 = 32'd850
; 
32'd128712: dataIn1 = 32'd854
; 
32'd128713: dataIn1 = 32'd1578
; 
32'd128714: dataIn1 = 32'd10442
; 
32'd128715: dataIn1 = 32'd10443
; 
32'd128716: dataIn1 = 32'd10912
; 
32'd128717: dataIn1 = 32'd10913
; 
32'd128718: dataIn1 = 32'd222
; 
32'd128719: dataIn1 = 32'd853
; 
32'd128720: dataIn1 = 32'd1579
; 
32'd128721: dataIn1 = 32'd1908
; 
32'd128722: dataIn1 = 32'd10443
; 
32'd128723: dataIn1 = 32'd10444
; 
32'd128724: dataIn1 = 32'd424
; 
32'd128725: dataIn1 = 32'd853
; 
32'd128726: dataIn1 = 32'd1580
; 
32'd128727: dataIn1 = 32'd1907
; 
32'd128728: dataIn1 = 32'd10441
; 
32'd128729: dataIn1 = 32'd10442
; 
32'd128730: dataIn1 = 32'd841
; 
32'd128731: dataIn1 = 32'd854
; 
32'd128732: dataIn1 = 32'd1581
; 
32'd128733: dataIn1 = 32'd10444
; 
32'd128734: dataIn1 = 32'd10445
; 
32'd128735: dataIn1 = 32'd10914
; 
32'd128736: dataIn1 = 32'd10915
; 
32'd128737: dataIn1 = 32'd845
; 
32'd128738: dataIn1 = 32'd852
; 
32'd128739: dataIn1 = 32'd1582
; 
32'd128740: dataIn1 = 32'd10436
; 
32'd128741: dataIn1 = 32'd10437
; 
32'd128742: dataIn1 = 32'd10906
; 
32'd128743: dataIn1 = 32'd10907
; 
32'd128744: dataIn1 = 32'd855
; 
32'd128745: dataIn1 = 32'd856
; 
32'd128746: dataIn1 = 32'd1583
; 
32'd128747: dataIn1 = 32'd10424
; 
32'd128748: dataIn1 = 32'd10425
; 
32'd128749: dataIn1 = 32'd10894
; 
32'd128750: dataIn1 = 32'd10895
; 
32'd128751: dataIn1 = 32'd855
; 
32'd128752: dataIn1 = 32'd857
; 
32'd128753: dataIn1 = 32'd1584
; 
32'd128754: dataIn1 = 32'd10422
; 
32'd128755: dataIn1 = 32'd10423
; 
32'd128756: dataIn1 = 32'd10892
; 
32'd128757: dataIn1 = 32'd10893
; 
32'd128758: dataIn1 = 32'd425
; 
32'd128759: dataIn1 = 32'd858
; 
32'd128760: dataIn1 = 32'd1585
; 
32'd128761: dataIn1 = 32'd1910
; 
32'd128762: dataIn1 = 32'd10423
; 
32'd128763: dataIn1 = 32'd10424
; 
32'd128764: dataIn1 = 32'd226
; 
32'd128765: dataIn1 = 32'd858
; 
32'd128766: dataIn1 = 32'd1586
; 
32'd128767: dataIn1 = 32'd1909
; 
32'd128768: dataIn1 = 32'd10421
; 
32'd128769: dataIn1 = 32'd10422
; 
32'd128770: dataIn1 = 32'd856
; 
32'd128771: dataIn1 = 32'd859
; 
32'd128772: dataIn1 = 32'd1587
; 
32'd128773: dataIn1 = 32'd10426
; 
32'd128774: dataIn1 = 32'd10427
; 
32'd128775: dataIn1 = 32'd10896
; 
32'd128776: dataIn1 = 32'd10897
; 
32'd128777: dataIn1 = 32'd425
; 
32'd128778: dataIn1 = 32'd860
; 
32'd128779: dataIn1 = 32'd1588
; 
32'd128780: dataIn1 = 32'd1912
; 
32'd128781: dataIn1 = 32'd10425
; 
32'd128782: dataIn1 = 32'd10426
; 
32'd128783: dataIn1 = 32'd225
; 
32'd128784: dataIn1 = 32'd860
; 
32'd128785: dataIn1 = 32'd1589
; 
32'd128786: dataIn1 = 32'd1911
; 
32'd128787: dataIn1 = 32'd10427
; 
32'd128788: dataIn1 = 32'd10428
; 
32'd128789: dataIn1 = 32'd848
; 
32'd128790: dataIn1 = 32'd859
; 
32'd128791: dataIn1 = 32'd1590
; 
32'd128792: dataIn1 = 32'd10428
; 
32'd128793: dataIn1 = 32'd10429
; 
32'd128794: dataIn1 = 32'd10898
; 
32'd128795: dataIn1 = 32'd10899
; 
32'd128796: dataIn1 = 32'd857
; 
32'd128797: dataIn1 = 32'd861
; 
32'd128798: dataIn1 = 32'd1591
; 
32'd128799: dataIn1 = 32'd10420
; 
32'd128800: dataIn1 = 32'd10421
; 
32'd128801: dataIn1 = 32'd10890
; 
32'd128802: dataIn1 = 32'd10891
; 
32'd128803: dataIn1 = 32'd862
; 
32'd128804: dataIn1 = 32'd863
; 
32'd128805: dataIn1 = 32'd1592
; 
32'd128806: dataIn1 = 32'd10416
; 
32'd128807: dataIn1 = 32'd10417
; 
32'd128808: dataIn1 = 32'd10886
; 
32'd128809: dataIn1 = 32'd10887
; 
32'd128810: dataIn1 = 32'd861
; 
32'd128811: dataIn1 = 32'd862
; 
32'd128812: dataIn1 = 32'd1593
; 
32'd128813: dataIn1 = 32'd10418
; 
32'd128814: dataIn1 = 32'd10419
; 
32'd128815: dataIn1 = 32'd10888
; 
32'd128816: dataIn1 = 32'd10889
; 
32'd128817: dataIn1 = 32'd426
; 
32'd128818: dataIn1 = 32'd864
; 
32'd128819: dataIn1 = 32'd1594
; 
32'd128820: dataIn1 = 32'd1914
; 
32'd128821: dataIn1 = 32'd10417
; 
32'd128822: dataIn1 = 32'd10418
; 
32'd128823: dataIn1 = 32'd226
; 
32'd128824: dataIn1 = 32'd864
; 
32'd128825: dataIn1 = 32'd1595
; 
32'd128826: dataIn1 = 32'd1913
; 
32'd128827: dataIn1 = 32'd10419
; 
32'd128828: dataIn1 = 32'd10420
; 
32'd128829: dataIn1 = 32'd863
; 
32'd128830: dataIn1 = 32'd865
; 
32'd128831: dataIn1 = 32'd1596
; 
32'd128832: dataIn1 = 32'd10414
; 
32'd128833: dataIn1 = 32'd10415
; 
32'd128834: dataIn1 = 32'd10884
; 
32'd128835: dataIn1 = 32'd10885
; 
32'd128836: dataIn1 = 32'd426
; 
32'd128837: dataIn1 = 32'd866
; 
32'd128838: dataIn1 = 32'd1597
; 
32'd128839: dataIn1 = 32'd1916
; 
32'd128840: dataIn1 = 32'd10415
; 
32'd128841: dataIn1 = 32'd10416
; 
32'd128842: dataIn1 = 32'd228
; 
32'd128843: dataIn1 = 32'd866
; 
32'd128844: dataIn1 = 32'd1598
; 
32'd128845: dataIn1 = 32'd1915
; 
32'd128846: dataIn1 = 32'd10413
; 
32'd128847: dataIn1 = 32'd10414
; 
32'd128848: dataIn1 = 32'd867
; 
32'd128849: dataIn1 = 32'd868
; 
32'd128850: dataIn1 = 32'd1599
; 
32'd128851: dataIn1 = 32'd10400
; 
32'd128852: dataIn1 = 32'd10401
; 
32'd128853: dataIn1 = 32'd10870
; 
32'd128854: dataIn1 = 32'd10871
; 
32'd128855: dataIn1 = 32'd867
; 
32'd128856: dataIn1 = 32'd869
; 
32'd128857: dataIn1 = 32'd1600
; 
32'd128858: dataIn1 = 32'd10402
; 
32'd128859: dataIn1 = 32'd10403
; 
32'd128860: dataIn1 = 32'd10872
; 
32'd128861: dataIn1 = 32'd10873
; 
32'd128862: dataIn1 = 32'd229
; 
32'd128863: dataIn1 = 32'd870
; 
32'd128864: dataIn1 = 32'd1601
; 
32'd128865: dataIn1 = 32'd1918
; 
32'd128866: dataIn1 = 32'd10403
; 
32'd128867: dataIn1 = 32'd10404
; 
32'd128868: dataIn1 = 32'd427
; 
32'd128869: dataIn1 = 32'd870
; 
32'd128870: dataIn1 = 32'd1602
; 
32'd128871: dataIn1 = 32'd1917
; 
32'd128872: dataIn1 = 32'd10401
; 
32'd128873: dataIn1 = 32'd10402
; 
32'd128874: dataIn1 = 32'd868
; 
32'd128875: dataIn1 = 32'd872
; 
32'd128876: dataIn1 = 32'd1603
; 
32'd128877: dataIn1 = 32'd10398
; 
32'd128878: dataIn1 = 32'd10399
; 
32'd128879: dataIn1 = 32'd10868
; 
32'd128880: dataIn1 = 32'd10869
; 
32'd128881: dataIn1 = 32'd427
; 
32'd128882: dataIn1 = 32'd871
; 
32'd128883: dataIn1 = 32'd1604
; 
32'd128884: dataIn1 = 32'd1920
; 
32'd128885: dataIn1 = 32'd10399
; 
32'd128886: dataIn1 = 32'd10400
; 
32'd128887: dataIn1 = 32'd231
; 
32'd128888: dataIn1 = 32'd871
; 
32'd128889: dataIn1 = 32'd1605
; 
32'd128890: dataIn1 = 32'd1919
; 
32'd128891: dataIn1 = 32'd10397
; 
32'd128892: dataIn1 = 32'd10398
; 
32'd128893: dataIn1 = 32'd873
; 
32'd128894: dataIn1 = 32'd874
; 
32'd128895: dataIn1 = 32'd1606
; 
32'd128896: dataIn1 = 32'd10408
; 
32'd128897: dataIn1 = 32'd10409
; 
32'd128898: dataIn1 = 32'd10878
; 
32'd128899: dataIn1 = 32'd10879
; 
32'd128900: dataIn1 = 32'd873
; 
32'd128901: dataIn1 = 32'd876
; 
32'd128902: dataIn1 = 32'd1607
; 
32'd128903: dataIn1 = 32'd10406
; 
32'd128904: dataIn1 = 32'd10407
; 
32'd128905: dataIn1 = 32'd10876
; 
32'd128906: dataIn1 = 32'd10877
; 
32'd128907: dataIn1 = 32'd229
; 
32'd128908: dataIn1 = 32'd875
; 
32'd128909: dataIn1 = 32'd1608
; 
32'd128910: dataIn1 = 32'd1922
; 
32'd128911: dataIn1 = 32'd10405
; 
32'd128912: dataIn1 = 32'd10406
; 
32'd128913: dataIn1 = 32'd428
; 
32'd128914: dataIn1 = 32'd875
; 
32'd128915: dataIn1 = 32'd1609
; 
32'd128916: dataIn1 = 32'd1921
; 
32'd128917: dataIn1 = 32'd10407
; 
32'd128918: dataIn1 = 32'd10408
; 
32'd128919: dataIn1 = 32'd874
; 
32'd128920: dataIn1 = 32'd878
; 
32'd128921: dataIn1 = 32'd1610
; 
32'd128922: dataIn1 = 32'd10410
; 
32'd128923: dataIn1 = 32'd10411
; 
32'd128924: dataIn1 = 32'd10880
; 
32'd128925: dataIn1 = 32'd10881
; 
32'd128926: dataIn1 = 32'd228
; 
32'd128927: dataIn1 = 32'd877
; 
32'd128928: dataIn1 = 32'd1611
; 
32'd128929: dataIn1 = 32'd1924
; 
32'd128930: dataIn1 = 32'd10411
; 
32'd128931: dataIn1 = 32'd10412
; 
32'd128932: dataIn1 = 32'd428
; 
32'd128933: dataIn1 = 32'd877
; 
32'd128934: dataIn1 = 32'd1612
; 
32'd128935: dataIn1 = 32'd1923
; 
32'd128936: dataIn1 = 32'd10409
; 
32'd128937: dataIn1 = 32'd10410
; 
32'd128938: dataIn1 = 32'd865
; 
32'd128939: dataIn1 = 32'd878
; 
32'd128940: dataIn1 = 32'd1613
; 
32'd128941: dataIn1 = 32'd10412
; 
32'd128942: dataIn1 = 32'd10413
; 
32'd128943: dataIn1 = 32'd10882
; 
32'd128944: dataIn1 = 32'd10883
; 
32'd128945: dataIn1 = 32'd869
; 
32'd128946: dataIn1 = 32'd876
; 
32'd128947: dataIn1 = 32'd1614
; 
32'd128948: dataIn1 = 32'd10404
; 
32'd128949: dataIn1 = 32'd10405
; 
32'd128950: dataIn1 = 32'd10874
; 
32'd128951: dataIn1 = 32'd10875
; 
32'd128952: dataIn1 = 32'd879
; 
32'd128953: dataIn1 = 32'd880
; 
32'd128954: dataIn1 = 32'd1615
; 
32'd128955: dataIn1 = 32'd10392
; 
32'd128956: dataIn1 = 32'd10393
; 
32'd128957: dataIn1 = 32'd10862
; 
32'd128958: dataIn1 = 32'd10863
; 
32'd128959: dataIn1 = 32'd879
; 
32'd128960: dataIn1 = 32'd881
; 
32'd128961: dataIn1 = 32'd1616
; 
32'd128962: dataIn1 = 32'd10390
; 
32'd128963: dataIn1 = 32'd10391
; 
32'd128964: dataIn1 = 32'd10860
; 
32'd128965: dataIn1 = 32'd10861
; 
32'd128966: dataIn1 = 32'd429
; 
32'd128967: dataIn1 = 32'd882
; 
32'd128968: dataIn1 = 32'd1617
; 
32'd128969: dataIn1 = 32'd1926
; 
32'd128970: dataIn1 = 32'd10391
; 
32'd128971: dataIn1 = 32'd10392
; 
32'd128972: dataIn1 = 32'd232
; 
32'd128973: dataIn1 = 32'd882
; 
32'd128974: dataIn1 = 32'd1618
; 
32'd128975: dataIn1 = 32'd1925
; 
32'd128976: dataIn1 = 32'd10389
; 
32'd128977: dataIn1 = 32'd10390
; 
32'd128978: dataIn1 = 32'd880
; 
32'd128979: dataIn1 = 32'd883
; 
32'd128980: dataIn1 = 32'd1619
; 
32'd128981: dataIn1 = 32'd10394
; 
32'd128982: dataIn1 = 32'd10395
; 
32'd128983: dataIn1 = 32'd10864
; 
32'd128984: dataIn1 = 32'd10865
; 
32'd128985: dataIn1 = 32'd429
; 
32'd128986: dataIn1 = 32'd884
; 
32'd128987: dataIn1 = 32'd1620
; 
32'd128988: dataIn1 = 32'd1928
; 
32'd128989: dataIn1 = 32'd10393
; 
32'd128990: dataIn1 = 32'd10394
; 
32'd128991: dataIn1 = 32'd231
; 
32'd128992: dataIn1 = 32'd884
; 
32'd128993: dataIn1 = 32'd1621
; 
32'd128994: dataIn1 = 32'd1927
; 
32'd128995: dataIn1 = 32'd10395
; 
32'd128996: dataIn1 = 32'd10396
; 
32'd128997: dataIn1 = 32'd872
; 
32'd128998: dataIn1 = 32'd883
; 
32'd128999: dataIn1 = 32'd1622
; 
32'd129000: dataIn1 = 32'd10396
; 
32'd129001: dataIn1 = 32'd10397
; 
32'd129002: dataIn1 = 32'd10866
; 
32'd129003: dataIn1 = 32'd10867
; 
32'd129004: dataIn1 = 32'd881
; 
32'd129005: dataIn1 = 32'd885
; 
32'd129006: dataIn1 = 32'd1623
; 
32'd129007: dataIn1 = 32'd10388
; 
32'd129008: dataIn1 = 32'd10389
; 
32'd129009: dataIn1 = 32'd10858
; 
32'd129010: dataIn1 = 32'd10859
; 
32'd129011: dataIn1 = 32'd886
; 
32'd129012: dataIn1 = 32'd887
; 
32'd129013: dataIn1 = 32'd1624
; 
32'd129014: dataIn1 = 32'd10384
; 
32'd129015: dataIn1 = 32'd10385
; 
32'd129016: dataIn1 = 32'd10854
; 
32'd129017: dataIn1 = 32'd10855
; 
32'd129018: dataIn1 = 32'd885
; 
32'd129019: dataIn1 = 32'd886
; 
32'd129020: dataIn1 = 32'd1625
; 
32'd129021: dataIn1 = 32'd10386
; 
32'd129022: dataIn1 = 32'd10387
; 
32'd129023: dataIn1 = 32'd10856
; 
32'd129024: dataIn1 = 32'd10857
; 
32'd129025: dataIn1 = 32'd430
; 
32'd129026: dataIn1 = 32'd888
; 
32'd129027: dataIn1 = 32'd1626
; 
32'd129028: dataIn1 = 32'd1930
; 
32'd129029: dataIn1 = 32'd10385
; 
32'd129030: dataIn1 = 32'd10386
; 
32'd129031: dataIn1 = 32'd232
; 
32'd129032: dataIn1 = 32'd888
; 
32'd129033: dataIn1 = 32'd1627
; 
32'd129034: dataIn1 = 32'd1929
; 
32'd129035: dataIn1 = 32'd10387
; 
32'd129036: dataIn1 = 32'd10388
; 
32'd129037: dataIn1 = 32'd887
; 
32'd129038: dataIn1 = 32'd889
; 
32'd129039: dataIn1 = 32'd1628
; 
32'd129040: dataIn1 = 32'd10382
; 
32'd129041: dataIn1 = 32'd10383
; 
32'd129042: dataIn1 = 32'd10852
; 
32'd129043: dataIn1 = 32'd10853
; 
32'd129044: dataIn1 = 32'd430
; 
32'd129045: dataIn1 = 32'd890
; 
32'd129046: dataIn1 = 32'd1629
; 
32'd129047: dataIn1 = 32'd1932
; 
32'd129048: dataIn1 = 32'd10383
; 
32'd129049: dataIn1 = 32'd10384
; 
32'd129050: dataIn1 = 32'd234
; 
32'd129051: dataIn1 = 32'd890
; 
32'd129052: dataIn1 = 32'd1630
; 
32'd129053: dataIn1 = 32'd1931
; 
32'd129054: dataIn1 = 32'd10381
; 
32'd129055: dataIn1 = 32'd10382
; 
32'd129056: dataIn1 = 32'd891
; 
32'd129057: dataIn1 = 32'd892
; 
32'd129058: dataIn1 = 32'd1631
; 
32'd129059: dataIn1 = 32'd10368
; 
32'd129060: dataIn1 = 32'd10369
; 
32'd129061: dataIn1 = 32'd10838
; 
32'd129062: dataIn1 = 32'd10839
; 
32'd129063: dataIn1 = 32'd891
; 
32'd129064: dataIn1 = 32'd893
; 
32'd129065: dataIn1 = 32'd1632
; 
32'd129066: dataIn1 = 32'd10370
; 
32'd129067: dataIn1 = 32'd10371
; 
32'd129068: dataIn1 = 32'd10840
; 
32'd129069: dataIn1 = 32'd10841
; 
32'd129070: dataIn1 = 32'd235
; 
32'd129071: dataIn1 = 32'd894
; 
32'd129072: dataIn1 = 32'd1633
; 
32'd129073: dataIn1 = 32'd1934
; 
32'd129074: dataIn1 = 32'd10371
; 
32'd129075: dataIn1 = 32'd10372
; 
32'd129076: dataIn1 = 32'd431
; 
32'd129077: dataIn1 = 32'd894
; 
32'd129078: dataIn1 = 32'd1634
; 
32'd129079: dataIn1 = 32'd1933
; 
32'd129080: dataIn1 = 32'd10369
; 
32'd129081: dataIn1 = 32'd10370
; 
32'd129082: dataIn1 = 32'd892
; 
32'd129083: dataIn1 = 32'd896
; 
32'd129084: dataIn1 = 32'd1635
; 
32'd129085: dataIn1 = 32'd10366
; 
32'd129086: dataIn1 = 32'd10367
; 
32'd129087: dataIn1 = 32'd10836
; 
32'd129088: dataIn1 = 32'd10837
; 
32'd129089: dataIn1 = 32'd431
; 
32'd129090: dataIn1 = 32'd895
; 
32'd129091: dataIn1 = 32'd1636
; 
32'd129092: dataIn1 = 32'd1936
; 
32'd129093: dataIn1 = 32'd10367
; 
32'd129094: dataIn1 = 32'd10368
; 
32'd129095: dataIn1 = 32'd237
; 
32'd129096: dataIn1 = 32'd895
; 
32'd129097: dataIn1 = 32'd1637
; 
32'd129098: dataIn1 = 32'd1935
; 
32'd129099: dataIn1 = 32'd10365
; 
32'd129100: dataIn1 = 32'd10366
; 
32'd129101: dataIn1 = 32'd897
; 
32'd129102: dataIn1 = 32'd898
; 
32'd129103: dataIn1 = 32'd1638
; 
32'd129104: dataIn1 = 32'd10376
; 
32'd129105: dataIn1 = 32'd10377
; 
32'd129106: dataIn1 = 32'd10846
; 
32'd129107: dataIn1 = 32'd10847
; 
32'd129108: dataIn1 = 32'd897
; 
32'd129109: dataIn1 = 32'd900
; 
32'd129110: dataIn1 = 32'd1639
; 
32'd129111: dataIn1 = 32'd10374
; 
32'd129112: dataIn1 = 32'd10375
; 
32'd129113: dataIn1 = 32'd10844
; 
32'd129114: dataIn1 = 32'd10845
; 
32'd129115: dataIn1 = 32'd235
; 
32'd129116: dataIn1 = 32'd899
; 
32'd129117: dataIn1 = 32'd1640
; 
32'd129118: dataIn1 = 32'd1938
; 
32'd129119: dataIn1 = 32'd10373
; 
32'd129120: dataIn1 = 32'd10374
; 
32'd129121: dataIn1 = 32'd432
; 
32'd129122: dataIn1 = 32'd899
; 
32'd129123: dataIn1 = 32'd1641
; 
32'd129124: dataIn1 = 32'd1937
; 
32'd129125: dataIn1 = 32'd10375
; 
32'd129126: dataIn1 = 32'd10376
; 
32'd129127: dataIn1 = 32'd898
; 
32'd129128: dataIn1 = 32'd902
; 
32'd129129: dataIn1 = 32'd1642
; 
32'd129130: dataIn1 = 32'd10378
; 
32'd129131: dataIn1 = 32'd10379
; 
32'd129132: dataIn1 = 32'd10848
; 
32'd129133: dataIn1 = 32'd10849
; 
32'd129134: dataIn1 = 32'd234
; 
32'd129135: dataIn1 = 32'd901
; 
32'd129136: dataIn1 = 32'd1643
; 
32'd129137: dataIn1 = 32'd1940
; 
32'd129138: dataIn1 = 32'd10379
; 
32'd129139: dataIn1 = 32'd10380
; 
32'd129140: dataIn1 = 32'd432
; 
32'd129141: dataIn1 = 32'd901
; 
32'd129142: dataIn1 = 32'd1644
; 
32'd129143: dataIn1 = 32'd1939
; 
32'd129144: dataIn1 = 32'd10377
; 
32'd129145: dataIn1 = 32'd10378
; 
32'd129146: dataIn1 = 32'd889
; 
32'd129147: dataIn1 = 32'd902
; 
32'd129148: dataIn1 = 32'd1645
; 
32'd129149: dataIn1 = 32'd10380
; 
32'd129150: dataIn1 = 32'd10381
; 
32'd129151: dataIn1 = 32'd10850
; 
32'd129152: dataIn1 = 32'd10851
; 
32'd129153: dataIn1 = 32'd893
; 
32'd129154: dataIn1 = 32'd900
; 
32'd129155: dataIn1 = 32'd1646
; 
32'd129156: dataIn1 = 32'd10372
; 
32'd129157: dataIn1 = 32'd10373
; 
32'd129158: dataIn1 = 32'd10842
; 
32'd129159: dataIn1 = 32'd10843
; 
32'd129160: dataIn1 = 32'd903
; 
32'd129161: dataIn1 = 32'd904
; 
32'd129162: dataIn1 = 32'd1647
; 
32'd129163: dataIn1 = 32'd10360
; 
32'd129164: dataIn1 = 32'd10361
; 
32'd129165: dataIn1 = 32'd10830
; 
32'd129166: dataIn1 = 32'd10831
; 
32'd129167: dataIn1 = 32'd903
; 
32'd129168: dataIn1 = 32'd905
; 
32'd129169: dataIn1 = 32'd1648
; 
32'd129170: dataIn1 = 32'd10358
; 
32'd129171: dataIn1 = 32'd10359
; 
32'd129172: dataIn1 = 32'd10828
; 
32'd129173: dataIn1 = 32'd10829
; 
32'd129174: dataIn1 = 32'd433
; 
32'd129175: dataIn1 = 32'd906
; 
32'd129176: dataIn1 = 32'd1649
; 
32'd129177: dataIn1 = 32'd1942
; 
32'd129178: dataIn1 = 32'd10359
; 
32'd129179: dataIn1 = 32'd10360
; 
32'd129180: dataIn1 = 32'd238
; 
32'd129181: dataIn1 = 32'd906
; 
32'd129182: dataIn1 = 32'd1650
; 
32'd129183: dataIn1 = 32'd1941
; 
32'd129184: dataIn1 = 32'd10357
; 
32'd129185: dataIn1 = 32'd10358
; 
32'd129186: dataIn1 = 32'd904
; 
32'd129187: dataIn1 = 32'd907
; 
32'd129188: dataIn1 = 32'd1651
; 
32'd129189: dataIn1 = 32'd10362
; 
32'd129190: dataIn1 = 32'd10363
; 
32'd129191: dataIn1 = 32'd10832
; 
32'd129192: dataIn1 = 32'd10833
; 
32'd129193: dataIn1 = 32'd433
; 
32'd129194: dataIn1 = 32'd908
; 
32'd129195: dataIn1 = 32'd1652
; 
32'd129196: dataIn1 = 32'd1944
; 
32'd129197: dataIn1 = 32'd10361
; 
32'd129198: dataIn1 = 32'd10362
; 
32'd129199: dataIn1 = 32'd237
; 
32'd129200: dataIn1 = 32'd908
; 
32'd129201: dataIn1 = 32'd1653
; 
32'd129202: dataIn1 = 32'd1943
; 
32'd129203: dataIn1 = 32'd10363
; 
32'd129204: dataIn1 = 32'd10364
; 
32'd129205: dataIn1 = 32'd896
; 
32'd129206: dataIn1 = 32'd907
; 
32'd129207: dataIn1 = 32'd1654
; 
32'd129208: dataIn1 = 32'd10364
; 
32'd129209: dataIn1 = 32'd10365
; 
32'd129210: dataIn1 = 32'd10834
; 
32'd129211: dataIn1 = 32'd10835
; 
32'd129212: dataIn1 = 32'd905
; 
32'd129213: dataIn1 = 32'd909
; 
32'd129214: dataIn1 = 32'd1655
; 
32'd129215: dataIn1 = 32'd10356
; 
32'd129216: dataIn1 = 32'd10357
; 
32'd129217: dataIn1 = 32'd10826
; 
32'd129218: dataIn1 = 32'd10827
; 
32'd129219: dataIn1 = 32'd910
; 
32'd129220: dataIn1 = 32'd911
; 
32'd129221: dataIn1 = 32'd1656
; 
32'd129222: dataIn1 = 32'd10352
; 
32'd129223: dataIn1 = 32'd10353
; 
32'd129224: dataIn1 = 32'd10822
; 
32'd129225: dataIn1 = 32'd10823
; 
32'd129226: dataIn1 = 32'd909
; 
32'd129227: dataIn1 = 32'd910
; 
32'd129228: dataIn1 = 32'd1657
; 
32'd129229: dataIn1 = 32'd10354
; 
32'd129230: dataIn1 = 32'd10355
; 
32'd129231: dataIn1 = 32'd10824
; 
32'd129232: dataIn1 = 32'd10825
; 
32'd129233: dataIn1 = 32'd434
; 
32'd129234: dataIn1 = 32'd912
; 
32'd129235: dataIn1 = 32'd1658
; 
32'd129236: dataIn1 = 32'd1946
; 
32'd129237: dataIn1 = 32'd10353
; 
32'd129238: dataIn1 = 32'd10354
; 
32'd129239: dataIn1 = 32'd238
; 
32'd129240: dataIn1 = 32'd912
; 
32'd129241: dataIn1 = 32'd1659
; 
32'd129242: dataIn1 = 32'd1945
; 
32'd129243: dataIn1 = 32'd10355
; 
32'd129244: dataIn1 = 32'd10356
; 
32'd129245: dataIn1 = 32'd911
; 
32'd129246: dataIn1 = 32'd913
; 
32'd129247: dataIn1 = 32'd1660
; 
32'd129248: dataIn1 = 32'd10350
; 
32'd129249: dataIn1 = 32'd10351
; 
32'd129250: dataIn1 = 32'd10820
; 
32'd129251: dataIn1 = 32'd10821
; 
32'd129252: dataIn1 = 32'd434
; 
32'd129253: dataIn1 = 32'd914
; 
32'd129254: dataIn1 = 32'd1661
; 
32'd129255: dataIn1 = 32'd1948
; 
32'd129256: dataIn1 = 32'd10351
; 
32'd129257: dataIn1 = 32'd10352
; 
32'd129258: dataIn1 = 32'd240
; 
32'd129259: dataIn1 = 32'd914
; 
32'd129260: dataIn1 = 32'd1662
; 
32'd129261: dataIn1 = 32'd1947
; 
32'd129262: dataIn1 = 32'd10349
; 
32'd129263: dataIn1 = 32'd10350
; 
32'd129264: dataIn1 = 32'd915
; 
32'd129265: dataIn1 = 32'd916
; 
32'd129266: dataIn1 = 32'd1663
; 
32'd129267: dataIn1 = 32'd10336
; 
32'd129268: dataIn1 = 32'd10337
; 
32'd129269: dataIn1 = 32'd10806
; 
32'd129270: dataIn1 = 32'd10807
; 
32'd129271: dataIn1 = 32'd915
; 
32'd129272: dataIn1 = 32'd917
; 
32'd129273: dataIn1 = 32'd1664
; 
32'd129274: dataIn1 = 32'd10338
; 
32'd129275: dataIn1 = 32'd10339
; 
32'd129276: dataIn1 = 32'd10808
; 
32'd129277: dataIn1 = 32'd10809
; 
32'd129278: dataIn1 = 32'd241
; 
32'd129279: dataIn1 = 32'd918
; 
32'd129280: dataIn1 = 32'd1665
; 
32'd129281: dataIn1 = 32'd1950
; 
32'd129282: dataIn1 = 32'd10339
; 
32'd129283: dataIn1 = 32'd10340
; 
32'd129284: dataIn1 = 32'd435
; 
32'd129285: dataIn1 = 32'd918
; 
32'd129286: dataIn1 = 32'd1666
; 
32'd129287: dataIn1 = 32'd1949
; 
32'd129288: dataIn1 = 32'd10337
; 
32'd129289: dataIn1 = 32'd10338
; 
32'd129290: dataIn1 = 32'd916
; 
32'd129291: dataIn1 = 32'd920
; 
32'd129292: dataIn1 = 32'd1667
; 
32'd129293: dataIn1 = 32'd10334
; 
32'd129294: dataIn1 = 32'd10335
; 
32'd129295: dataIn1 = 32'd10804
; 
32'd129296: dataIn1 = 32'd10805
; 
32'd129297: dataIn1 = 32'd435
; 
32'd129298: dataIn1 = 32'd919
; 
32'd129299: dataIn1 = 32'd1668
; 
32'd129300: dataIn1 = 32'd1952
; 
32'd129301: dataIn1 = 32'd10335
; 
32'd129302: dataIn1 = 32'd10336
; 
32'd129303: dataIn1 = 32'd243
; 
32'd129304: dataIn1 = 32'd919
; 
32'd129305: dataIn1 = 32'd1669
; 
32'd129306: dataIn1 = 32'd1951
; 
32'd129307: dataIn1 = 32'd10333
; 
32'd129308: dataIn1 = 32'd10334
; 
32'd129309: dataIn1 = 32'd921
; 
32'd129310: dataIn1 = 32'd922
; 
32'd129311: dataIn1 = 32'd1670
; 
32'd129312: dataIn1 = 32'd10344
; 
32'd129313: dataIn1 = 32'd10345
; 
32'd129314: dataIn1 = 32'd10814
; 
32'd129315: dataIn1 = 32'd10815
; 
32'd129316: dataIn1 = 32'd921
; 
32'd129317: dataIn1 = 32'd924
; 
32'd129318: dataIn1 = 32'd1671
; 
32'd129319: dataIn1 = 32'd10342
; 
32'd129320: dataIn1 = 32'd10343
; 
32'd129321: dataIn1 = 32'd10812
; 
32'd129322: dataIn1 = 32'd10813
; 
32'd129323: dataIn1 = 32'd241
; 
32'd129324: dataIn1 = 32'd923
; 
32'd129325: dataIn1 = 32'd1672
; 
32'd129326: dataIn1 = 32'd1954
; 
32'd129327: dataIn1 = 32'd10341
; 
32'd129328: dataIn1 = 32'd10342
; 
32'd129329: dataIn1 = 32'd436
; 
32'd129330: dataIn1 = 32'd923
; 
32'd129331: dataIn1 = 32'd1673
; 
32'd129332: dataIn1 = 32'd1953
; 
32'd129333: dataIn1 = 32'd10343
; 
32'd129334: dataIn1 = 32'd10344
; 
32'd129335: dataIn1 = 32'd922
; 
32'd129336: dataIn1 = 32'd926
; 
32'd129337: dataIn1 = 32'd1674
; 
32'd129338: dataIn1 = 32'd10346
; 
32'd129339: dataIn1 = 32'd10347
; 
32'd129340: dataIn1 = 32'd10816
; 
32'd129341: dataIn1 = 32'd10817
; 
32'd129342: dataIn1 = 32'd240
; 
32'd129343: dataIn1 = 32'd925
; 
32'd129344: dataIn1 = 32'd1675
; 
32'd129345: dataIn1 = 32'd1956
; 
32'd129346: dataIn1 = 32'd10347
; 
32'd129347: dataIn1 = 32'd10348
; 
32'd129348: dataIn1 = 32'd436
; 
32'd129349: dataIn1 = 32'd925
; 
32'd129350: dataIn1 = 32'd1676
; 
32'd129351: dataIn1 = 32'd1955
; 
32'd129352: dataIn1 = 32'd10345
; 
32'd129353: dataIn1 = 32'd10346
; 
32'd129354: dataIn1 = 32'd913
; 
32'd129355: dataIn1 = 32'd926
; 
32'd129356: dataIn1 = 32'd1677
; 
32'd129357: dataIn1 = 32'd10348
; 
32'd129358: dataIn1 = 32'd10349
; 
32'd129359: dataIn1 = 32'd10818
; 
32'd129360: dataIn1 = 32'd10819
; 
32'd129361: dataIn1 = 32'd917
; 
32'd129362: dataIn1 = 32'd924
; 
32'd129363: dataIn1 = 32'd1678
; 
32'd129364: dataIn1 = 32'd10340
; 
32'd129365: dataIn1 = 32'd10341
; 
32'd129366: dataIn1 = 32'd10810
; 
32'd129367: dataIn1 = 32'd10811
; 
32'd129368: dataIn1 = 32'd927
; 
32'd129369: dataIn1 = 32'd928
; 
32'd129370: dataIn1 = 32'd1679
; 
32'd129371: dataIn1 = 32'd10328
; 
32'd129372: dataIn1 = 32'd10329
; 
32'd129373: dataIn1 = 32'd10798
; 
32'd129374: dataIn1 = 32'd10799
; 
32'd129375: dataIn1 = 32'd927
; 
32'd129376: dataIn1 = 32'd929
; 
32'd129377: dataIn1 = 32'd1680
; 
32'd129378: dataIn1 = 32'd10326
; 
32'd129379: dataIn1 = 32'd10327
; 
32'd129380: dataIn1 = 32'd10796
; 
32'd129381: dataIn1 = 32'd10797
; 
32'd129382: dataIn1 = 32'd437
; 
32'd129383: dataIn1 = 32'd930
; 
32'd129384: dataIn1 = 32'd1681
; 
32'd129385: dataIn1 = 32'd1958
; 
32'd129386: dataIn1 = 32'd10327
; 
32'd129387: dataIn1 = 32'd10328
; 
32'd129388: dataIn1 = 32'd244
; 
32'd129389: dataIn1 = 32'd930
; 
32'd129390: dataIn1 = 32'd1682
; 
32'd129391: dataIn1 = 32'd1957
; 
32'd129392: dataIn1 = 32'd10325
; 
32'd129393: dataIn1 = 32'd10326
; 
32'd129394: dataIn1 = 32'd928
; 
32'd129395: dataIn1 = 32'd931
; 
32'd129396: dataIn1 = 32'd1683
; 
32'd129397: dataIn1 = 32'd10330
; 
32'd129398: dataIn1 = 32'd10331
; 
32'd129399: dataIn1 = 32'd10800
; 
32'd129400: dataIn1 = 32'd10801
; 
32'd129401: dataIn1 = 32'd437
; 
32'd129402: dataIn1 = 32'd932
; 
32'd129403: dataIn1 = 32'd1684
; 
32'd129404: dataIn1 = 32'd1960
; 
32'd129405: dataIn1 = 32'd10329
; 
32'd129406: dataIn1 = 32'd10330
; 
32'd129407: dataIn1 = 32'd243
; 
32'd129408: dataIn1 = 32'd932
; 
32'd129409: dataIn1 = 32'd1685
; 
32'd129410: dataIn1 = 32'd1959
; 
32'd129411: dataIn1 = 32'd10331
; 
32'd129412: dataIn1 = 32'd10332
; 
32'd129413: dataIn1 = 32'd920
; 
32'd129414: dataIn1 = 32'd931
; 
32'd129415: dataIn1 = 32'd1686
; 
32'd129416: dataIn1 = 32'd10332
; 
32'd129417: dataIn1 = 32'd10333
; 
32'd129418: dataIn1 = 32'd10802
; 
32'd129419: dataIn1 = 32'd10803
; 
32'd129420: dataIn1 = 32'd929
; 
32'd129421: dataIn1 = 32'd933
; 
32'd129422: dataIn1 = 32'd1687
; 
32'd129423: dataIn1 = 32'd10324
; 
32'd129424: dataIn1 = 32'd10325
; 
32'd129425: dataIn1 = 32'd10794
; 
32'd129426: dataIn1 = 32'd10795
; 
32'd129427: dataIn1 = 32'd934
; 
32'd129428: dataIn1 = 32'd935
; 
32'd129429: dataIn1 = 32'd1688
; 
32'd129430: dataIn1 = 32'd10320
; 
32'd129431: dataIn1 = 32'd10321
; 
32'd129432: dataIn1 = 32'd10790
; 
32'd129433: dataIn1 = 32'd10791
; 
32'd129434: dataIn1 = 32'd933
; 
32'd129435: dataIn1 = 32'd934
; 
32'd129436: dataIn1 = 32'd1689
; 
32'd129437: dataIn1 = 32'd10322
; 
32'd129438: dataIn1 = 32'd10323
; 
32'd129439: dataIn1 = 32'd10792
; 
32'd129440: dataIn1 = 32'd10793
; 
32'd129441: dataIn1 = 32'd438
; 
32'd129442: dataIn1 = 32'd936
; 
32'd129443: dataIn1 = 32'd1690
; 
32'd129444: dataIn1 = 32'd1962
; 
32'd129445: dataIn1 = 32'd10321
; 
32'd129446: dataIn1 = 32'd10322
; 
32'd129447: dataIn1 = 32'd244
; 
32'd129448: dataIn1 = 32'd936
; 
32'd129449: dataIn1 = 32'd1691
; 
32'd129450: dataIn1 = 32'd1961
; 
32'd129451: dataIn1 = 32'd10323
; 
32'd129452: dataIn1 = 32'd10324
; 
32'd129453: dataIn1 = 32'd935
; 
32'd129454: dataIn1 = 32'd937
; 
32'd129455: dataIn1 = 32'd1692
; 
32'd129456: dataIn1 = 32'd10318
; 
32'd129457: dataIn1 = 32'd10319
; 
32'd129458: dataIn1 = 32'd10788
; 
32'd129459: dataIn1 = 32'd10789
; 
32'd129460: dataIn1 = 32'd438
; 
32'd129461: dataIn1 = 32'd938
; 
32'd129462: dataIn1 = 32'd1693
; 
32'd129463: dataIn1 = 32'd1964
; 
32'd129464: dataIn1 = 32'd10319
; 
32'd129465: dataIn1 = 32'd10320
; 
32'd129466: dataIn1 = 32'd246
; 
32'd129467: dataIn1 = 32'd938
; 
32'd129468: dataIn1 = 32'd1694
; 
32'd129469: dataIn1 = 32'd1963
; 
32'd129470: dataIn1 = 32'd10317
; 
32'd129471: dataIn1 = 32'd10318
; 
32'd129472: dataIn1 = 32'd939
; 
32'd129473: dataIn1 = 32'd940
; 
32'd129474: dataIn1 = 32'd1695
; 
32'd129475: dataIn1 = 32'd10304
; 
32'd129476: dataIn1 = 32'd10305
; 
32'd129477: dataIn1 = 32'd10774
; 
32'd129478: dataIn1 = 32'd10775
; 
32'd129479: dataIn1 = 32'd939
; 
32'd129480: dataIn1 = 32'd941
; 
32'd129481: dataIn1 = 32'd1696
; 
32'd129482: dataIn1 = 32'd10306
; 
32'd129483: dataIn1 = 32'd10307
; 
32'd129484: dataIn1 = 32'd10308
; 
32'd129485: dataIn1 = 32'd10776
; 
32'd129486: dataIn1 = 32'd10777
; 
32'd129487: dataIn1 = 32'd247
; 
32'd129488: dataIn1 = 32'd942
; 
32'd129489: dataIn1 = 32'd1697
; 
32'd129490: dataIn1 = 32'd1966
; 
32'd129491: dataIn1 = 32'd1970
; 
32'd129492: dataIn1 = 32'd10307
; 
32'd129493: dataIn1 = 32'd439
; 
32'd129494: dataIn1 = 32'd942
; 
32'd129495: dataIn1 = 32'd1698
; 
32'd129496: dataIn1 = 32'd1965
; 
32'd129497: dataIn1 = 32'd1966
; 
32'd129498: dataIn1 = 32'd10305
; 
32'd129499: dataIn1 = 32'd10306
; 
32'd129500: dataIn1 = 32'd940
; 
32'd129501: dataIn1 = 32'd944
; 
32'd129502: dataIn1 = 32'd1699
; 
32'd129503: dataIn1 = 32'd10302
; 
32'd129504: dataIn1 = 32'd10303
; 
32'd129505: dataIn1 = 32'd10772
; 
32'd129506: dataIn1 = 32'd10773
; 
32'd129507: dataIn1 = 32'd439
; 
32'd129508: dataIn1 = 32'd943
; 
32'd129509: dataIn1 = 32'd1700
; 
32'd129510: dataIn1 = 32'd1965
; 
32'd129511: dataIn1 = 32'd1968
; 
32'd129512: dataIn1 = 32'd10303
; 
32'd129513: dataIn1 = 32'd10304
; 
32'd129514: dataIn1 = 32'd249
; 
32'd129515: dataIn1 = 32'd943
; 
32'd129516: dataIn1 = 32'd1701
; 
32'd129517: dataIn1 = 32'd1967
; 
32'd129518: dataIn1 = 32'd1968
; 
32'd129519: dataIn1 = 32'd10301
; 
32'd129520: dataIn1 = 32'd10302
; 
32'd129521: dataIn1 = 32'd945
; 
32'd129522: dataIn1 = 32'd946
; 
32'd129523: dataIn1 = 32'd1702
; 
32'd129524: dataIn1 = 32'd10313
; 
32'd129525: dataIn1 = 32'd10314
; 
32'd129526: dataIn1 = 32'd10782
; 
32'd129527: dataIn1 = 32'd10783
; 
32'd129528: dataIn1 = 32'd945
; 
32'd129529: dataIn1 = 32'd948
; 
32'd129530: dataIn1 = 32'd1703
; 
32'd129531: dataIn1 = 32'd10310
; 
32'd129532: dataIn1 = 32'd10311
; 
32'd129533: dataIn1 = 32'd10780
; 
32'd129534: dataIn1 = 32'd10781
; 
32'd129535: dataIn1 = 32'd247
; 
32'd129536: dataIn1 = 32'd947
; 
32'd129537: dataIn1 = 32'd1704
; 
32'd129538: dataIn1 = 32'd1969
; 
32'd129539: dataIn1 = 32'd1970
; 
32'd129540: dataIn1 = 32'd10308
; 
32'd129541: dataIn1 = 32'd10309
; 
32'd129542: dataIn1 = 32'd10310
; 
32'd129543: dataIn1 = 32'd440
; 
32'd129544: dataIn1 = 32'd947
; 
32'd129545: dataIn1 = 32'd1705
; 
32'd129546: dataIn1 = 32'd1969
; 
32'd129547: dataIn1 = 32'd1971
; 
32'd129548: dataIn1 = 32'd10311
; 
32'd129549: dataIn1 = 32'd10312
; 
32'd129550: dataIn1 = 32'd946
; 
32'd129551: dataIn1 = 32'd950
; 
32'd129552: dataIn1 = 32'd1706
; 
32'd129553: dataIn1 = 32'd10315
; 
32'd129554: dataIn1 = 32'd10316
; 
32'd129555: dataIn1 = 32'd10784
; 
32'd129556: dataIn1 = 32'd10785
; 
32'd129557: dataIn1 = 32'd246
; 
32'd129558: dataIn1 = 32'd949
; 
32'd129559: dataIn1 = 32'd1707
; 
32'd129560: dataIn1 = 32'd1972
; 
32'd129561: dataIn1 = 32'd10314
; 
32'd129562: dataIn1 = 32'd10315
; 
32'd129563: dataIn1 = 32'd440
; 
32'd129564: dataIn1 = 32'd949
; 
32'd129565: dataIn1 = 32'd1708
; 
32'd129566: dataIn1 = 32'd1971
; 
32'd129567: dataIn1 = 32'd1972
; 
32'd129568: dataIn1 = 32'd10312
; 
32'd129569: dataIn1 = 32'd10313
; 
32'd129570: dataIn1 = 32'd937
; 
32'd129571: dataIn1 = 32'd950
; 
32'd129572: dataIn1 = 32'd1709
; 
32'd129573: dataIn1 = 32'd10316
; 
32'd129574: dataIn1 = 32'd10317
; 
32'd129575: dataIn1 = 32'd10786
; 
32'd129576: dataIn1 = 32'd10787
; 
32'd129577: dataIn1 = 32'd941
; 
32'd129578: dataIn1 = 32'd948
; 
32'd129579: dataIn1 = 32'd1710
; 
32'd129580: dataIn1 = 32'd10309
; 
32'd129581: dataIn1 = 32'd10778
; 
32'd129582: dataIn1 = 32'd10779
; 
32'd129583: dataIn1 = 32'd951
; 
32'd129584: dataIn1 = 32'd952
; 
32'd129585: dataIn1 = 32'd1711
; 
32'd129586: dataIn1 = 32'd10296
; 
32'd129587: dataIn1 = 32'd10297
; 
32'd129588: dataIn1 = 32'd10766
; 
32'd129589: dataIn1 = 32'd10767
; 
32'd129590: dataIn1 = 32'd951
; 
32'd129591: dataIn1 = 32'd953
; 
32'd129592: dataIn1 = 32'd1712
; 
32'd129593: dataIn1 = 32'd10294
; 
32'd129594: dataIn1 = 32'd10295
; 
32'd129595: dataIn1 = 32'd10764
; 
32'd129596: dataIn1 = 32'd10765
; 
32'd129597: dataIn1 = 32'd441
; 
32'd129598: dataIn1 = 32'd954
; 
32'd129599: dataIn1 = 32'd1713
; 
32'd129600: dataIn1 = 32'd1974
; 
32'd129601: dataIn1 = 32'd1976
; 
32'd129602: dataIn1 = 32'd10295
; 
32'd129603: dataIn1 = 32'd10296
; 
32'd129604: dataIn1 = 32'd250
; 
32'd129605: dataIn1 = 32'd954
; 
32'd129606: dataIn1 = 32'd1714
; 
32'd129607: dataIn1 = 32'd1973
; 
32'd129608: dataIn1 = 32'd1974
; 
32'd129609: dataIn1 = 32'd10293
; 
32'd129610: dataIn1 = 32'd952
; 
32'd129611: dataIn1 = 32'd955
; 
32'd129612: dataIn1 = 32'd1715
; 
32'd129613: dataIn1 = 32'd10298
; 
32'd129614: dataIn1 = 32'd10299
; 
32'd129615: dataIn1 = 32'd10768
; 
32'd129616: dataIn1 = 32'd10769
; 
32'd129617: dataIn1 = 32'd441
; 
32'd129618: dataIn1 = 32'd956
; 
32'd129619: dataIn1 = 32'd1716
; 
32'd129620: dataIn1 = 32'd1975
; 
32'd129621: dataIn1 = 32'd1976
; 
32'd129622: dataIn1 = 32'd10297
; 
32'd129623: dataIn1 = 32'd10298
; 
32'd129624: dataIn1 = 32'd249
; 
32'd129625: dataIn1 = 32'd956
; 
32'd129626: dataIn1 = 32'd1717
; 
32'd129627: dataIn1 = 32'd1967
; 
32'd129628: dataIn1 = 32'd1975
; 
32'd129629: dataIn1 = 32'd10299
; 
32'd129630: dataIn1 = 32'd10300
; 
32'd129631: dataIn1 = 32'd944
; 
32'd129632: dataIn1 = 32'd955
; 
32'd129633: dataIn1 = 32'd1718
; 
32'd129634: dataIn1 = 32'd10300
; 
32'd129635: dataIn1 = 32'd10301
; 
32'd129636: dataIn1 = 32'd10770
; 
32'd129637: dataIn1 = 32'd10771
; 
32'd129638: dataIn1 = 32'd953
; 
32'd129639: dataIn1 = 32'd957
; 
32'd129640: dataIn1 = 32'd1719
; 
32'd129641: dataIn1 = 32'd10293
; 
32'd129642: dataIn1 = 32'd10294
; 
32'd129643: dataIn1 = 32'd10562
; 
32'd129644: dataIn1 = 32'd10762
; 
32'd129645: dataIn1 = 32'd108
; 
32'd129646: dataIn1 = 32'd274
; 
32'd129647: dataIn1 = 32'd561
; 
32'd129648: dataIn1 = 32'd1720
; 
32'd129649: dataIn1 = 32'd1721
; 
32'd129650: dataIn1 = 32'd5526
; 
32'd129651: dataIn1 = 32'd5527
; 
32'd129652: dataIn1 = 32'd108
; 
32'd129653: dataIn1 = 32'd273
; 
32'd129654: dataIn1 = 32'd561
; 
32'd129655: dataIn1 = 32'd572
; 
32'd129656: dataIn1 = 32'd1278
; 
32'd129657: dataIn1 = 32'd1292
; 
32'd129658: dataIn1 = 32'd1720
; 
32'd129659: dataIn1 = 32'd1721
; 
32'd129660: dataIn1 = 32'd1722
; 
32'd129661: dataIn1 = 32'd108
; 
32'd129662: dataIn1 = 32'd278
; 
32'd129663: dataIn1 = 32'd572
; 
32'd129664: dataIn1 = 32'd1721
; 
32'd129665: dataIn1 = 32'd1722
; 
32'd129666: dataIn1 = 32'd5529
; 
32'd129667: dataIn1 = 32'd5530
; 
32'd129668: dataIn1 = 32'd1723
; 
32'd129669: dataIn1 = 32'd2761
; 
32'd129670: dataIn1 = 32'd2763
; 
32'd129671: dataIn1 = 32'd2765
; 
32'd129672: dataIn1 = 32'd3048
; 
32'd129673: dataIn1 = 32'd3050
; 
32'd129674: dataIn1 = 32'd3053
; 
32'd129675: dataIn1 = 32'd1724
; 
32'd129676: dataIn1 = 32'd2761
; 
32'd129677: dataIn1 = 32'd2762
; 
32'd129678: dataIn1 = 32'd2764
; 
32'd129679: dataIn1 = 32'd3041
; 
32'd129680: dataIn1 = 32'd3042
; 
32'd129681: dataIn1 = 32'd3045
; 
32'd129682: dataIn1 = 32'd1725
; 
32'd129683: dataIn1 = 32'd2767
; 
32'd129684: dataIn1 = 32'd2768
; 
32'd129685: dataIn1 = 32'd2771
; 
32'd129686: dataIn1 = 32'd3049
; 
32'd129687: dataIn1 = 32'd3050
; 
32'd129688: dataIn1 = 32'd3054
; 
32'd129689: dataIn1 = 32'd1726
; 
32'd129690: dataIn1 = 32'd2766
; 
32'd129691: dataIn1 = 32'd2767
; 
32'd129692: dataIn1 = 32'd2769
; 
32'd129693: dataIn1 = 32'd2770
; 
32'd129694: dataIn1 = 32'd3868
; 
32'd129695: dataIn1 = 32'd3869
; 
32'd129696: dataIn1 = 32'd1727
; 
32'd129697: dataIn1 = 32'd2773
; 
32'd129698: dataIn1 = 32'd2774
; 
32'd129699: dataIn1 = 32'd2776
; 
32'd129700: dataIn1 = 32'd3063
; 
32'd129701: dataIn1 = 32'd3064
; 
32'd129702: dataIn1 = 32'd3068
; 
32'd129703: dataIn1 = 32'd1728
; 
32'd129704: dataIn1 = 32'd2772
; 
32'd129705: dataIn1 = 32'd2773
; 
32'd129706: dataIn1 = 32'd2775
; 
32'd129707: dataIn1 = 32'd3055
; 
32'd129708: dataIn1 = 32'd3056
; 
32'd129709: dataIn1 = 32'd3058
; 
32'd129710: dataIn1 = 32'd1729
; 
32'd129711: dataIn1 = 32'd2778
; 
32'd129712: dataIn1 = 32'd2779
; 
32'd129713: dataIn1 = 32'd2781
; 
32'd129714: dataIn1 = 32'd3042
; 
32'd129715: dataIn1 = 32'd3043
; 
32'd129716: dataIn1 = 32'd3046
; 
32'd129717: dataIn1 = 32'd1730
; 
32'd129718: dataIn1 = 32'd2777
; 
32'd129719: dataIn1 = 32'd2779
; 
32'd129720: dataIn1 = 32'd2780
; 
32'd129721: dataIn1 = 32'd3055
; 
32'd129722: dataIn1 = 32'd3057
; 
32'd129723: dataIn1 = 32'd3059
; 
32'd129724: dataIn1 = 32'd1731
; 
32'd129725: dataIn1 = 32'd2782
; 
32'd129726: dataIn1 = 32'd2784
; 
32'd129727: dataIn1 = 32'd2786
; 
32'd129728: dataIn1 = 32'd3062
; 
32'd129729: dataIn1 = 32'd3064
; 
32'd129730: dataIn1 = 32'd3067
; 
32'd129731: dataIn1 = 32'd1732
; 
32'd129732: dataIn1 = 32'd2782
; 
32'd129733: dataIn1 = 32'd2783
; 
32'd129734: dataIn1 = 32'd2785
; 
32'd129735: dataIn1 = 32'd3069
; 
32'd129736: dataIn1 = 32'd3071
; 
32'd129737: dataIn1 = 32'd3074
; 
32'd129738: dataIn1 = 32'd1733
; 
32'd129739: dataIn1 = 32'd2788
; 
32'd129740: dataIn1 = 32'd2789
; 
32'd129741: dataIn1 = 32'd2791
; 
32'd129742: dataIn1 = 32'd3070
; 
32'd129743: dataIn1 = 32'd3071
; 
32'd129744: dataIn1 = 32'd3075
; 
32'd129745: dataIn1 = 32'd1734
; 
32'd129746: dataIn1 = 32'd2787
; 
32'd129747: dataIn1 = 32'd2788
; 
32'd129748: dataIn1 = 32'd2790
; 
32'd129749: dataIn1 = 32'd3076
; 
32'd129750: dataIn1 = 32'd3077
; 
32'd129751: dataIn1 = 32'd3079
; 
32'd129752: dataIn1 = 32'd1735
; 
32'd129753: dataIn1 = 32'd2792
; 
32'd129754: dataIn1 = 32'd2794
; 
32'd129755: dataIn1 = 32'd2796
; 
32'd129756: dataIn1 = 32'd3090
; 
32'd129757: dataIn1 = 32'd3092
; 
32'd129758: dataIn1 = 32'd3095
; 
32'd129759: dataIn1 = 32'd1736
; 
32'd129760: dataIn1 = 32'd2792
; 
32'd129761: dataIn1 = 32'd2793
; 
32'd129762: dataIn1 = 32'd2795
; 
32'd129763: dataIn1 = 32'd3083
; 
32'd129764: dataIn1 = 32'd3084
; 
32'd129765: dataIn1 = 32'd3087
; 
32'd129766: dataIn1 = 32'd1737
; 
32'd129767: dataIn1 = 32'd2798
; 
32'd129768: dataIn1 = 32'd2799
; 
32'd129769: dataIn1 = 32'd2801
; 
32'd129770: dataIn1 = 32'd3105
; 
32'd129771: dataIn1 = 32'd3106
; 
32'd129772: dataIn1 = 32'd3109
; 
32'd129773: dataIn1 = 32'd1738
; 
32'd129774: dataIn1 = 32'd2797
; 
32'd129775: dataIn1 = 32'd2799
; 
32'd129776: dataIn1 = 32'd2800
; 
32'd129777: dataIn1 = 32'd3097
; 
32'd129778: dataIn1 = 32'd3099
; 
32'd129779: dataIn1 = 32'd3101
; 
32'd129780: dataIn1 = 32'd1739
; 
32'd129781: dataIn1 = 32'd2803
; 
32'd129782: dataIn1 = 32'd2804
; 
32'd129783: dataIn1 = 32'd2806
; 
32'd129784: dataIn1 = 32'd3091
; 
32'd129785: dataIn1 = 32'd3092
; 
32'd129786: dataIn1 = 32'd3096
; 
32'd129787: dataIn1 = 32'd1740
; 
32'd129788: dataIn1 = 32'd2802
; 
32'd129789: dataIn1 = 32'd2803
; 
32'd129790: dataIn1 = 32'd2805
; 
32'd129791: dataIn1 = 32'd3097
; 
32'd129792: dataIn1 = 32'd3098
; 
32'd129793: dataIn1 = 32'd3100
; 
32'd129794: dataIn1 = 32'd1741
; 
32'd129795: dataIn1 = 32'd2807
; 
32'd129796: dataIn1 = 32'd2809
; 
32'd129797: dataIn1 = 32'd2811
; 
32'd129798: dataIn1 = 32'd3076
; 
32'd129799: dataIn1 = 32'd3078
; 
32'd129800: dataIn1 = 32'd3080
; 
32'd129801: dataIn1 = 32'd1742
; 
32'd129802: dataIn1 = 32'd2807
; 
32'd129803: dataIn1 = 32'd2808
; 
32'd129804: dataIn1 = 32'd2810
; 
32'd129805: dataIn1 = 32'd3104
; 
32'd129806: dataIn1 = 32'd3105
; 
32'd129807: dataIn1 = 32'd3108
; 
32'd129808: dataIn1 = 32'd1743
; 
32'd129809: dataIn1 = 32'd2813
; 
32'd129810: dataIn1 = 32'd2814
; 
32'd129811: dataIn1 = 32'd2816
; 
32'd129812: dataIn1 = 32'd3119
; 
32'd129813: dataIn1 = 32'd3120
; 
32'd129814: dataIn1 = 32'd3124
; 
32'd129815: dataIn1 = 32'd1744
; 
32'd129816: dataIn1 = 32'd2812
; 
32'd129817: dataIn1 = 32'd2813
; 
32'd129818: dataIn1 = 32'd2815
; 
32'd129819: dataIn1 = 32'd3111
; 
32'd129820: dataIn1 = 32'd3112
; 
32'd129821: dataIn1 = 32'd3114
; 
32'd129822: dataIn1 = 32'd1745
; 
32'd129823: dataIn1 = 32'd2818
; 
32'd129824: dataIn1 = 32'd2819
; 
32'd129825: dataIn1 = 32'd2821
; 
32'd129826: dataIn1 = 32'd3084
; 
32'd129827: dataIn1 = 32'd3085
; 
32'd129828: dataIn1 = 32'd3088
; 
32'd129829: dataIn1 = 32'd1746
; 
32'd129830: dataIn1 = 32'd2817
; 
32'd129831: dataIn1 = 32'd2819
; 
32'd129832: dataIn1 = 32'd2820
; 
32'd129833: dataIn1 = 32'd3111
; 
32'd129834: dataIn1 = 32'd3113
; 
32'd129835: dataIn1 = 32'd3115
; 
32'd129836: dataIn1 = 32'd1747
; 
32'd129837: dataIn1 = 32'd2822
; 
32'd129838: dataIn1 = 32'd2824
; 
32'd129839: dataIn1 = 32'd2826
; 
32'd129840: dataIn1 = 32'd3118
; 
32'd129841: dataIn1 = 32'd3120
; 
32'd129842: dataIn1 = 32'd3123
; 
32'd129843: dataIn1 = 32'd1748
; 
32'd129844: dataIn1 = 32'd2822
; 
32'd129845: dataIn1 = 32'd2823
; 
32'd129846: dataIn1 = 32'd2825
; 
32'd129847: dataIn1 = 32'd3125
; 
32'd129848: dataIn1 = 32'd3127
; 
32'd129849: dataIn1 = 32'd3130
; 
32'd129850: dataIn1 = 32'd1749
; 
32'd129851: dataIn1 = 32'd2828
; 
32'd129852: dataIn1 = 32'd2829
; 
32'd129853: dataIn1 = 32'd2831
; 
32'd129854: dataIn1 = 32'd3126
; 
32'd129855: dataIn1 = 32'd3127
; 
32'd129856: dataIn1 = 32'd3131
; 
32'd129857: dataIn1 = 32'd1750
; 
32'd129858: dataIn1 = 32'd2827
; 
32'd129859: dataIn1 = 32'd2828
; 
32'd129860: dataIn1 = 32'd2830
; 
32'd129861: dataIn1 = 32'd3132
; 
32'd129862: dataIn1 = 32'd3133
; 
32'd129863: dataIn1 = 32'd3135
; 
32'd129864: dataIn1 = 32'd1751
; 
32'd129865: dataIn1 = 32'd2832
; 
32'd129866: dataIn1 = 32'd2834
; 
32'd129867: dataIn1 = 32'd2836
; 
32'd129868: dataIn1 = 32'd3146
; 
32'd129869: dataIn1 = 32'd3148
; 
32'd129870: dataIn1 = 32'd3151
; 
32'd129871: dataIn1 = 32'd1752
; 
32'd129872: dataIn1 = 32'd2832
; 
32'd129873: dataIn1 = 32'd2833
; 
32'd129874: dataIn1 = 32'd2835
; 
32'd129875: dataIn1 = 32'd3139
; 
32'd129876: dataIn1 = 32'd3140
; 
32'd129877: dataIn1 = 32'd3143
; 
32'd129878: dataIn1 = 32'd1753
; 
32'd129879: dataIn1 = 32'd2838
; 
32'd129880: dataIn1 = 32'd2839
; 
32'd129881: dataIn1 = 32'd2841
; 
32'd129882: dataIn1 = 32'd3161
; 
32'd129883: dataIn1 = 32'd3162
; 
32'd129884: dataIn1 = 32'd3165
; 
32'd129885: dataIn1 = 32'd1754
; 
32'd129886: dataIn1 = 32'd2837
; 
32'd129887: dataIn1 = 32'd2839
; 
32'd129888: dataIn1 = 32'd2840
; 
32'd129889: dataIn1 = 32'd3153
; 
32'd129890: dataIn1 = 32'd3155
; 
32'd129891: dataIn1 = 32'd3157
; 
32'd129892: dataIn1 = 32'd1755
; 
32'd129893: dataIn1 = 32'd2843
; 
32'd129894: dataIn1 = 32'd2844
; 
32'd129895: dataIn1 = 32'd2846
; 
32'd129896: dataIn1 = 32'd3147
; 
32'd129897: dataIn1 = 32'd3148
; 
32'd129898: dataIn1 = 32'd3152
; 
32'd129899: dataIn1 = 32'd1756
; 
32'd129900: dataIn1 = 32'd2842
; 
32'd129901: dataIn1 = 32'd2843
; 
32'd129902: dataIn1 = 32'd2845
; 
32'd129903: dataIn1 = 32'd3153
; 
32'd129904: dataIn1 = 32'd3154
; 
32'd129905: dataIn1 = 32'd3156
; 
32'd129906: dataIn1 = 32'd1757
; 
32'd129907: dataIn1 = 32'd2847
; 
32'd129908: dataIn1 = 32'd2849
; 
32'd129909: dataIn1 = 32'd2851
; 
32'd129910: dataIn1 = 32'd3132
; 
32'd129911: dataIn1 = 32'd3134
; 
32'd129912: dataIn1 = 32'd3136
; 
32'd129913: dataIn1 = 32'd1758
; 
32'd129914: dataIn1 = 32'd2847
; 
32'd129915: dataIn1 = 32'd2848
; 
32'd129916: dataIn1 = 32'd2850
; 
32'd129917: dataIn1 = 32'd3160
; 
32'd129918: dataIn1 = 32'd3161
; 
32'd129919: dataIn1 = 32'd3164
; 
32'd129920: dataIn1 = 32'd1759
; 
32'd129921: dataIn1 = 32'd2853
; 
32'd129922: dataIn1 = 32'd2854
; 
32'd129923: dataIn1 = 32'd2856
; 
32'd129924: dataIn1 = 32'd3175
; 
32'd129925: dataIn1 = 32'd3176
; 
32'd129926: dataIn1 = 32'd3180
; 
32'd129927: dataIn1 = 32'd1760
; 
32'd129928: dataIn1 = 32'd2852
; 
32'd129929: dataIn1 = 32'd2853
; 
32'd129930: dataIn1 = 32'd2855
; 
32'd129931: dataIn1 = 32'd3167
; 
32'd129932: dataIn1 = 32'd3168
; 
32'd129933: dataIn1 = 32'd3170
; 
32'd129934: dataIn1 = 32'd1761
; 
32'd129935: dataIn1 = 32'd2858
; 
32'd129936: dataIn1 = 32'd2859
; 
32'd129937: dataIn1 = 32'd2861
; 
32'd129938: dataIn1 = 32'd3140
; 
32'd129939: dataIn1 = 32'd3141
; 
32'd129940: dataIn1 = 32'd3144
; 
32'd129941: dataIn1 = 32'd1762
; 
32'd129942: dataIn1 = 32'd2857
; 
32'd129943: dataIn1 = 32'd2859
; 
32'd129944: dataIn1 = 32'd2860
; 
32'd129945: dataIn1 = 32'd3167
; 
32'd129946: dataIn1 = 32'd3169
; 
32'd129947: dataIn1 = 32'd3171
; 
32'd129948: dataIn1 = 32'd1763
; 
32'd129949: dataIn1 = 32'd2862
; 
32'd129950: dataIn1 = 32'd2864
; 
32'd129951: dataIn1 = 32'd2866
; 
32'd129952: dataIn1 = 32'd3174
; 
32'd129953: dataIn1 = 32'd3176
; 
32'd129954: dataIn1 = 32'd3179
; 
32'd129955: dataIn1 = 32'd1764
; 
32'd129956: dataIn1 = 32'd2862
; 
32'd129957: dataIn1 = 32'd2863
; 
32'd129958: dataIn1 = 32'd2865
; 
32'd129959: dataIn1 = 32'd3181
; 
32'd129960: dataIn1 = 32'd3183
; 
32'd129961: dataIn1 = 32'd3186
; 
32'd129962: dataIn1 = 32'd1765
; 
32'd129963: dataIn1 = 32'd2868
; 
32'd129964: dataIn1 = 32'd2869
; 
32'd129965: dataIn1 = 32'd2871
; 
32'd129966: dataIn1 = 32'd3182
; 
32'd129967: dataIn1 = 32'd3183
; 
32'd129968: dataIn1 = 32'd3187
; 
32'd129969: dataIn1 = 32'd1766
; 
32'd129970: dataIn1 = 32'd2867
; 
32'd129971: dataIn1 = 32'd2868
; 
32'd129972: dataIn1 = 32'd2870
; 
32'd129973: dataIn1 = 32'd3188
; 
32'd129974: dataIn1 = 32'd3189
; 
32'd129975: dataIn1 = 32'd3191
; 
32'd129976: dataIn1 = 32'd1767
; 
32'd129977: dataIn1 = 32'd2872
; 
32'd129978: dataIn1 = 32'd2874
; 
32'd129979: dataIn1 = 32'd2876
; 
32'd129980: dataIn1 = 32'd3202
; 
32'd129981: dataIn1 = 32'd3204
; 
32'd129982: dataIn1 = 32'd3207
; 
32'd129983: dataIn1 = 32'd1768
; 
32'd129984: dataIn1 = 32'd2872
; 
32'd129985: dataIn1 = 32'd2873
; 
32'd129986: dataIn1 = 32'd2875
; 
32'd129987: dataIn1 = 32'd3195
; 
32'd129988: dataIn1 = 32'd3196
; 
32'd129989: dataIn1 = 32'd3199
; 
32'd129990: dataIn1 = 32'd1769
; 
32'd129991: dataIn1 = 32'd2878
; 
32'd129992: dataIn1 = 32'd2879
; 
32'd129993: dataIn1 = 32'd2881
; 
32'd129994: dataIn1 = 32'd3217
; 
32'd129995: dataIn1 = 32'd3218
; 
32'd129996: dataIn1 = 32'd3221
; 
32'd129997: dataIn1 = 32'd1770
; 
32'd129998: dataIn1 = 32'd2877
; 
32'd129999: dataIn1 = 32'd2879
; 
32'd130000: dataIn1 = 32'd2880
; 
32'd130001: dataIn1 = 32'd3209
; 
32'd130002: dataIn1 = 32'd3211
; 
32'd130003: dataIn1 = 32'd3213
; 
32'd130004: dataIn1 = 32'd1771
; 
32'd130005: dataIn1 = 32'd2883
; 
32'd130006: dataIn1 = 32'd2884
; 
32'd130007: dataIn1 = 32'd2886
; 
32'd130008: dataIn1 = 32'd3203
; 
32'd130009: dataIn1 = 32'd3204
; 
32'd130010: dataIn1 = 32'd3208
; 
32'd130011: dataIn1 = 32'd1772
; 
32'd130012: dataIn1 = 32'd2882
; 
32'd130013: dataIn1 = 32'd2883
; 
32'd130014: dataIn1 = 32'd2885
; 
32'd130015: dataIn1 = 32'd3209
; 
32'd130016: dataIn1 = 32'd3210
; 
32'd130017: dataIn1 = 32'd3212
; 
32'd130018: dataIn1 = 32'd1773
; 
32'd130019: dataIn1 = 32'd2887
; 
32'd130020: dataIn1 = 32'd2889
; 
32'd130021: dataIn1 = 32'd2891
; 
32'd130022: dataIn1 = 32'd3188
; 
32'd130023: dataIn1 = 32'd3190
; 
32'd130024: dataIn1 = 32'd3192
; 
32'd130025: dataIn1 = 32'd1774
; 
32'd130026: dataIn1 = 32'd2887
; 
32'd130027: dataIn1 = 32'd2888
; 
32'd130028: dataIn1 = 32'd2890
; 
32'd130029: dataIn1 = 32'd3216
; 
32'd130030: dataIn1 = 32'd3217
; 
32'd130031: dataIn1 = 32'd3220
; 
32'd130032: dataIn1 = 32'd1775
; 
32'd130033: dataIn1 = 32'd2893
; 
32'd130034: dataIn1 = 32'd2894
; 
32'd130035: dataIn1 = 32'd2896
; 
32'd130036: dataIn1 = 32'd3231
; 
32'd130037: dataIn1 = 32'd3232
; 
32'd130038: dataIn1 = 32'd3236
; 
32'd130039: dataIn1 = 32'd1776
; 
32'd130040: dataIn1 = 32'd2892
; 
32'd130041: dataIn1 = 32'd2893
; 
32'd130042: dataIn1 = 32'd2895
; 
32'd130043: dataIn1 = 32'd3223
; 
32'd130044: dataIn1 = 32'd3224
; 
32'd130045: dataIn1 = 32'd3226
; 
32'd130046: dataIn1 = 32'd1777
; 
32'd130047: dataIn1 = 32'd2898
; 
32'd130048: dataIn1 = 32'd2899
; 
32'd130049: dataIn1 = 32'd2901
; 
32'd130050: dataIn1 = 32'd3196
; 
32'd130051: dataIn1 = 32'd3197
; 
32'd130052: dataIn1 = 32'd3200
; 
32'd130053: dataIn1 = 32'd1778
; 
32'd130054: dataIn1 = 32'd2897
; 
32'd130055: dataIn1 = 32'd2899
; 
32'd130056: dataIn1 = 32'd2900
; 
32'd130057: dataIn1 = 32'd3223
; 
32'd130058: dataIn1 = 32'd3225
; 
32'd130059: dataIn1 = 32'd3227
; 
32'd130060: dataIn1 = 32'd1779
; 
32'd130061: dataIn1 = 32'd2902
; 
32'd130062: dataIn1 = 32'd2904
; 
32'd130063: dataIn1 = 32'd2906
; 
32'd130064: dataIn1 = 32'd3230
; 
32'd130065: dataIn1 = 32'd3232
; 
32'd130066: dataIn1 = 32'd3235
; 
32'd130067: dataIn1 = 32'd1780
; 
32'd130068: dataIn1 = 32'd2902
; 
32'd130069: dataIn1 = 32'd2903
; 
32'd130070: dataIn1 = 32'd2905
; 
32'd130071: dataIn1 = 32'd3237
; 
32'd130072: dataIn1 = 32'd3239
; 
32'd130073: dataIn1 = 32'd3242
; 
32'd130074: dataIn1 = 32'd1781
; 
32'd130075: dataIn1 = 32'd2908
; 
32'd130076: dataIn1 = 32'd2909
; 
32'd130077: dataIn1 = 32'd2911
; 
32'd130078: dataIn1 = 32'd3238
; 
32'd130079: dataIn1 = 32'd3239
; 
32'd130080: dataIn1 = 32'd3243
; 
32'd130081: dataIn1 = 32'd1782
; 
32'd130082: dataIn1 = 32'd2907
; 
32'd130083: dataIn1 = 32'd2908
; 
32'd130084: dataIn1 = 32'd2910
; 
32'd130085: dataIn1 = 32'd3244
; 
32'd130086: dataIn1 = 32'd3245
; 
32'd130087: dataIn1 = 32'd3247
; 
32'd130088: dataIn1 = 32'd1783
; 
32'd130089: dataIn1 = 32'd2912
; 
32'd130090: dataIn1 = 32'd2914
; 
32'd130091: dataIn1 = 32'd2916
; 
32'd130092: dataIn1 = 32'd3258
; 
32'd130093: dataIn1 = 32'd3260
; 
32'd130094: dataIn1 = 32'd3263
; 
32'd130095: dataIn1 = 32'd1784
; 
32'd130096: dataIn1 = 32'd2912
; 
32'd130097: dataIn1 = 32'd2913
; 
32'd130098: dataIn1 = 32'd2915
; 
32'd130099: dataIn1 = 32'd3251
; 
32'd130100: dataIn1 = 32'd3252
; 
32'd130101: dataIn1 = 32'd3255
; 
32'd130102: dataIn1 = 32'd1785
; 
32'd130103: dataIn1 = 32'd2918
; 
32'd130104: dataIn1 = 32'd2919
; 
32'd130105: dataIn1 = 32'd2921
; 
32'd130106: dataIn1 = 32'd3273
; 
32'd130107: dataIn1 = 32'd3274
; 
32'd130108: dataIn1 = 32'd3277
; 
32'd130109: dataIn1 = 32'd1786
; 
32'd130110: dataIn1 = 32'd2917
; 
32'd130111: dataIn1 = 32'd2919
; 
32'd130112: dataIn1 = 32'd2920
; 
32'd130113: dataIn1 = 32'd3265
; 
32'd130114: dataIn1 = 32'd3267
; 
32'd130115: dataIn1 = 32'd3269
; 
32'd130116: dataIn1 = 32'd1787
; 
32'd130117: dataIn1 = 32'd2923
; 
32'd130118: dataIn1 = 32'd2924
; 
32'd130119: dataIn1 = 32'd2926
; 
32'd130120: dataIn1 = 32'd3259
; 
32'd130121: dataIn1 = 32'd3260
; 
32'd130122: dataIn1 = 32'd3264
; 
32'd130123: dataIn1 = 32'd1788
; 
32'd130124: dataIn1 = 32'd2922
; 
32'd130125: dataIn1 = 32'd2923
; 
32'd130126: dataIn1 = 32'd2925
; 
32'd130127: dataIn1 = 32'd3265
; 
32'd130128: dataIn1 = 32'd3266
; 
32'd130129: dataIn1 = 32'd3268
; 
32'd130130: dataIn1 = 32'd1789
; 
32'd130131: dataIn1 = 32'd2927
; 
32'd130132: dataIn1 = 32'd2929
; 
32'd130133: dataIn1 = 32'd2931
; 
32'd130134: dataIn1 = 32'd3244
; 
32'd130135: dataIn1 = 32'd3246
; 
32'd130136: dataIn1 = 32'd3248
; 
32'd130137: dataIn1 = 32'd1790
; 
32'd130138: dataIn1 = 32'd2927
; 
32'd130139: dataIn1 = 32'd2928
; 
32'd130140: dataIn1 = 32'd2930
; 
32'd130141: dataIn1 = 32'd3272
; 
32'd130142: dataIn1 = 32'd3273
; 
32'd130143: dataIn1 = 32'd3276
; 
32'd130144: dataIn1 = 32'd1791
; 
32'd130145: dataIn1 = 32'd2933
; 
32'd130146: dataIn1 = 32'd2934
; 
32'd130147: dataIn1 = 32'd2936
; 
32'd130148: dataIn1 = 32'd3287
; 
32'd130149: dataIn1 = 32'd3288
; 
32'd130150: dataIn1 = 32'd3292
; 
32'd130151: dataIn1 = 32'd1792
; 
32'd130152: dataIn1 = 32'd2932
; 
32'd130153: dataIn1 = 32'd2933
; 
32'd130154: dataIn1 = 32'd2935
; 
32'd130155: dataIn1 = 32'd3279
; 
32'd130156: dataIn1 = 32'd3280
; 
32'd130157: dataIn1 = 32'd3282
; 
32'd130158: dataIn1 = 32'd1793
; 
32'd130159: dataIn1 = 32'd2938
; 
32'd130160: dataIn1 = 32'd2939
; 
32'd130161: dataIn1 = 32'd2941
; 
32'd130162: dataIn1 = 32'd3252
; 
32'd130163: dataIn1 = 32'd3253
; 
32'd130164: dataIn1 = 32'd3256
; 
32'd130165: dataIn1 = 32'd1794
; 
32'd130166: dataIn1 = 32'd2937
; 
32'd130167: dataIn1 = 32'd2939
; 
32'd130168: dataIn1 = 32'd2940
; 
32'd130169: dataIn1 = 32'd3279
; 
32'd130170: dataIn1 = 32'd3281
; 
32'd130171: dataIn1 = 32'd3283
; 
32'd130172: dataIn1 = 32'd1795
; 
32'd130173: dataIn1 = 32'd2942
; 
32'd130174: dataIn1 = 32'd2944
; 
32'd130175: dataIn1 = 32'd2946
; 
32'd130176: dataIn1 = 32'd3286
; 
32'd130177: dataIn1 = 32'd3288
; 
32'd130178: dataIn1 = 32'd3291
; 
32'd130179: dataIn1 = 32'd1796
; 
32'd130180: dataIn1 = 32'd2942
; 
32'd130181: dataIn1 = 32'd2943
; 
32'd130182: dataIn1 = 32'd2945
; 
32'd130183: dataIn1 = 32'd3293
; 
32'd130184: dataIn1 = 32'd3295
; 
32'd130185: dataIn1 = 32'd3298
; 
32'd130186: dataIn1 = 32'd1797
; 
32'd130187: dataIn1 = 32'd2948
; 
32'd130188: dataIn1 = 32'd2949
; 
32'd130189: dataIn1 = 32'd2951
; 
32'd130190: dataIn1 = 32'd3294
; 
32'd130191: dataIn1 = 32'd3295
; 
32'd130192: dataIn1 = 32'd3299
; 
32'd130193: dataIn1 = 32'd1798
; 
32'd130194: dataIn1 = 32'd2947
; 
32'd130195: dataIn1 = 32'd2948
; 
32'd130196: dataIn1 = 32'd2950
; 
32'd130197: dataIn1 = 32'd3300
; 
32'd130198: dataIn1 = 32'd3301
; 
32'd130199: dataIn1 = 32'd3303
; 
32'd130200: dataIn1 = 32'd1799
; 
32'd130201: dataIn1 = 32'd2952
; 
32'd130202: dataIn1 = 32'd2954
; 
32'd130203: dataIn1 = 32'd2956
; 
32'd130204: dataIn1 = 32'd3314
; 
32'd130205: dataIn1 = 32'd3316
; 
32'd130206: dataIn1 = 32'd3319
; 
32'd130207: dataIn1 = 32'd1800
; 
32'd130208: dataIn1 = 32'd2952
; 
32'd130209: dataIn1 = 32'd2953
; 
32'd130210: dataIn1 = 32'd2955
; 
32'd130211: dataIn1 = 32'd3307
; 
32'd130212: dataIn1 = 32'd3308
; 
32'd130213: dataIn1 = 32'd3311
; 
32'd130214: dataIn1 = 32'd1801
; 
32'd130215: dataIn1 = 32'd2958
; 
32'd130216: dataIn1 = 32'd2959
; 
32'd130217: dataIn1 = 32'd2961
; 
32'd130218: dataIn1 = 32'd3329
; 
32'd130219: dataIn1 = 32'd3330
; 
32'd130220: dataIn1 = 32'd3333
; 
32'd130221: dataIn1 = 32'd1802
; 
32'd130222: dataIn1 = 32'd2957
; 
32'd130223: dataIn1 = 32'd2959
; 
32'd130224: dataIn1 = 32'd2960
; 
32'd130225: dataIn1 = 32'd3321
; 
32'd130226: dataIn1 = 32'd3323
; 
32'd130227: dataIn1 = 32'd3325
; 
32'd130228: dataIn1 = 32'd1803
; 
32'd130229: dataIn1 = 32'd2963
; 
32'd130230: dataIn1 = 32'd2964
; 
32'd130231: dataIn1 = 32'd2966
; 
32'd130232: dataIn1 = 32'd3315
; 
32'd130233: dataIn1 = 32'd3316
; 
32'd130234: dataIn1 = 32'd3320
; 
32'd130235: dataIn1 = 32'd1804
; 
32'd130236: dataIn1 = 32'd2962
; 
32'd130237: dataIn1 = 32'd2963
; 
32'd130238: dataIn1 = 32'd2965
; 
32'd130239: dataIn1 = 32'd3321
; 
32'd130240: dataIn1 = 32'd3322
; 
32'd130241: dataIn1 = 32'd3324
; 
32'd130242: dataIn1 = 32'd1805
; 
32'd130243: dataIn1 = 32'd2967
; 
32'd130244: dataIn1 = 32'd2969
; 
32'd130245: dataIn1 = 32'd2971
; 
32'd130246: dataIn1 = 32'd3300
; 
32'd130247: dataIn1 = 32'd3302
; 
32'd130248: dataIn1 = 32'd3304
; 
32'd130249: dataIn1 = 32'd1806
; 
32'd130250: dataIn1 = 32'd2967
; 
32'd130251: dataIn1 = 32'd2968
; 
32'd130252: dataIn1 = 32'd2970
; 
32'd130253: dataIn1 = 32'd3328
; 
32'd130254: dataIn1 = 32'd3329
; 
32'd130255: dataIn1 = 32'd3332
; 
32'd130256: dataIn1 = 32'd1807
; 
32'd130257: dataIn1 = 32'd2973
; 
32'd130258: dataIn1 = 32'd2974
; 
32'd130259: dataIn1 = 32'd2976
; 
32'd130260: dataIn1 = 32'd3343
; 
32'd130261: dataIn1 = 32'd3344
; 
32'd130262: dataIn1 = 32'd3348
; 
32'd130263: dataIn1 = 32'd1808
; 
32'd130264: dataIn1 = 32'd2972
; 
32'd130265: dataIn1 = 32'd2973
; 
32'd130266: dataIn1 = 32'd2975
; 
32'd130267: dataIn1 = 32'd3335
; 
32'd130268: dataIn1 = 32'd3336
; 
32'd130269: dataIn1 = 32'd3338
; 
32'd130270: dataIn1 = 32'd1809
; 
32'd130271: dataIn1 = 32'd2978
; 
32'd130272: dataIn1 = 32'd2979
; 
32'd130273: dataIn1 = 32'd2981
; 
32'd130274: dataIn1 = 32'd3308
; 
32'd130275: dataIn1 = 32'd3309
; 
32'd130276: dataIn1 = 32'd3312
; 
32'd130277: dataIn1 = 32'd1810
; 
32'd130278: dataIn1 = 32'd2977
; 
32'd130279: dataIn1 = 32'd2979
; 
32'd130280: dataIn1 = 32'd2980
; 
32'd130281: dataIn1 = 32'd3335
; 
32'd130282: dataIn1 = 32'd3337
; 
32'd130283: dataIn1 = 32'd3339
; 
32'd130284: dataIn1 = 32'd1811
; 
32'd130285: dataIn1 = 32'd2982
; 
32'd130286: dataIn1 = 32'd2984
; 
32'd130287: dataIn1 = 32'd2986
; 
32'd130288: dataIn1 = 32'd3342
; 
32'd130289: dataIn1 = 32'd3344
; 
32'd130290: dataIn1 = 32'd3347
; 
32'd130291: dataIn1 = 32'd1812
; 
32'd130292: dataIn1 = 32'd2982
; 
32'd130293: dataIn1 = 32'd2983
; 
32'd130294: dataIn1 = 32'd2985
; 
32'd130295: dataIn1 = 32'd3349
; 
32'd130296: dataIn1 = 32'd3351
; 
32'd130297: dataIn1 = 32'd3354
; 
32'd130298: dataIn1 = 32'd1813
; 
32'd130299: dataIn1 = 32'd2988
; 
32'd130300: dataIn1 = 32'd2989
; 
32'd130301: dataIn1 = 32'd2991
; 
32'd130302: dataIn1 = 32'd3350
; 
32'd130303: dataIn1 = 32'd3351
; 
32'd130304: dataIn1 = 32'd3355
; 
32'd130305: dataIn1 = 32'd1814
; 
32'd130306: dataIn1 = 32'd2987
; 
32'd130307: dataIn1 = 32'd2988
; 
32'd130308: dataIn1 = 32'd2990
; 
32'd130309: dataIn1 = 32'd3356
; 
32'd130310: dataIn1 = 32'd3357
; 
32'd130311: dataIn1 = 32'd3359
; 
32'd130312: dataIn1 = 32'd1815
; 
32'd130313: dataIn1 = 32'd2992
; 
32'd130314: dataIn1 = 32'd2994
; 
32'd130315: dataIn1 = 32'd2996
; 
32'd130316: dataIn1 = 32'd3370
; 
32'd130317: dataIn1 = 32'd3372
; 
32'd130318: dataIn1 = 32'd3375
; 
32'd130319: dataIn1 = 32'd1816
; 
32'd130320: dataIn1 = 32'd2992
; 
32'd130321: dataIn1 = 32'd2993
; 
32'd130322: dataIn1 = 32'd2995
; 
32'd130323: dataIn1 = 32'd3363
; 
32'd130324: dataIn1 = 32'd3364
; 
32'd130325: dataIn1 = 32'd3367
; 
32'd130326: dataIn1 = 32'd1817
; 
32'd130327: dataIn1 = 32'd2998
; 
32'd130328: dataIn1 = 32'd2999
; 
32'd130329: dataIn1 = 32'd3001
; 
32'd130330: dataIn1 = 32'd3385
; 
32'd130331: dataIn1 = 32'd3386
; 
32'd130332: dataIn1 = 32'd3389
; 
32'd130333: dataIn1 = 32'd1818
; 
32'd130334: dataIn1 = 32'd2997
; 
32'd130335: dataIn1 = 32'd2999
; 
32'd130336: dataIn1 = 32'd3000
; 
32'd130337: dataIn1 = 32'd3377
; 
32'd130338: dataIn1 = 32'd3379
; 
32'd130339: dataIn1 = 32'd3381
; 
32'd130340: dataIn1 = 32'd1819
; 
32'd130341: dataIn1 = 32'd3003
; 
32'd130342: dataIn1 = 32'd3004
; 
32'd130343: dataIn1 = 32'd3006
; 
32'd130344: dataIn1 = 32'd3371
; 
32'd130345: dataIn1 = 32'd3372
; 
32'd130346: dataIn1 = 32'd3376
; 
32'd130347: dataIn1 = 32'd1820
; 
32'd130348: dataIn1 = 32'd3002
; 
32'd130349: dataIn1 = 32'd3003
; 
32'd130350: dataIn1 = 32'd3005
; 
32'd130351: dataIn1 = 32'd3377
; 
32'd130352: dataIn1 = 32'd3378
; 
32'd130353: dataIn1 = 32'd3380
; 
32'd130354: dataIn1 = 32'd1821
; 
32'd130355: dataIn1 = 32'd3007
; 
32'd130356: dataIn1 = 32'd3009
; 
32'd130357: dataIn1 = 32'd3011
; 
32'd130358: dataIn1 = 32'd3356
; 
32'd130359: dataIn1 = 32'd3358
; 
32'd130360: dataIn1 = 32'd3360
; 
32'd130361: dataIn1 = 32'd1822
; 
32'd130362: dataIn1 = 32'd3007
; 
32'd130363: dataIn1 = 32'd3008
; 
32'd130364: dataIn1 = 32'd3010
; 
32'd130365: dataIn1 = 32'd3384
; 
32'd130366: dataIn1 = 32'd3385
; 
32'd130367: dataIn1 = 32'd3388
; 
32'd130368: dataIn1 = 32'd1823
; 
32'd130369: dataIn1 = 32'd3013
; 
32'd130370: dataIn1 = 32'd3014
; 
32'd130371: dataIn1 = 32'd3016
; 
32'd130372: dataIn1 = 32'd3399
; 
32'd130373: dataIn1 = 32'd3400
; 
32'd130374: dataIn1 = 32'd3404
; 
32'd130375: dataIn1 = 32'd1824
; 
32'd130376: dataIn1 = 32'd3012
; 
32'd130377: dataIn1 = 32'd3013
; 
32'd130378: dataIn1 = 32'd3015
; 
32'd130379: dataIn1 = 32'd3391
; 
32'd130380: dataIn1 = 32'd3392
; 
32'd130381: dataIn1 = 32'd3394
; 
32'd130382: dataIn1 = 32'd1825
; 
32'd130383: dataIn1 = 32'd3018
; 
32'd130384: dataIn1 = 32'd3019
; 
32'd130385: dataIn1 = 32'd3021
; 
32'd130386: dataIn1 = 32'd3364
; 
32'd130387: dataIn1 = 32'd3365
; 
32'd130388: dataIn1 = 32'd3368
; 
32'd130389: dataIn1 = 32'd1826
; 
32'd130390: dataIn1 = 32'd3017
; 
32'd130391: dataIn1 = 32'd3019
; 
32'd130392: dataIn1 = 32'd3020
; 
32'd130393: dataIn1 = 32'd3391
; 
32'd130394: dataIn1 = 32'd3393
; 
32'd130395: dataIn1 = 32'd3395
; 
32'd130396: dataIn1 = 32'd1827
; 
32'd130397: dataIn1 = 32'd3022
; 
32'd130398: dataIn1 = 32'd3024
; 
32'd130399: dataIn1 = 32'd3026
; 
32'd130400: dataIn1 = 32'd3398
; 
32'd130401: dataIn1 = 32'd3400
; 
32'd130402: dataIn1 = 32'd3403
; 
32'd130403: dataIn1 = 32'd1828
; 
32'd130404: dataIn1 = 32'd3022
; 
32'd130405: dataIn1 = 32'd3023
; 
32'd130406: dataIn1 = 32'd3025
; 
32'd130407: dataIn1 = 32'd3441
; 
32'd130408: dataIn1 = 32'd731
; 
32'd130409: dataIn1 = 32'd962
; 
32'd130410: dataIn1 = 32'd1397
; 
32'd130411: dataIn1 = 32'd1398
; 
32'd130412: dataIn1 = 32'd1829
; 
32'd130413: dataIn1 = 32'd1830
; 
32'd130414: dataIn1 = 32'd1832
; 
32'd130415: dataIn1 = 32'd2030
; 
32'd130416: dataIn1 = 32'd194
; 
32'd130417: dataIn1 = 32'd962
; 
32'd130418: dataIn1 = 32'd1397
; 
32'd130419: dataIn1 = 32'd1401
; 
32'd130420: dataIn1 = 32'd1829
; 
32'd130421: dataIn1 = 32'd1830
; 
32'd130422: dataIn1 = 32'd1834
; 
32'd130423: dataIn1 = 32'd2029
; 
32'd130424: dataIn1 = 32'd732
; 
32'd130425: dataIn1 = 32'd961
; 
32'd130426: dataIn1 = 32'd1399
; 
32'd130427: dataIn1 = 32'd1400
; 
32'd130428: dataIn1 = 32'd1831
; 
32'd130429: dataIn1 = 32'd1832
; 
32'd130430: dataIn1 = 32'd1839
; 
32'd130431: dataIn1 = 32'd2031
; 
32'd130432: dataIn1 = 32'd383
; 
32'd130433: dataIn1 = 32'd961
; 
32'd130434: dataIn1 = 32'd1398
; 
32'd130435: dataIn1 = 32'd1399
; 
32'd130436: dataIn1 = 32'd1829
; 
32'd130437: dataIn1 = 32'd1831
; 
32'd130438: dataIn1 = 32'd1832
; 
32'd130439: dataIn1 = 32'd2030
; 
32'd130440: dataIn1 = 32'd384
; 
32'd130441: dataIn1 = 32'd964
; 
32'd130442: dataIn1 = 32'd1402
; 
32'd130443: dataIn1 = 32'd1404
; 
32'd130444: dataIn1 = 32'd1833
; 
32'd130445: dataIn1 = 32'd1834
; 
32'd130446: dataIn1 = 32'd1835
; 
32'd130447: dataIn1 = 32'd2032
; 
32'd130448: dataIn1 = 32'd733
; 
32'd130449: dataIn1 = 32'd964
; 
32'd130450: dataIn1 = 32'd1401
; 
32'd130451: dataIn1 = 32'd1402
; 
32'd130452: dataIn1 = 32'd1830
; 
32'd130453: dataIn1 = 32'd1833
; 
32'd130454: dataIn1 = 32'd1834
; 
32'd130455: dataIn1 = 32'd2029
; 
32'd130456: dataIn1 = 32'd734
; 
32'd130457: dataIn1 = 32'd963
; 
32'd130458: dataIn1 = 32'd1403
; 
32'd130459: dataIn1 = 32'd1404
; 
32'd130460: dataIn1 = 32'd1833
; 
32'd130461: dataIn1 = 32'd1835
; 
32'd130462: dataIn1 = 32'd1836
; 
32'd130463: dataIn1 = 32'd2032
; 
32'd130464: dataIn1 = 32'd197
; 
32'd130465: dataIn1 = 32'd963
; 
32'd130466: dataIn1 = 32'd1403
; 
32'd130467: dataIn1 = 32'd1835
; 
32'd130468: dataIn1 = 32'd1836
; 
32'd130469: dataIn1 = 32'd198
; 
32'd130470: dataIn1 = 32'd735
; 
32'd130471: dataIn1 = 32'd966
; 
32'd130472: dataIn1 = 32'd1405
; 
32'd130473: dataIn1 = 32'd1406
; 
32'd130474: dataIn1 = 32'd1837
; 
32'd130475: dataIn1 = 32'd1838
; 
32'd130476: dataIn1 = 32'd1841
; 
32'd130477: dataIn1 = 32'd2034
; 
32'd130478: dataIn1 = 32'd385
; 
32'd130479: dataIn1 = 32'd966
; 
32'd130480: dataIn1 = 32'd1405
; 
32'd130481: dataIn1 = 32'd1407
; 
32'd130482: dataIn1 = 32'd1837
; 
32'd130483: dataIn1 = 32'd1838
; 
32'd130484: dataIn1 = 32'd1840
; 
32'd130485: dataIn1 = 32'd2033
; 
32'd130486: dataIn1 = 32'd196
; 
32'd130487: dataIn1 = 32'd965
; 
32'd130488: dataIn1 = 32'd1400
; 
32'd130489: dataIn1 = 32'd1408
; 
32'd130490: dataIn1 = 32'd1831
; 
32'd130491: dataIn1 = 32'd1839
; 
32'd130492: dataIn1 = 32'd1840
; 
32'd130493: dataIn1 = 32'd2031
; 
32'd130494: dataIn1 = 32'd736
; 
32'd130495: dataIn1 = 32'd965
; 
32'd130496: dataIn1 = 32'd1407
; 
32'd130497: dataIn1 = 32'd1408
; 
32'd130498: dataIn1 = 32'd1838
; 
32'd130499: dataIn1 = 32'd1839
; 
32'd130500: dataIn1 = 32'd1840
; 
32'd130501: dataIn1 = 32'd2033
; 
32'd130502: dataIn1 = 32'd198
; 
32'd130503: dataIn1 = 32'd737
; 
32'd130504: dataIn1 = 32'd968
; 
32'd130505: dataIn1 = 32'd1410
; 
32'd130506: dataIn1 = 32'd1837
; 
32'd130507: dataIn1 = 32'd1841
; 
32'd130508: dataIn1 = 32'd1842
; 
32'd130509: dataIn1 = 32'd2034
; 
32'd130510: dataIn1 = 32'd386
; 
32'd130511: dataIn1 = 32'd737
; 
32'd130512: dataIn1 = 32'd968
; 
32'd130513: dataIn1 = 32'd1409
; 
32'd130514: dataIn1 = 32'd1841
; 
32'd130515: dataIn1 = 32'd1842
; 
32'd130516: dataIn1 = 32'd1844
; 
32'd130517: dataIn1 = 32'd2035
; 
32'd130518: dataIn1 = 32'd200
; 
32'd130519: dataIn1 = 32'd738
; 
32'd130520: dataIn1 = 32'd967
; 
32'd130521: dataIn1 = 32'd1412
; 
32'd130522: dataIn1 = 32'd1843
; 
32'd130523: dataIn1 = 32'd1844
; 
32'd130524: dataIn1 = 32'd1852
; 
32'd130525: dataIn1 = 32'd2036
; 
32'd130526: dataIn1 = 32'd386
; 
32'd130527: dataIn1 = 32'd738
; 
32'd130528: dataIn1 = 32'd967
; 
32'd130529: dataIn1 = 32'd1411
; 
32'd130530: dataIn1 = 32'd1842
; 
32'd130531: dataIn1 = 32'd1843
; 
32'd130532: dataIn1 = 32'd1844
; 
32'd130533: dataIn1 = 32'd2035
; 
32'd130534: dataIn1 = 32'd387
; 
32'd130535: dataIn1 = 32'd739
; 
32'd130536: dataIn1 = 32'd970
; 
32'd130537: dataIn1 = 32'd1414
; 
32'd130538: dataIn1 = 32'd1845
; 
32'd130539: dataIn1 = 32'd1846
; 
32'd130540: dataIn1 = 32'd1848
; 
32'd130541: dataIn1 = 32'd2038
; 
32'd130542: dataIn1 = 32'd201
; 
32'd130543: dataIn1 = 32'd739
; 
32'd130544: dataIn1 = 32'd970
; 
32'd130545: dataIn1 = 32'd1413
; 
32'd130546: dataIn1 = 32'd1845
; 
32'd130547: dataIn1 = 32'd1846
; 
32'd130548: dataIn1 = 32'd1850
; 
32'd130549: dataIn1 = 32'd2037
; 
32'd130550: dataIn1 = 32'd969
; 
32'd130551: dataIn1 = 32'd1847
; 
32'd130552: dataIn1 = 32'd1848
; 
32'd130553: dataIn1 = 32'd3405
; 
32'd130554: dataIn1 = 32'd3407
; 
32'd130555: dataIn1 = 32'd3409
; 
32'd130556: dataIn1 = 32'd3446
; 
32'd130557: dataIn1 = 32'd387
; 
32'd130558: dataIn1 = 32'd740
; 
32'd130559: dataIn1 = 32'd969
; 
32'd130560: dataIn1 = 32'd1415
; 
32'd130561: dataIn1 = 32'd1845
; 
32'd130562: dataIn1 = 32'd1847
; 
32'd130563: dataIn1 = 32'd1848
; 
32'd130564: dataIn1 = 32'd2038
; 
32'd130565: dataIn1 = 32'd3446
; 
32'd130566: dataIn1 = 32'd388
; 
32'd130567: dataIn1 = 32'd741
; 
32'd130568: dataIn1 = 32'd972
; 
32'd130569: dataIn1 = 32'd1418
; 
32'd130570: dataIn1 = 32'd1849
; 
32'd130571: dataIn1 = 32'd1850
; 
32'd130572: dataIn1 = 32'd1851
; 
32'd130573: dataIn1 = 32'd2040
; 
32'd130574: dataIn1 = 32'd201
; 
32'd130575: dataIn1 = 32'd741
; 
32'd130576: dataIn1 = 32'd972
; 
32'd130577: dataIn1 = 32'd1417
; 
32'd130578: dataIn1 = 32'd1846
; 
32'd130579: dataIn1 = 32'd1849
; 
32'd130580: dataIn1 = 32'd1850
; 
32'd130581: dataIn1 = 32'd2037
; 
32'd130582: dataIn1 = 32'd388
; 
32'd130583: dataIn1 = 32'd742
; 
32'd130584: dataIn1 = 32'd971
; 
32'd130585: dataIn1 = 32'd1420
; 
32'd130586: dataIn1 = 32'd1849
; 
32'd130587: dataIn1 = 32'd1851
; 
32'd130588: dataIn1 = 32'd1852
; 
32'd130589: dataIn1 = 32'd2040
; 
32'd130590: dataIn1 = 32'd200
; 
32'd130591: dataIn1 = 32'd742
; 
32'd130592: dataIn1 = 32'd971
; 
32'd130593: dataIn1 = 32'd1419
; 
32'd130594: dataIn1 = 32'd1843
; 
32'd130595: dataIn1 = 32'd1851
; 
32'd130596: dataIn1 = 32'd1852
; 
32'd130597: dataIn1 = 32'd2036
; 
32'd130598: dataIn1 = 32'd1853
; 
32'd130599: dataIn1 = 32'd3028
; 
32'd130600: dataIn1 = 32'd3029
; 
32'd130601: dataIn1 = 32'd3031
; 
32'd130602: dataIn1 = 32'd3406
; 
32'd130603: dataIn1 = 32'd3407
; 
32'd130604: dataIn1 = 32'd3410
; 
32'd130605: dataIn1 = 32'd1854
; 
32'd130606: dataIn1 = 32'd3027
; 
32'd130607: dataIn1 = 32'd3028
; 
32'd130608: dataIn1 = 32'd3030
; 
32'd130609: dataIn1 = 32'd3442
; 
32'd130610: dataIn1 = 32'd3460
; 
32'd130611: dataIn1 = 32'd10256
; 
32'd130612: dataIn1 = 32'd392
; 
32'd130613: dataIn1 = 32'd1855
; 
32'd130614: dataIn1 = 32'd10256
; 
32'd130615: dataIn1 = 32'd10257
; 
32'd130616: dataIn1 = 32'd10263
; 
32'd130617: dataIn1 = 32'd10271
; 
32'd130618: dataIn1 = 32'd10272
; 
32'd130619: dataIn1 = 32'd393
; 
32'd130620: dataIn1 = 32'd1856
; 
32'd130621: dataIn1 = 32'd2041
; 
32'd130622: dataIn1 = 32'd3033
; 
32'd130623: dataIn1 = 32'd3034
; 
32'd130624: dataIn1 = 32'd3414
; 
32'd130625: dataIn1 = 32'd3415
; 
32'd130626: dataIn1 = 32'd393
; 
32'd130627: dataIn1 = 32'd1857
; 
32'd130628: dataIn1 = 32'd3032
; 
32'd130629: dataIn1 = 32'd3034
; 
32'd130630: dataIn1 = 32'd3411
; 
32'd130631: dataIn1 = 32'd3413
; 
32'd130632: dataIn1 = 32'd10270
; 
32'd130633: dataIn1 = 32'd393
; 
32'd130634: dataIn1 = 32'd1858
; 
32'd130635: dataIn1 = 32'd1859
; 
32'd130636: dataIn1 = 32'd10258
; 
32'd130637: dataIn1 = 32'd10259
; 
32'd130638: dataIn1 = 32'd10270
; 
32'd130639: dataIn1 = 32'd10284
; 
32'd130640: dataIn1 = 32'd1
; 
32'd130641: dataIn1 = 32'd393
; 
32'd130642: dataIn1 = 32'd771
; 
32'd130643: dataIn1 = 32'd959
; 
32'd130644: dataIn1 = 32'd1469
; 
32'd130645: dataIn1 = 32'd1858
; 
32'd130646: dataIn1 = 32'd1859
; 
32'd130647: dataIn1 = 32'd2042
; 
32'd130648: dataIn1 = 32'd10284
; 
32'd130649: dataIn1 = 32'd208
; 
32'd130650: dataIn1 = 32'd779
; 
32'd130651: dataIn1 = 32'd975
; 
32'd130652: dataIn1 = 32'd1484
; 
32'd130653: dataIn1 = 32'd1860
; 
32'd130654: dataIn1 = 32'd1861
; 
32'd130655: dataIn1 = 32'd1864
; 
32'd130656: dataIn1 = 32'd2044
; 
32'd130657: dataIn1 = 32'd406
; 
32'd130658: dataIn1 = 32'd779
; 
32'd130659: dataIn1 = 32'd975
; 
32'd130660: dataIn1 = 32'd1483
; 
32'd130661: dataIn1 = 32'd1860
; 
32'd130662: dataIn1 = 32'd1861
; 
32'd130663: dataIn1 = 32'd1863
; 
32'd130664: dataIn1 = 32'd2043
; 
32'd130665: dataIn1 = 32'd207
; 
32'd130666: dataIn1 = 32'd767
; 
32'd130667: dataIn1 = 32'd781
; 
32'd130668: dataIn1 = 32'd973
; 
32'd130669: dataIn1 = 32'd1487
; 
32'd130670: dataIn1 = 32'd1862
; 
32'd130671: dataIn1 = 32'd1863
; 
32'd130672: dataIn1 = 32'd2045
; 
32'd130673: dataIn1 = 32'd406
; 
32'd130674: dataIn1 = 32'd781
; 
32'd130675: dataIn1 = 32'd973
; 
32'd130676: dataIn1 = 32'd1486
; 
32'd130677: dataIn1 = 32'd1861
; 
32'd130678: dataIn1 = 32'd1862
; 
32'd130679: dataIn1 = 32'd1863
; 
32'd130680: dataIn1 = 32'd2043
; 
32'd130681: dataIn1 = 32'd208
; 
32'd130682: dataIn1 = 32'd789
; 
32'd130683: dataIn1 = 32'd978
; 
32'd130684: dataIn1 = 32'd1495
; 
32'd130685: dataIn1 = 32'd1860
; 
32'd130686: dataIn1 = 32'd1864
; 
32'd130687: dataIn1 = 32'd1865
; 
32'd130688: dataIn1 = 32'd2044
; 
32'd130689: dataIn1 = 32'd410
; 
32'd130690: dataIn1 = 32'd789
; 
32'd130691: dataIn1 = 32'd978
; 
32'd130692: dataIn1 = 32'd1494
; 
32'd130693: dataIn1 = 32'd1864
; 
32'd130694: dataIn1 = 32'd1865
; 
32'd130695: dataIn1 = 32'd1867
; 
32'd130696: dataIn1 = 32'd2046
; 
32'd130697: dataIn1 = 32'd210
; 
32'd130698: dataIn1 = 32'd791
; 
32'd130699: dataIn1 = 32'd977
; 
32'd130700: dataIn1 = 32'd1498
; 
32'd130701: dataIn1 = 32'd1866
; 
32'd130702: dataIn1 = 32'd1867
; 
32'd130703: dataIn1 = 32'd1876
; 
32'd130704: dataIn1 = 32'd2047
; 
32'd130705: dataIn1 = 32'd410
; 
32'd130706: dataIn1 = 32'd791
; 
32'd130707: dataIn1 = 32'd977
; 
32'd130708: dataIn1 = 32'd1497
; 
32'd130709: dataIn1 = 32'd1865
; 
32'd130710: dataIn1 = 32'd1866
; 
32'd130711: dataIn1 = 32'd1867
; 
32'd130712: dataIn1 = 32'd2046
; 
32'd130713: dataIn1 = 32'd1868
; 
32'd130714: dataIn1 = 32'd1871
; 
32'd130715: dataIn1 = 32'd2049
; 
32'd130716: dataIn1 = 32'd3036
; 
32'd130717: dataIn1 = 32'd3037
; 
32'd130718: dataIn1 = 32'd3039
; 
32'd130719: dataIn1 = 32'd3443
; 
32'd130720: dataIn1 = 32'd1869
; 
32'd130721: dataIn1 = 32'd3035
; 
32'd130722: dataIn1 = 32'd3037
; 
32'd130723: dataIn1 = 32'd3038
; 
32'd130724: dataIn1 = 32'd3418
; 
32'd130725: dataIn1 = 32'd3444
; 
32'd130726: dataIn1 = 32'd10260
; 
32'd130727: dataIn1 = 32'd213
; 
32'd130728: dataIn1 = 32'd796
; 
32'd130729: dataIn1 = 32'd979
; 
32'd130730: dataIn1 = 32'd1505
; 
32'd130731: dataIn1 = 32'd1870
; 
32'd130732: dataIn1 = 32'd1871
; 
32'd130733: dataIn1 = 32'd1879
; 
32'd130734: dataIn1 = 32'd2050
; 
32'd130735: dataIn1 = 32'd412
; 
32'd130736: dataIn1 = 32'd796
; 
32'd130737: dataIn1 = 32'd979
; 
32'd130738: dataIn1 = 32'd1504
; 
32'd130739: dataIn1 = 32'd1868
; 
32'd130740: dataIn1 = 32'd1870
; 
32'd130741: dataIn1 = 32'd1871
; 
32'd130742: dataIn1 = 32'd2049
; 
32'd130743: dataIn1 = 32'd3443
; 
32'd130744: dataIn1 = 32'd414
; 
32'd130745: dataIn1 = 32'd798
; 
32'd130746: dataIn1 = 32'd1507
; 
32'd130747: dataIn1 = 32'd1517
; 
32'd130748: dataIn1 = 32'd1872
; 
32'd130749: dataIn1 = 32'd2759
; 
32'd130750: dataIn1 = 32'd3040
; 
32'd130751: dataIn1 = 32'd415
; 
32'd130752: dataIn1 = 32'd801
; 
32'd130753: dataIn1 = 32'd983
; 
32'd130754: dataIn1 = 32'd1509
; 
32'd130755: dataIn1 = 32'd1873
; 
32'd130756: dataIn1 = 32'd1874
; 
32'd130757: dataIn1 = 32'd1875
; 
32'd130758: dataIn1 = 32'd2051
; 
32'd130759: dataIn1 = 32'd10273
; 
32'd130760: dataIn1 = 32'd10285
; 
32'd130761: dataIn1 = 32'd1873
; 
32'd130762: dataIn1 = 32'd1874
; 
32'd130763: dataIn1 = 32'd10260
; 
32'd130764: dataIn1 = 32'd10261
; 
32'd130765: dataIn1 = 32'd10262
; 
32'd130766: dataIn1 = 32'd10273
; 
32'd130767: dataIn1 = 32'd10285
; 
32'd130768: dataIn1 = 32'd415
; 
32'd130769: dataIn1 = 32'd803
; 
32'd130770: dataIn1 = 32'd982
; 
32'd130771: dataIn1 = 32'd1512
; 
32'd130772: dataIn1 = 32'd1873
; 
32'd130773: dataIn1 = 32'd1875
; 
32'd130774: dataIn1 = 32'd1876
; 
32'd130775: dataIn1 = 32'd2051
; 
32'd130776: dataIn1 = 32'd210
; 
32'd130777: dataIn1 = 32'd803
; 
32'd130778: dataIn1 = 32'd982
; 
32'd130779: dataIn1 = 32'd1511
; 
32'd130780: dataIn1 = 32'd1866
; 
32'd130781: dataIn1 = 32'd1875
; 
32'd130782: dataIn1 = 32'd1876
; 
32'd130783: dataIn1 = 32'd2047
; 
32'd130784: dataIn1 = 32'd214
; 
32'd130785: dataIn1 = 32'd810
; 
32'd130786: dataIn1 = 32'd985
; 
32'd130787: dataIn1 = 32'd1522
; 
32'd130788: dataIn1 = 32'd1877
; 
32'd130789: dataIn1 = 32'd1878
; 
32'd130790: dataIn1 = 32'd1881
; 
32'd130791: dataIn1 = 32'd2053
; 
32'd130792: dataIn1 = 32'd417
; 
32'd130793: dataIn1 = 32'd810
; 
32'd130794: dataIn1 = 32'd985
; 
32'd130795: dataIn1 = 32'd1521
; 
32'd130796: dataIn1 = 32'd1877
; 
32'd130797: dataIn1 = 32'd1878
; 
32'd130798: dataIn1 = 32'd1880
; 
32'd130799: dataIn1 = 32'd2052
; 
32'd130800: dataIn1 = 32'd213
; 
32'd130801: dataIn1 = 32'd812
; 
32'd130802: dataIn1 = 32'd984
; 
32'd130803: dataIn1 = 32'd1525
; 
32'd130804: dataIn1 = 32'd1870
; 
32'd130805: dataIn1 = 32'd1879
; 
32'd130806: dataIn1 = 32'd1880
; 
32'd130807: dataIn1 = 32'd2050
; 
32'd130808: dataIn1 = 32'd417
; 
32'd130809: dataIn1 = 32'd812
; 
32'd130810: dataIn1 = 32'd984
; 
32'd130811: dataIn1 = 32'd1524
; 
32'd130812: dataIn1 = 32'd1878
; 
32'd130813: dataIn1 = 32'd1879
; 
32'd130814: dataIn1 = 32'd1880
; 
32'd130815: dataIn1 = 32'd2052
; 
32'd130816: dataIn1 = 32'd214
; 
32'd130817: dataIn1 = 32'd816
; 
32'd130818: dataIn1 = 32'd987
; 
32'd130819: dataIn1 = 32'd1531
; 
32'd130820: dataIn1 = 32'd1877
; 
32'd130821: dataIn1 = 32'd1881
; 
32'd130822: dataIn1 = 32'd1882
; 
32'd130823: dataIn1 = 32'd2053
; 
32'd130824: dataIn1 = 32'd418
; 
32'd130825: dataIn1 = 32'd816
; 
32'd130826: dataIn1 = 32'd987
; 
32'd130827: dataIn1 = 32'd1530
; 
32'd130828: dataIn1 = 32'd1881
; 
32'd130829: dataIn1 = 32'd1882
; 
32'd130830: dataIn1 = 32'd1884
; 
32'd130831: dataIn1 = 32'd2054
; 
32'd130832: dataIn1 = 32'd216
; 
32'd130833: dataIn1 = 32'd818
; 
32'd130834: dataIn1 = 32'd986
; 
32'd130835: dataIn1 = 32'd1534
; 
32'd130836: dataIn1 = 32'd1883
; 
32'd130837: dataIn1 = 32'd1884
; 
32'd130838: dataIn1 = 32'd1892
; 
32'd130839: dataIn1 = 32'd2055
; 
32'd130840: dataIn1 = 32'd418
; 
32'd130841: dataIn1 = 32'd818
; 
32'd130842: dataIn1 = 32'd986
; 
32'd130843: dataIn1 = 32'd1533
; 
32'd130844: dataIn1 = 32'd1882
; 
32'd130845: dataIn1 = 32'd1883
; 
32'd130846: dataIn1 = 32'd1884
; 
32'd130847: dataIn1 = 32'd2054
; 
32'd130848: dataIn1 = 32'd419
; 
32'd130849: dataIn1 = 32'd822
; 
32'd130850: dataIn1 = 32'd989
; 
32'd130851: dataIn1 = 32'd1538
; 
32'd130852: dataIn1 = 32'd1885
; 
32'd130853: dataIn1 = 32'd1886
; 
32'd130854: dataIn1 = 32'd1888
; 
32'd130855: dataIn1 = 32'd2057
; 
32'd130856: dataIn1 = 32'd217
; 
32'd130857: dataIn1 = 32'd822
; 
32'd130858: dataIn1 = 32'd989
; 
32'd130859: dataIn1 = 32'd1537
; 
32'd130860: dataIn1 = 32'd1885
; 
32'd130861: dataIn1 = 32'd1886
; 
32'd130862: dataIn1 = 32'd1890
; 
32'd130863: dataIn1 = 32'd2056
; 
32'd130864: dataIn1 = 32'd219
; 
32'd130865: dataIn1 = 32'd823
; 
32'd130866: dataIn1 = 32'd988
; 
32'd130867: dataIn1 = 32'd1541
; 
32'd130868: dataIn1 = 32'd1887
; 
32'd130869: dataIn1 = 32'd1888
; 
32'd130870: dataIn1 = 32'd1895
; 
32'd130871: dataIn1 = 32'd2058
; 
32'd130872: dataIn1 = 32'd419
; 
32'd130873: dataIn1 = 32'd823
; 
32'd130874: dataIn1 = 32'd988
; 
32'd130875: dataIn1 = 32'd1540
; 
32'd130876: dataIn1 = 32'd1885
; 
32'd130877: dataIn1 = 32'd1887
; 
32'd130878: dataIn1 = 32'd1888
; 
32'd130879: dataIn1 = 32'd2057
; 
32'd130880: dataIn1 = 32'd420
; 
32'd130881: dataIn1 = 32'd827
; 
32'd130882: dataIn1 = 32'd991
; 
32'd130883: dataIn1 = 32'd1545
; 
32'd130884: dataIn1 = 32'd1889
; 
32'd130885: dataIn1 = 32'd1890
; 
32'd130886: dataIn1 = 32'd1891
; 
32'd130887: dataIn1 = 32'd2059
; 
32'd130888: dataIn1 = 32'd217
; 
32'd130889: dataIn1 = 32'd827
; 
32'd130890: dataIn1 = 32'd991
; 
32'd130891: dataIn1 = 32'd1544
; 
32'd130892: dataIn1 = 32'd1886
; 
32'd130893: dataIn1 = 32'd1889
; 
32'd130894: dataIn1 = 32'd1890
; 
32'd130895: dataIn1 = 32'd2056
; 
32'd130896: dataIn1 = 32'd420
; 
32'd130897: dataIn1 = 32'd829
; 
32'd130898: dataIn1 = 32'd990
; 
32'd130899: dataIn1 = 32'd1548
; 
32'd130900: dataIn1 = 32'd1889
; 
32'd130901: dataIn1 = 32'd1891
; 
32'd130902: dataIn1 = 32'd1892
; 
32'd130903: dataIn1 = 32'd2059
; 
32'd130904: dataIn1 = 32'd216
; 
32'd130905: dataIn1 = 32'd829
; 
32'd130906: dataIn1 = 32'd990
; 
32'd130907: dataIn1 = 32'd1547
; 
32'd130908: dataIn1 = 32'd1883
; 
32'd130909: dataIn1 = 32'd1891
; 
32'd130910: dataIn1 = 32'd1892
; 
32'd130911: dataIn1 = 32'd2055
; 
32'd130912: dataIn1 = 32'd220
; 
32'd130913: dataIn1 = 32'd834
; 
32'd130914: dataIn1 = 32'd993
; 
32'd130915: dataIn1 = 32'd1554
; 
32'd130916: dataIn1 = 32'd1893
; 
32'd130917: dataIn1 = 32'd1894
; 
32'd130918: dataIn1 = 32'd1897
; 
32'd130919: dataIn1 = 32'd2061
; 
32'd130920: dataIn1 = 32'd421
; 
32'd130921: dataIn1 = 32'd834
; 
32'd130922: dataIn1 = 32'd993
; 
32'd130923: dataIn1 = 32'd1553
; 
32'd130924: dataIn1 = 32'd1893
; 
32'd130925: dataIn1 = 32'd1894
; 
32'd130926: dataIn1 = 32'd1896
; 
32'd130927: dataIn1 = 32'd2060
; 
32'd130928: dataIn1 = 32'd219
; 
32'd130929: dataIn1 = 32'd836
; 
32'd130930: dataIn1 = 32'd992
; 
32'd130931: dataIn1 = 32'd1557
; 
32'd130932: dataIn1 = 32'd1887
; 
32'd130933: dataIn1 = 32'd1895
; 
32'd130934: dataIn1 = 32'd1896
; 
32'd130935: dataIn1 = 32'd2058
; 
32'd130936: dataIn1 = 32'd421
; 
32'd130937: dataIn1 = 32'd836
; 
32'd130938: dataIn1 = 32'd992
; 
32'd130939: dataIn1 = 32'd1556
; 
32'd130940: dataIn1 = 32'd1894
; 
32'd130941: dataIn1 = 32'd1895
; 
32'd130942: dataIn1 = 32'd1896
; 
32'd130943: dataIn1 = 32'd2060
; 
32'd130944: dataIn1 = 32'd220
; 
32'd130945: dataIn1 = 32'd840
; 
32'd130946: dataIn1 = 32'd995
; 
32'd130947: dataIn1 = 32'd1563
; 
32'd130948: dataIn1 = 32'd1893
; 
32'd130949: dataIn1 = 32'd1897
; 
32'd130950: dataIn1 = 32'd1898
; 
32'd130951: dataIn1 = 32'd2061
; 
32'd130952: dataIn1 = 32'd422
; 
32'd130953: dataIn1 = 32'd840
; 
32'd130954: dataIn1 = 32'd995
; 
32'd130955: dataIn1 = 32'd1562
; 
32'd130956: dataIn1 = 32'd1897
; 
32'd130957: dataIn1 = 32'd1898
; 
32'd130958: dataIn1 = 32'd1900
; 
32'd130959: dataIn1 = 32'd2062
; 
32'd130960: dataIn1 = 32'd222
; 
32'd130961: dataIn1 = 32'd842
; 
32'd130962: dataIn1 = 32'd994
; 
32'd130963: dataIn1 = 32'd1566
; 
32'd130964: dataIn1 = 32'd1899
; 
32'd130965: dataIn1 = 32'd1900
; 
32'd130966: dataIn1 = 32'd1908
; 
32'd130967: dataIn1 = 32'd2063
; 
32'd130968: dataIn1 = 32'd422
; 
32'd130969: dataIn1 = 32'd842
; 
32'd130970: dataIn1 = 32'd994
; 
32'd130971: dataIn1 = 32'd1565
; 
32'd130972: dataIn1 = 32'd1898
; 
32'd130973: dataIn1 = 32'd1899
; 
32'd130974: dataIn1 = 32'd1900
; 
32'd130975: dataIn1 = 32'd2062
; 
32'd130976: dataIn1 = 32'd423
; 
32'd130977: dataIn1 = 32'd846
; 
32'd130978: dataIn1 = 32'd997
; 
32'd130979: dataIn1 = 32'd1570
; 
32'd130980: dataIn1 = 32'd1901
; 
32'd130981: dataIn1 = 32'd1902
; 
32'd130982: dataIn1 = 32'd1904
; 
32'd130983: dataIn1 = 32'd2065
; 
32'd130984: dataIn1 = 32'd223
; 
32'd130985: dataIn1 = 32'd846
; 
32'd130986: dataIn1 = 32'd997
; 
32'd130987: dataIn1 = 32'd1569
; 
32'd130988: dataIn1 = 32'd1901
; 
32'd130989: dataIn1 = 32'd1902
; 
32'd130990: dataIn1 = 32'd1906
; 
32'd130991: dataIn1 = 32'd2064
; 
32'd130992: dataIn1 = 32'd225
; 
32'd130993: dataIn1 = 32'd847
; 
32'd130994: dataIn1 = 32'd996
; 
32'd130995: dataIn1 = 32'd1573
; 
32'd130996: dataIn1 = 32'd1903
; 
32'd130997: dataIn1 = 32'd1904
; 
32'd130998: dataIn1 = 32'd1911
; 
32'd130999: dataIn1 = 32'd2066
; 
32'd131000: dataIn1 = 32'd423
; 
32'd131001: dataIn1 = 32'd847
; 
32'd131002: dataIn1 = 32'd996
; 
32'd131003: dataIn1 = 32'd1572
; 
32'd131004: dataIn1 = 32'd1901
; 
32'd131005: dataIn1 = 32'd1903
; 
32'd131006: dataIn1 = 32'd1904
; 
32'd131007: dataIn1 = 32'd2065
; 
32'd131008: dataIn1 = 32'd424
; 
32'd131009: dataIn1 = 32'd851
; 
32'd131010: dataIn1 = 32'd999
; 
32'd131011: dataIn1 = 32'd1577
; 
32'd131012: dataIn1 = 32'd1905
; 
32'd131013: dataIn1 = 32'd1906
; 
32'd131014: dataIn1 = 32'd1907
; 
32'd131015: dataIn1 = 32'd2067
; 
32'd131016: dataIn1 = 32'd223
; 
32'd131017: dataIn1 = 32'd851
; 
32'd131018: dataIn1 = 32'd999
; 
32'd131019: dataIn1 = 32'd1576
; 
32'd131020: dataIn1 = 32'd1902
; 
32'd131021: dataIn1 = 32'd1905
; 
32'd131022: dataIn1 = 32'd1906
; 
32'd131023: dataIn1 = 32'd2064
; 
32'd131024: dataIn1 = 32'd424
; 
32'd131025: dataIn1 = 32'd853
; 
32'd131026: dataIn1 = 32'd998
; 
32'd131027: dataIn1 = 32'd1580
; 
32'd131028: dataIn1 = 32'd1905
; 
32'd131029: dataIn1 = 32'd1907
; 
32'd131030: dataIn1 = 32'd1908
; 
32'd131031: dataIn1 = 32'd2067
; 
32'd131032: dataIn1 = 32'd222
; 
32'd131033: dataIn1 = 32'd853
; 
32'd131034: dataIn1 = 32'd998
; 
32'd131035: dataIn1 = 32'd1579
; 
32'd131036: dataIn1 = 32'd1899
; 
32'd131037: dataIn1 = 32'd1907
; 
32'd131038: dataIn1 = 32'd1908
; 
32'd131039: dataIn1 = 32'd2063
; 
32'd131040: dataIn1 = 32'd226
; 
32'd131041: dataIn1 = 32'd858
; 
32'd131042: dataIn1 = 32'd1001
; 
32'd131043: dataIn1 = 32'd1586
; 
32'd131044: dataIn1 = 32'd1909
; 
32'd131045: dataIn1 = 32'd1910
; 
32'd131046: dataIn1 = 32'd1913
; 
32'd131047: dataIn1 = 32'd2069
; 
32'd131048: dataIn1 = 32'd425
; 
32'd131049: dataIn1 = 32'd858
; 
32'd131050: dataIn1 = 32'd1001
; 
32'd131051: dataIn1 = 32'd1585
; 
32'd131052: dataIn1 = 32'd1909
; 
32'd131053: dataIn1 = 32'd1910
; 
32'd131054: dataIn1 = 32'd1912
; 
32'd131055: dataIn1 = 32'd2068
; 
32'd131056: dataIn1 = 32'd225
; 
32'd131057: dataIn1 = 32'd860
; 
32'd131058: dataIn1 = 32'd1000
; 
32'd131059: dataIn1 = 32'd1589
; 
32'd131060: dataIn1 = 32'd1903
; 
32'd131061: dataIn1 = 32'd1911
; 
32'd131062: dataIn1 = 32'd1912
; 
32'd131063: dataIn1 = 32'd2066
; 
32'd131064: dataIn1 = 32'd425
; 
32'd131065: dataIn1 = 32'd860
; 
32'd131066: dataIn1 = 32'd1000
; 
32'd131067: dataIn1 = 32'd1588
; 
32'd131068: dataIn1 = 32'd1910
; 
32'd131069: dataIn1 = 32'd1911
; 
32'd131070: dataIn1 = 32'd1912
; 
32'd131071: dataIn1 = 32'd2068
; 
32'd131072: dataIn1 = 32'd226
; 
32'd131073: dataIn1 = 32'd864
; 
32'd131074: dataIn1 = 32'd1003
; 
32'd131075: dataIn1 = 32'd1595
; 
32'd131076: dataIn1 = 32'd1909
; 
32'd131077: dataIn1 = 32'd1913
; 
32'd131078: dataIn1 = 32'd1914
; 
32'd131079: dataIn1 = 32'd2069
; 
32'd131080: dataIn1 = 32'd426
; 
32'd131081: dataIn1 = 32'd864
; 
32'd131082: dataIn1 = 32'd1003
; 
32'd131083: dataIn1 = 32'd1594
; 
32'd131084: dataIn1 = 32'd1913
; 
32'd131085: dataIn1 = 32'd1914
; 
32'd131086: dataIn1 = 32'd1916
; 
32'd131087: dataIn1 = 32'd2070
; 
32'd131088: dataIn1 = 32'd228
; 
32'd131089: dataIn1 = 32'd866
; 
32'd131090: dataIn1 = 32'd1002
; 
32'd131091: dataIn1 = 32'd1598
; 
32'd131092: dataIn1 = 32'd1915
; 
32'd131093: dataIn1 = 32'd1916
; 
32'd131094: dataIn1 = 32'd1924
; 
32'd131095: dataIn1 = 32'd2071
; 
32'd131096: dataIn1 = 32'd426
; 
32'd131097: dataIn1 = 32'd866
; 
32'd131098: dataIn1 = 32'd1002
; 
32'd131099: dataIn1 = 32'd1597
; 
32'd131100: dataIn1 = 32'd1914
; 
32'd131101: dataIn1 = 32'd1915
; 
32'd131102: dataIn1 = 32'd1916
; 
32'd131103: dataIn1 = 32'd2070
; 
32'd131104: dataIn1 = 32'd427
; 
32'd131105: dataIn1 = 32'd870
; 
32'd131106: dataIn1 = 32'd1005
; 
32'd131107: dataIn1 = 32'd1602
; 
32'd131108: dataIn1 = 32'd1917
; 
32'd131109: dataIn1 = 32'd1918
; 
32'd131110: dataIn1 = 32'd1920
; 
32'd131111: dataIn1 = 32'd2073
; 
32'd131112: dataIn1 = 32'd229
; 
32'd131113: dataIn1 = 32'd870
; 
32'd131114: dataIn1 = 32'd1005
; 
32'd131115: dataIn1 = 32'd1601
; 
32'd131116: dataIn1 = 32'd1917
; 
32'd131117: dataIn1 = 32'd1918
; 
32'd131118: dataIn1 = 32'd1922
; 
32'd131119: dataIn1 = 32'd2072
; 
32'd131120: dataIn1 = 32'd231
; 
32'd131121: dataIn1 = 32'd871
; 
32'd131122: dataIn1 = 32'd1004
; 
32'd131123: dataIn1 = 32'd1605
; 
32'd131124: dataIn1 = 32'd1919
; 
32'd131125: dataIn1 = 32'd1920
; 
32'd131126: dataIn1 = 32'd1927
; 
32'd131127: dataIn1 = 32'd2074
; 
32'd131128: dataIn1 = 32'd427
; 
32'd131129: dataIn1 = 32'd871
; 
32'd131130: dataIn1 = 32'd1004
; 
32'd131131: dataIn1 = 32'd1604
; 
32'd131132: dataIn1 = 32'd1917
; 
32'd131133: dataIn1 = 32'd1919
; 
32'd131134: dataIn1 = 32'd1920
; 
32'd131135: dataIn1 = 32'd2073
; 
32'd131136: dataIn1 = 32'd428
; 
32'd131137: dataIn1 = 32'd875
; 
32'd131138: dataIn1 = 32'd1007
; 
32'd131139: dataIn1 = 32'd1609
; 
32'd131140: dataIn1 = 32'd1921
; 
32'd131141: dataIn1 = 32'd1922
; 
32'd131142: dataIn1 = 32'd1923
; 
32'd131143: dataIn1 = 32'd2075
; 
32'd131144: dataIn1 = 32'd229
; 
32'd131145: dataIn1 = 32'd875
; 
32'd131146: dataIn1 = 32'd1007
; 
32'd131147: dataIn1 = 32'd1608
; 
32'd131148: dataIn1 = 32'd1918
; 
32'd131149: dataIn1 = 32'd1921
; 
32'd131150: dataIn1 = 32'd1922
; 
32'd131151: dataIn1 = 32'd2072
; 
32'd131152: dataIn1 = 32'd428
; 
32'd131153: dataIn1 = 32'd877
; 
32'd131154: dataIn1 = 32'd1006
; 
32'd131155: dataIn1 = 32'd1612
; 
32'd131156: dataIn1 = 32'd1921
; 
32'd131157: dataIn1 = 32'd1923
; 
32'd131158: dataIn1 = 32'd1924
; 
32'd131159: dataIn1 = 32'd2075
; 
32'd131160: dataIn1 = 32'd228
; 
32'd131161: dataIn1 = 32'd877
; 
32'd131162: dataIn1 = 32'd1006
; 
32'd131163: dataIn1 = 32'd1611
; 
32'd131164: dataIn1 = 32'd1915
; 
32'd131165: dataIn1 = 32'd1923
; 
32'd131166: dataIn1 = 32'd1924
; 
32'd131167: dataIn1 = 32'd2071
; 
32'd131168: dataIn1 = 32'd232
; 
32'd131169: dataIn1 = 32'd882
; 
32'd131170: dataIn1 = 32'd1009
; 
32'd131171: dataIn1 = 32'd1618
; 
32'd131172: dataIn1 = 32'd1925
; 
32'd131173: dataIn1 = 32'd1926
; 
32'd131174: dataIn1 = 32'd1929
; 
32'd131175: dataIn1 = 32'd2077
; 
32'd131176: dataIn1 = 32'd429
; 
32'd131177: dataIn1 = 32'd882
; 
32'd131178: dataIn1 = 32'd1009
; 
32'd131179: dataIn1 = 32'd1617
; 
32'd131180: dataIn1 = 32'd1925
; 
32'd131181: dataIn1 = 32'd1926
; 
32'd131182: dataIn1 = 32'd1928
; 
32'd131183: dataIn1 = 32'd2076
; 
32'd131184: dataIn1 = 32'd231
; 
32'd131185: dataIn1 = 32'd884
; 
32'd131186: dataIn1 = 32'd1008
; 
32'd131187: dataIn1 = 32'd1621
; 
32'd131188: dataIn1 = 32'd1919
; 
32'd131189: dataIn1 = 32'd1927
; 
32'd131190: dataIn1 = 32'd1928
; 
32'd131191: dataIn1 = 32'd2074
; 
32'd131192: dataIn1 = 32'd429
; 
32'd131193: dataIn1 = 32'd884
; 
32'd131194: dataIn1 = 32'd1008
; 
32'd131195: dataIn1 = 32'd1620
; 
32'd131196: dataIn1 = 32'd1926
; 
32'd131197: dataIn1 = 32'd1927
; 
32'd131198: dataIn1 = 32'd1928
; 
32'd131199: dataIn1 = 32'd2076
; 
32'd131200: dataIn1 = 32'd232
; 
32'd131201: dataIn1 = 32'd888
; 
32'd131202: dataIn1 = 32'd1011
; 
32'd131203: dataIn1 = 32'd1627
; 
32'd131204: dataIn1 = 32'd1925
; 
32'd131205: dataIn1 = 32'd1929
; 
32'd131206: dataIn1 = 32'd1930
; 
32'd131207: dataIn1 = 32'd2077
; 
32'd131208: dataIn1 = 32'd430
; 
32'd131209: dataIn1 = 32'd888
; 
32'd131210: dataIn1 = 32'd1011
; 
32'd131211: dataIn1 = 32'd1626
; 
32'd131212: dataIn1 = 32'd1929
; 
32'd131213: dataIn1 = 32'd1930
; 
32'd131214: dataIn1 = 32'd1932
; 
32'd131215: dataIn1 = 32'd2078
; 
32'd131216: dataIn1 = 32'd234
; 
32'd131217: dataIn1 = 32'd890
; 
32'd131218: dataIn1 = 32'd1010
; 
32'd131219: dataIn1 = 32'd1630
; 
32'd131220: dataIn1 = 32'd1931
; 
32'd131221: dataIn1 = 32'd1932
; 
32'd131222: dataIn1 = 32'd1940
; 
32'd131223: dataIn1 = 32'd2079
; 
32'd131224: dataIn1 = 32'd430
; 
32'd131225: dataIn1 = 32'd890
; 
32'd131226: dataIn1 = 32'd1010
; 
32'd131227: dataIn1 = 32'd1629
; 
32'd131228: dataIn1 = 32'd1930
; 
32'd131229: dataIn1 = 32'd1931
; 
32'd131230: dataIn1 = 32'd1932
; 
32'd131231: dataIn1 = 32'd2078
; 
32'd131232: dataIn1 = 32'd431
; 
32'd131233: dataIn1 = 32'd894
; 
32'd131234: dataIn1 = 32'd1013
; 
32'd131235: dataIn1 = 32'd1634
; 
32'd131236: dataIn1 = 32'd1933
; 
32'd131237: dataIn1 = 32'd1934
; 
32'd131238: dataIn1 = 32'd1936
; 
32'd131239: dataIn1 = 32'd2081
; 
32'd131240: dataIn1 = 32'd235
; 
32'd131241: dataIn1 = 32'd894
; 
32'd131242: dataIn1 = 32'd1013
; 
32'd131243: dataIn1 = 32'd1633
; 
32'd131244: dataIn1 = 32'd1933
; 
32'd131245: dataIn1 = 32'd1934
; 
32'd131246: dataIn1 = 32'd1938
; 
32'd131247: dataIn1 = 32'd2080
; 
32'd131248: dataIn1 = 32'd237
; 
32'd131249: dataIn1 = 32'd895
; 
32'd131250: dataIn1 = 32'd1012
; 
32'd131251: dataIn1 = 32'd1637
; 
32'd131252: dataIn1 = 32'd1935
; 
32'd131253: dataIn1 = 32'd1936
; 
32'd131254: dataIn1 = 32'd1943
; 
32'd131255: dataIn1 = 32'd2082
; 
32'd131256: dataIn1 = 32'd431
; 
32'd131257: dataIn1 = 32'd895
; 
32'd131258: dataIn1 = 32'd1012
; 
32'd131259: dataIn1 = 32'd1636
; 
32'd131260: dataIn1 = 32'd1933
; 
32'd131261: dataIn1 = 32'd1935
; 
32'd131262: dataIn1 = 32'd1936
; 
32'd131263: dataIn1 = 32'd2081
; 
32'd131264: dataIn1 = 32'd432
; 
32'd131265: dataIn1 = 32'd899
; 
32'd131266: dataIn1 = 32'd1015
; 
32'd131267: dataIn1 = 32'd1641
; 
32'd131268: dataIn1 = 32'd1937
; 
32'd131269: dataIn1 = 32'd1938
; 
32'd131270: dataIn1 = 32'd1939
; 
32'd131271: dataIn1 = 32'd2083
; 
32'd131272: dataIn1 = 32'd235
; 
32'd131273: dataIn1 = 32'd899
; 
32'd131274: dataIn1 = 32'd1015
; 
32'd131275: dataIn1 = 32'd1640
; 
32'd131276: dataIn1 = 32'd1934
; 
32'd131277: dataIn1 = 32'd1937
; 
32'd131278: dataIn1 = 32'd1938
; 
32'd131279: dataIn1 = 32'd2080
; 
32'd131280: dataIn1 = 32'd432
; 
32'd131281: dataIn1 = 32'd901
; 
32'd131282: dataIn1 = 32'd1014
; 
32'd131283: dataIn1 = 32'd1644
; 
32'd131284: dataIn1 = 32'd1937
; 
32'd131285: dataIn1 = 32'd1939
; 
32'd131286: dataIn1 = 32'd1940
; 
32'd131287: dataIn1 = 32'd2083
; 
32'd131288: dataIn1 = 32'd234
; 
32'd131289: dataIn1 = 32'd901
; 
32'd131290: dataIn1 = 32'd1014
; 
32'd131291: dataIn1 = 32'd1643
; 
32'd131292: dataIn1 = 32'd1931
; 
32'd131293: dataIn1 = 32'd1939
; 
32'd131294: dataIn1 = 32'd1940
; 
32'd131295: dataIn1 = 32'd2079
; 
32'd131296: dataIn1 = 32'd238
; 
32'd131297: dataIn1 = 32'd906
; 
32'd131298: dataIn1 = 32'd1017
; 
32'd131299: dataIn1 = 32'd1650
; 
32'd131300: dataIn1 = 32'd1941
; 
32'd131301: dataIn1 = 32'd1942
; 
32'd131302: dataIn1 = 32'd1945
; 
32'd131303: dataIn1 = 32'd2085
; 
32'd131304: dataIn1 = 32'd433
; 
32'd131305: dataIn1 = 32'd906
; 
32'd131306: dataIn1 = 32'd1017
; 
32'd131307: dataIn1 = 32'd1649
; 
32'd131308: dataIn1 = 32'd1941
; 
32'd131309: dataIn1 = 32'd1942
; 
32'd131310: dataIn1 = 32'd1944
; 
32'd131311: dataIn1 = 32'd2084
; 
32'd131312: dataIn1 = 32'd237
; 
32'd131313: dataIn1 = 32'd908
; 
32'd131314: dataIn1 = 32'd1016
; 
32'd131315: dataIn1 = 32'd1653
; 
32'd131316: dataIn1 = 32'd1935
; 
32'd131317: dataIn1 = 32'd1943
; 
32'd131318: dataIn1 = 32'd1944
; 
32'd131319: dataIn1 = 32'd2082
; 
32'd131320: dataIn1 = 32'd433
; 
32'd131321: dataIn1 = 32'd908
; 
32'd131322: dataIn1 = 32'd1016
; 
32'd131323: dataIn1 = 32'd1652
; 
32'd131324: dataIn1 = 32'd1942
; 
32'd131325: dataIn1 = 32'd1943
; 
32'd131326: dataIn1 = 32'd1944
; 
32'd131327: dataIn1 = 32'd2084
; 
32'd131328: dataIn1 = 32'd238
; 
32'd131329: dataIn1 = 32'd912
; 
32'd131330: dataIn1 = 32'd1019
; 
32'd131331: dataIn1 = 32'd1659
; 
32'd131332: dataIn1 = 32'd1941
; 
32'd131333: dataIn1 = 32'd1945
; 
32'd131334: dataIn1 = 32'd1946
; 
32'd131335: dataIn1 = 32'd2085
; 
32'd131336: dataIn1 = 32'd434
; 
32'd131337: dataIn1 = 32'd912
; 
32'd131338: dataIn1 = 32'd1019
; 
32'd131339: dataIn1 = 32'd1658
; 
32'd131340: dataIn1 = 32'd1945
; 
32'd131341: dataIn1 = 32'd1946
; 
32'd131342: dataIn1 = 32'd1948
; 
32'd131343: dataIn1 = 32'd2086
; 
32'd131344: dataIn1 = 32'd240
; 
32'd131345: dataIn1 = 32'd914
; 
32'd131346: dataIn1 = 32'd1018
; 
32'd131347: dataIn1 = 32'd1662
; 
32'd131348: dataIn1 = 32'd1947
; 
32'd131349: dataIn1 = 32'd1948
; 
32'd131350: dataIn1 = 32'd1956
; 
32'd131351: dataIn1 = 32'd2087
; 
32'd131352: dataIn1 = 32'd434
; 
32'd131353: dataIn1 = 32'd914
; 
32'd131354: dataIn1 = 32'd1018
; 
32'd131355: dataIn1 = 32'd1661
; 
32'd131356: dataIn1 = 32'd1946
; 
32'd131357: dataIn1 = 32'd1947
; 
32'd131358: dataIn1 = 32'd1948
; 
32'd131359: dataIn1 = 32'd2086
; 
32'd131360: dataIn1 = 32'd435
; 
32'd131361: dataIn1 = 32'd918
; 
32'd131362: dataIn1 = 32'd1021
; 
32'd131363: dataIn1 = 32'd1666
; 
32'd131364: dataIn1 = 32'd1949
; 
32'd131365: dataIn1 = 32'd1950
; 
32'd131366: dataIn1 = 32'd1952
; 
32'd131367: dataIn1 = 32'd2089
; 
32'd131368: dataIn1 = 32'd241
; 
32'd131369: dataIn1 = 32'd918
; 
32'd131370: dataIn1 = 32'd1021
; 
32'd131371: dataIn1 = 32'd1665
; 
32'd131372: dataIn1 = 32'd1949
; 
32'd131373: dataIn1 = 32'd1950
; 
32'd131374: dataIn1 = 32'd1954
; 
32'd131375: dataIn1 = 32'd2088
; 
32'd131376: dataIn1 = 32'd243
; 
32'd131377: dataIn1 = 32'd919
; 
32'd131378: dataIn1 = 32'd1020
; 
32'd131379: dataIn1 = 32'd1669
; 
32'd131380: dataIn1 = 32'd1951
; 
32'd131381: dataIn1 = 32'd1952
; 
32'd131382: dataIn1 = 32'd1959
; 
32'd131383: dataIn1 = 32'd2090
; 
32'd131384: dataIn1 = 32'd435
; 
32'd131385: dataIn1 = 32'd919
; 
32'd131386: dataIn1 = 32'd1020
; 
32'd131387: dataIn1 = 32'd1668
; 
32'd131388: dataIn1 = 32'd1949
; 
32'd131389: dataIn1 = 32'd1951
; 
32'd131390: dataIn1 = 32'd1952
; 
32'd131391: dataIn1 = 32'd2089
; 
32'd131392: dataIn1 = 32'd436
; 
32'd131393: dataIn1 = 32'd923
; 
32'd131394: dataIn1 = 32'd1023
; 
32'd131395: dataIn1 = 32'd1673
; 
32'd131396: dataIn1 = 32'd1953
; 
32'd131397: dataIn1 = 32'd1954
; 
32'd131398: dataIn1 = 32'd1955
; 
32'd131399: dataIn1 = 32'd2091
; 
32'd131400: dataIn1 = 32'd241
; 
32'd131401: dataIn1 = 32'd923
; 
32'd131402: dataIn1 = 32'd1023
; 
32'd131403: dataIn1 = 32'd1672
; 
32'd131404: dataIn1 = 32'd1950
; 
32'd131405: dataIn1 = 32'd1953
; 
32'd131406: dataIn1 = 32'd1954
; 
32'd131407: dataIn1 = 32'd2088
; 
32'd131408: dataIn1 = 32'd436
; 
32'd131409: dataIn1 = 32'd925
; 
32'd131410: dataIn1 = 32'd1022
; 
32'd131411: dataIn1 = 32'd1676
; 
32'd131412: dataIn1 = 32'd1953
; 
32'd131413: dataIn1 = 32'd1955
; 
32'd131414: dataIn1 = 32'd1956
; 
32'd131415: dataIn1 = 32'd2091
; 
32'd131416: dataIn1 = 32'd240
; 
32'd131417: dataIn1 = 32'd925
; 
32'd131418: dataIn1 = 32'd1022
; 
32'd131419: dataIn1 = 32'd1675
; 
32'd131420: dataIn1 = 32'd1947
; 
32'd131421: dataIn1 = 32'd1955
; 
32'd131422: dataIn1 = 32'd1956
; 
32'd131423: dataIn1 = 32'd2087
; 
32'd131424: dataIn1 = 32'd244
; 
32'd131425: dataIn1 = 32'd930
; 
32'd131426: dataIn1 = 32'd1025
; 
32'd131427: dataIn1 = 32'd1682
; 
32'd131428: dataIn1 = 32'd1957
; 
32'd131429: dataIn1 = 32'd1958
; 
32'd131430: dataIn1 = 32'd1961
; 
32'd131431: dataIn1 = 32'd2093
; 
32'd131432: dataIn1 = 32'd437
; 
32'd131433: dataIn1 = 32'd930
; 
32'd131434: dataIn1 = 32'd1025
; 
32'd131435: dataIn1 = 32'd1681
; 
32'd131436: dataIn1 = 32'd1957
; 
32'd131437: dataIn1 = 32'd1958
; 
32'd131438: dataIn1 = 32'd1960
; 
32'd131439: dataIn1 = 32'd2092
; 
32'd131440: dataIn1 = 32'd243
; 
32'd131441: dataIn1 = 32'd932
; 
32'd131442: dataIn1 = 32'd1024
; 
32'd131443: dataIn1 = 32'd1685
; 
32'd131444: dataIn1 = 32'd1951
; 
32'd131445: dataIn1 = 32'd1959
; 
32'd131446: dataIn1 = 32'd1960
; 
32'd131447: dataIn1 = 32'd2090
; 
32'd131448: dataIn1 = 32'd437
; 
32'd131449: dataIn1 = 32'd932
; 
32'd131450: dataIn1 = 32'd1024
; 
32'd131451: dataIn1 = 32'd1684
; 
32'd131452: dataIn1 = 32'd1958
; 
32'd131453: dataIn1 = 32'd1959
; 
32'd131454: dataIn1 = 32'd1960
; 
32'd131455: dataIn1 = 32'd2092
; 
32'd131456: dataIn1 = 32'd244
; 
32'd131457: dataIn1 = 32'd936
; 
32'd131458: dataIn1 = 32'd1027
; 
32'd131459: dataIn1 = 32'd1691
; 
32'd131460: dataIn1 = 32'd1957
; 
32'd131461: dataIn1 = 32'd1961
; 
32'd131462: dataIn1 = 32'd1962
; 
32'd131463: dataIn1 = 32'd2093
; 
32'd131464: dataIn1 = 32'd438
; 
32'd131465: dataIn1 = 32'd936
; 
32'd131466: dataIn1 = 32'd1027
; 
32'd131467: dataIn1 = 32'd1690
; 
32'd131468: dataIn1 = 32'd1961
; 
32'd131469: dataIn1 = 32'd1962
; 
32'd131470: dataIn1 = 32'd1964
; 
32'd131471: dataIn1 = 32'd2094
; 
32'd131472: dataIn1 = 32'd246
; 
32'd131473: dataIn1 = 32'd938
; 
32'd131474: dataIn1 = 32'd1026
; 
32'd131475: dataIn1 = 32'd1694
; 
32'd131476: dataIn1 = 32'd1963
; 
32'd131477: dataIn1 = 32'd1964
; 
32'd131478: dataIn1 = 32'd1972
; 
32'd131479: dataIn1 = 32'd2095
; 
32'd131480: dataIn1 = 32'd438
; 
32'd131481: dataIn1 = 32'd938
; 
32'd131482: dataIn1 = 32'd1026
; 
32'd131483: dataIn1 = 32'd1693
; 
32'd131484: dataIn1 = 32'd1962
; 
32'd131485: dataIn1 = 32'd1963
; 
32'd131486: dataIn1 = 32'd1964
; 
32'd131487: dataIn1 = 32'd2094
; 
32'd131488: dataIn1 = 32'd439
; 
32'd131489: dataIn1 = 32'd1029
; 
32'd131490: dataIn1 = 32'd1698
; 
32'd131491: dataIn1 = 32'd1700
; 
32'd131492: dataIn1 = 32'd1965
; 
32'd131493: dataIn1 = 32'd1966
; 
32'd131494: dataIn1 = 32'd1968
; 
32'd131495: dataIn1 = 32'd2097
; 
32'd131496: dataIn1 = 32'd942
; 
32'd131497: dataIn1 = 32'd1029
; 
32'd131498: dataIn1 = 32'd1697
; 
32'd131499: dataIn1 = 32'd1698
; 
32'd131500: dataIn1 = 32'd1965
; 
32'd131501: dataIn1 = 32'd1966
; 
32'd131502: dataIn1 = 32'd1970
; 
32'd131503: dataIn1 = 32'd2096
; 
32'd131504: dataIn1 = 32'd249
; 
32'd131505: dataIn1 = 32'd1028
; 
32'd131506: dataIn1 = 32'd1701
; 
32'd131507: dataIn1 = 32'd1717
; 
32'd131508: dataIn1 = 32'd1967
; 
32'd131509: dataIn1 = 32'd1968
; 
32'd131510: dataIn1 = 32'd1975
; 
32'd131511: dataIn1 = 32'd2098
; 
32'd131512: dataIn1 = 32'd943
; 
32'd131513: dataIn1 = 32'd1028
; 
32'd131514: dataIn1 = 32'd1700
; 
32'd131515: dataIn1 = 32'd1701
; 
32'd131516: dataIn1 = 32'd1965
; 
32'd131517: dataIn1 = 32'd1967
; 
32'd131518: dataIn1 = 32'd1968
; 
32'd131519: dataIn1 = 32'd2097
; 
32'd131520: dataIn1 = 32'd947
; 
32'd131521: dataIn1 = 32'd1031
; 
32'd131522: dataIn1 = 32'd1704
; 
32'd131523: dataIn1 = 32'd1705
; 
32'd131524: dataIn1 = 32'd1969
; 
32'd131525: dataIn1 = 32'd1970
; 
32'd131526: dataIn1 = 32'd1971
; 
32'd131527: dataIn1 = 32'd2099
; 
32'd131528: dataIn1 = 32'd247
; 
32'd131529: dataIn1 = 32'd1031
; 
32'd131530: dataIn1 = 32'd1697
; 
32'd131531: dataIn1 = 32'd1704
; 
32'd131532: dataIn1 = 32'd1966
; 
32'd131533: dataIn1 = 32'd1969
; 
32'd131534: dataIn1 = 32'd1970
; 
32'd131535: dataIn1 = 32'd2096
; 
32'd131536: dataIn1 = 32'd440
; 
32'd131537: dataIn1 = 32'd1030
; 
32'd131538: dataIn1 = 32'd1705
; 
32'd131539: dataIn1 = 32'd1708
; 
32'd131540: dataIn1 = 32'd1969
; 
32'd131541: dataIn1 = 32'd1971
; 
32'd131542: dataIn1 = 32'd1972
; 
32'd131543: dataIn1 = 32'd2099
; 
32'd131544: dataIn1 = 32'd246
; 
32'd131545: dataIn1 = 32'd949
; 
32'd131546: dataIn1 = 32'd1030
; 
32'd131547: dataIn1 = 32'd1707
; 
32'd131548: dataIn1 = 32'd1708
; 
32'd131549: dataIn1 = 32'd1963
; 
32'd131550: dataIn1 = 32'd1971
; 
32'd131551: dataIn1 = 32'd1972
; 
32'd131552: dataIn1 = 32'd2095
; 
32'd131553: dataIn1 = 32'd250
; 
32'd131554: dataIn1 = 32'd1033
; 
32'd131555: dataIn1 = 32'd1714
; 
32'd131556: dataIn1 = 32'd1973
; 
32'd131557: dataIn1 = 32'd1974
; 
32'd131558: dataIn1 = 32'd954
; 
32'd131559: dataIn1 = 32'd1033
; 
32'd131560: dataIn1 = 32'd1713
; 
32'd131561: dataIn1 = 32'd1714
; 
32'd131562: dataIn1 = 32'd1973
; 
32'd131563: dataIn1 = 32'd1974
; 
32'd131564: dataIn1 = 32'd1976
; 
32'd131565: dataIn1 = 32'd2100
; 
32'd131566: dataIn1 = 32'd956
; 
32'd131567: dataIn1 = 32'd1032
; 
32'd131568: dataIn1 = 32'd1716
; 
32'd131569: dataIn1 = 32'd1717
; 
32'd131570: dataIn1 = 32'd1967
; 
32'd131571: dataIn1 = 32'd1975
; 
32'd131572: dataIn1 = 32'd1976
; 
32'd131573: dataIn1 = 32'd2098
; 
32'd131574: dataIn1 = 32'd441
; 
32'd131575: dataIn1 = 32'd1032
; 
32'd131576: dataIn1 = 32'd1713
; 
32'd131577: dataIn1 = 32'd1716
; 
32'd131578: dataIn1 = 32'd1974
; 
32'd131579: dataIn1 = 32'd1975
; 
32'd131580: dataIn1 = 32'd1976
; 
32'd131581: dataIn1 = 32'd2100
; 
32'd131582: dataIn1 = 32'd1977
; 
32'd131583: dataIn1 = 32'd3041
; 
32'd131584: dataIn1 = 32'd3043
; 
32'd131585: dataIn1 = 32'd3044
; 
32'd131586: dataIn1 = 32'd3047
; 
32'd131587: dataIn1 = 32'd3998
; 
32'd131588: dataIn1 = 32'd4000
; 
32'd131589: dataIn1 = 32'd1978
; 
32'd131590: dataIn1 = 32'd3048
; 
32'd131591: dataIn1 = 32'd3049
; 
32'd131592: dataIn1 = 32'd3051
; 
32'd131593: dataIn1 = 32'd3052
; 
32'd131594: dataIn1 = 32'd3995
; 
32'd131595: dataIn1 = 32'd3996
; 
32'd131596: dataIn1 = 32'd1979
; 
32'd131597: dataIn1 = 32'd3056
; 
32'd131598: dataIn1 = 32'd3057
; 
32'd131599: dataIn1 = 32'd3060
; 
32'd131600: dataIn1 = 32'd3061
; 
32'd131601: dataIn1 = 32'd4024
; 
32'd131602: dataIn1 = 32'd4025
; 
32'd131603: dataIn1 = 32'd1980
; 
32'd131604: dataIn1 = 32'd3062
; 
32'd131605: dataIn1 = 32'd3063
; 
32'd131606: dataIn1 = 32'd3065
; 
32'd131607: dataIn1 = 32'd3066
; 
32'd131608: dataIn1 = 32'd4019
; 
32'd131609: dataIn1 = 32'd4020
; 
32'd131610: dataIn1 = 32'd1981
; 
32'd131611: dataIn1 = 32'd3069
; 
32'd131612: dataIn1 = 32'd3070
; 
32'd131613: dataIn1 = 32'd3072
; 
32'd131614: dataIn1 = 32'd3073
; 
32'd131615: dataIn1 = 32'd4043
; 
32'd131616: dataIn1 = 32'd4044
; 
32'd131617: dataIn1 = 32'd1982
; 
32'd131618: dataIn1 = 32'd3077
; 
32'd131619: dataIn1 = 32'd3078
; 
32'd131620: dataIn1 = 32'd3081
; 
32'd131621: dataIn1 = 32'd3082
; 
32'd131622: dataIn1 = 32'd4047
; 
32'd131623: dataIn1 = 32'd4048
; 
32'd131624: dataIn1 = 32'd1983
; 
32'd131625: dataIn1 = 32'd3083
; 
32'd131626: dataIn1 = 32'd3085
; 
32'd131627: dataIn1 = 32'd3086
; 
32'd131628: dataIn1 = 32'd3089
; 
32'd131629: dataIn1 = 32'd4094
; 
32'd131630: dataIn1 = 32'd4096
; 
32'd131631: dataIn1 = 32'd1984
; 
32'd131632: dataIn1 = 32'd3090
; 
32'd131633: dataIn1 = 32'd3091
; 
32'd131634: dataIn1 = 32'd3093
; 
32'd131635: dataIn1 = 32'd3094
; 
32'd131636: dataIn1 = 32'd4091
; 
32'd131637: dataIn1 = 32'd4092
; 
32'd131638: dataIn1 = 32'd1985
; 
32'd131639: dataIn1 = 32'd3098
; 
32'd131640: dataIn1 = 32'd3099
; 
32'd131641: dataIn1 = 32'd3102
; 
32'd131642: dataIn1 = 32'd3103
; 
32'd131643: dataIn1 = 32'd4071
; 
32'd131644: dataIn1 = 32'd4072
; 
32'd131645: dataIn1 = 32'd1986
; 
32'd131646: dataIn1 = 32'd3104
; 
32'd131647: dataIn1 = 32'd3106
; 
32'd131648: dataIn1 = 32'd3107
; 
32'd131649: dataIn1 = 32'd3110
; 
32'd131650: dataIn1 = 32'd4067
; 
32'd131651: dataIn1 = 32'd4069
; 
32'd131652: dataIn1 = 32'd1987
; 
32'd131653: dataIn1 = 32'd3112
; 
32'd131654: dataIn1 = 32'd3113
; 
32'd131655: dataIn1 = 32'd3116
; 
32'd131656: dataIn1 = 32'd3117
; 
32'd131657: dataIn1 = 32'd4120
; 
32'd131658: dataIn1 = 32'd4121
; 
32'd131659: dataIn1 = 32'd1988
; 
32'd131660: dataIn1 = 32'd3118
; 
32'd131661: dataIn1 = 32'd3119
; 
32'd131662: dataIn1 = 32'd3121
; 
32'd131663: dataIn1 = 32'd3122
; 
32'd131664: dataIn1 = 32'd4115
; 
32'd131665: dataIn1 = 32'd4116
; 
32'd131666: dataIn1 = 32'd1989
; 
32'd131667: dataIn1 = 32'd3125
; 
32'd131668: dataIn1 = 32'd3126
; 
32'd131669: dataIn1 = 32'd3128
; 
32'd131670: dataIn1 = 32'd3129
; 
32'd131671: dataIn1 = 32'd4139
; 
32'd131672: dataIn1 = 32'd4140
; 
32'd131673: dataIn1 = 32'd1990
; 
32'd131674: dataIn1 = 32'd3133
; 
32'd131675: dataIn1 = 32'd3134
; 
32'd131676: dataIn1 = 32'd3137
; 
32'd131677: dataIn1 = 32'd3138
; 
32'd131678: dataIn1 = 32'd4143
; 
32'd131679: dataIn1 = 32'd4144
; 
32'd131680: dataIn1 = 32'd1991
; 
32'd131681: dataIn1 = 32'd3139
; 
32'd131682: dataIn1 = 32'd3141
; 
32'd131683: dataIn1 = 32'd3142
; 
32'd131684: dataIn1 = 32'd3145
; 
32'd131685: dataIn1 = 32'd4190
; 
32'd131686: dataIn1 = 32'd4192
; 
32'd131687: dataIn1 = 32'd1992
; 
32'd131688: dataIn1 = 32'd3146
; 
32'd131689: dataIn1 = 32'd3147
; 
32'd131690: dataIn1 = 32'd3149
; 
32'd131691: dataIn1 = 32'd3150
; 
32'd131692: dataIn1 = 32'd4187
; 
32'd131693: dataIn1 = 32'd4188
; 
32'd131694: dataIn1 = 32'd1993
; 
32'd131695: dataIn1 = 32'd3154
; 
32'd131696: dataIn1 = 32'd3155
; 
32'd131697: dataIn1 = 32'd3158
; 
32'd131698: dataIn1 = 32'd3159
; 
32'd131699: dataIn1 = 32'd4167
; 
32'd131700: dataIn1 = 32'd4168
; 
32'd131701: dataIn1 = 32'd1994
; 
32'd131702: dataIn1 = 32'd3160
; 
32'd131703: dataIn1 = 32'd3162
; 
32'd131704: dataIn1 = 32'd3163
; 
32'd131705: dataIn1 = 32'd3166
; 
32'd131706: dataIn1 = 32'd4163
; 
32'd131707: dataIn1 = 32'd4165
; 
32'd131708: dataIn1 = 32'd1995
; 
32'd131709: dataIn1 = 32'd3168
; 
32'd131710: dataIn1 = 32'd3169
; 
32'd131711: dataIn1 = 32'd3172
; 
32'd131712: dataIn1 = 32'd3173
; 
32'd131713: dataIn1 = 32'd4216
; 
32'd131714: dataIn1 = 32'd4217
; 
32'd131715: dataIn1 = 32'd1996
; 
32'd131716: dataIn1 = 32'd3174
; 
32'd131717: dataIn1 = 32'd3175
; 
32'd131718: dataIn1 = 32'd3177
; 
32'd131719: dataIn1 = 32'd3178
; 
32'd131720: dataIn1 = 32'd4211
; 
32'd131721: dataIn1 = 32'd4212
; 
32'd131722: dataIn1 = 32'd1997
; 
32'd131723: dataIn1 = 32'd3181
; 
32'd131724: dataIn1 = 32'd3182
; 
32'd131725: dataIn1 = 32'd3184
; 
32'd131726: dataIn1 = 32'd3185
; 
32'd131727: dataIn1 = 32'd4235
; 
32'd131728: dataIn1 = 32'd4236
; 
32'd131729: dataIn1 = 32'd1998
; 
32'd131730: dataIn1 = 32'd3189
; 
32'd131731: dataIn1 = 32'd3190
; 
32'd131732: dataIn1 = 32'd3193
; 
32'd131733: dataIn1 = 32'd3194
; 
32'd131734: dataIn1 = 32'd4239
; 
32'd131735: dataIn1 = 32'd4240
; 
32'd131736: dataIn1 = 32'd1999
; 
32'd131737: dataIn1 = 32'd3195
; 
32'd131738: dataIn1 = 32'd3197
; 
32'd131739: dataIn1 = 32'd3198
; 
32'd131740: dataIn1 = 32'd3201
; 
32'd131741: dataIn1 = 32'd4286
; 
32'd131742: dataIn1 = 32'd4288
; 
32'd131743: dataIn1 = 32'd2000
; 
32'd131744: dataIn1 = 32'd3202
; 
32'd131745: dataIn1 = 32'd3203
; 
32'd131746: dataIn1 = 32'd3205
; 
32'd131747: dataIn1 = 32'd3206
; 
32'd131748: dataIn1 = 32'd4283
; 
32'd131749: dataIn1 = 32'd4284
; 
32'd131750: dataIn1 = 32'd2001
; 
32'd131751: dataIn1 = 32'd3210
; 
32'd131752: dataIn1 = 32'd3211
; 
32'd131753: dataIn1 = 32'd3214
; 
32'd131754: dataIn1 = 32'd3215
; 
32'd131755: dataIn1 = 32'd4263
; 
32'd131756: dataIn1 = 32'd4264
; 
32'd131757: dataIn1 = 32'd2002
; 
32'd131758: dataIn1 = 32'd3216
; 
32'd131759: dataIn1 = 32'd3218
; 
32'd131760: dataIn1 = 32'd3219
; 
32'd131761: dataIn1 = 32'd3222
; 
32'd131762: dataIn1 = 32'd4259
; 
32'd131763: dataIn1 = 32'd4261
; 
32'd131764: dataIn1 = 32'd2003
; 
32'd131765: dataIn1 = 32'd3224
; 
32'd131766: dataIn1 = 32'd3225
; 
32'd131767: dataIn1 = 32'd3228
; 
32'd131768: dataIn1 = 32'd3229
; 
32'd131769: dataIn1 = 32'd4312
; 
32'd131770: dataIn1 = 32'd4313
; 
32'd131771: dataIn1 = 32'd2004
; 
32'd131772: dataIn1 = 32'd3230
; 
32'd131773: dataIn1 = 32'd3231
; 
32'd131774: dataIn1 = 32'd3233
; 
32'd131775: dataIn1 = 32'd3234
; 
32'd131776: dataIn1 = 32'd4307
; 
32'd131777: dataIn1 = 32'd4308
; 
32'd131778: dataIn1 = 32'd2005
; 
32'd131779: dataIn1 = 32'd3237
; 
32'd131780: dataIn1 = 32'd3238
; 
32'd131781: dataIn1 = 32'd3240
; 
32'd131782: dataIn1 = 32'd3241
; 
32'd131783: dataIn1 = 32'd4331
; 
32'd131784: dataIn1 = 32'd4332
; 
32'd131785: dataIn1 = 32'd2006
; 
32'd131786: dataIn1 = 32'd3245
; 
32'd131787: dataIn1 = 32'd3246
; 
32'd131788: dataIn1 = 32'd3249
; 
32'd131789: dataIn1 = 32'd3250
; 
32'd131790: dataIn1 = 32'd4335
; 
32'd131791: dataIn1 = 32'd4336
; 
32'd131792: dataIn1 = 32'd2007
; 
32'd131793: dataIn1 = 32'd3251
; 
32'd131794: dataIn1 = 32'd3253
; 
32'd131795: dataIn1 = 32'd3254
; 
32'd131796: dataIn1 = 32'd3257
; 
32'd131797: dataIn1 = 32'd4382
; 
32'd131798: dataIn1 = 32'd4384
; 
32'd131799: dataIn1 = 32'd2008
; 
32'd131800: dataIn1 = 32'd3258
; 
32'd131801: dataIn1 = 32'd3259
; 
32'd131802: dataIn1 = 32'd3261
; 
32'd131803: dataIn1 = 32'd3262
; 
32'd131804: dataIn1 = 32'd4379
; 
32'd131805: dataIn1 = 32'd4380
; 
32'd131806: dataIn1 = 32'd2009
; 
32'd131807: dataIn1 = 32'd3266
; 
32'd131808: dataIn1 = 32'd3267
; 
32'd131809: dataIn1 = 32'd3270
; 
32'd131810: dataIn1 = 32'd3271
; 
32'd131811: dataIn1 = 32'd4359
; 
32'd131812: dataIn1 = 32'd4360
; 
32'd131813: dataIn1 = 32'd2010
; 
32'd131814: dataIn1 = 32'd3272
; 
32'd131815: dataIn1 = 32'd3274
; 
32'd131816: dataIn1 = 32'd3275
; 
32'd131817: dataIn1 = 32'd3278
; 
32'd131818: dataIn1 = 32'd4355
; 
32'd131819: dataIn1 = 32'd4357
; 
32'd131820: dataIn1 = 32'd2011
; 
32'd131821: dataIn1 = 32'd3280
; 
32'd131822: dataIn1 = 32'd3281
; 
32'd131823: dataIn1 = 32'd3284
; 
32'd131824: dataIn1 = 32'd3285
; 
32'd131825: dataIn1 = 32'd4408
; 
32'd131826: dataIn1 = 32'd4409
; 
32'd131827: dataIn1 = 32'd2012
; 
32'd131828: dataIn1 = 32'd3286
; 
32'd131829: dataIn1 = 32'd3287
; 
32'd131830: dataIn1 = 32'd3289
; 
32'd131831: dataIn1 = 32'd3290
; 
32'd131832: dataIn1 = 32'd4403
; 
32'd131833: dataIn1 = 32'd4404
; 
32'd131834: dataIn1 = 32'd2013
; 
32'd131835: dataIn1 = 32'd3293
; 
32'd131836: dataIn1 = 32'd3294
; 
32'd131837: dataIn1 = 32'd3296
; 
32'd131838: dataIn1 = 32'd3297
; 
32'd131839: dataIn1 = 32'd4427
; 
32'd131840: dataIn1 = 32'd4428
; 
32'd131841: dataIn1 = 32'd2014
; 
32'd131842: dataIn1 = 32'd3301
; 
32'd131843: dataIn1 = 32'd3302
; 
32'd131844: dataIn1 = 32'd3305
; 
32'd131845: dataIn1 = 32'd3306
; 
32'd131846: dataIn1 = 32'd4431
; 
32'd131847: dataIn1 = 32'd4432
; 
32'd131848: dataIn1 = 32'd2015
; 
32'd131849: dataIn1 = 32'd3307
; 
32'd131850: dataIn1 = 32'd3309
; 
32'd131851: dataIn1 = 32'd3310
; 
32'd131852: dataIn1 = 32'd3313
; 
32'd131853: dataIn1 = 32'd4478
; 
32'd131854: dataIn1 = 32'd4480
; 
32'd131855: dataIn1 = 32'd2016
; 
32'd131856: dataIn1 = 32'd3314
; 
32'd131857: dataIn1 = 32'd3315
; 
32'd131858: dataIn1 = 32'd3317
; 
32'd131859: dataIn1 = 32'd3318
; 
32'd131860: dataIn1 = 32'd4475
; 
32'd131861: dataIn1 = 32'd4476
; 
32'd131862: dataIn1 = 32'd2017
; 
32'd131863: dataIn1 = 32'd3322
; 
32'd131864: dataIn1 = 32'd3323
; 
32'd131865: dataIn1 = 32'd3326
; 
32'd131866: dataIn1 = 32'd3327
; 
32'd131867: dataIn1 = 32'd4455
; 
32'd131868: dataIn1 = 32'd4456
; 
32'd131869: dataIn1 = 32'd2018
; 
32'd131870: dataIn1 = 32'd3328
; 
32'd131871: dataIn1 = 32'd3330
; 
32'd131872: dataIn1 = 32'd3331
; 
32'd131873: dataIn1 = 32'd3334
; 
32'd131874: dataIn1 = 32'd4451
; 
32'd131875: dataIn1 = 32'd4453
; 
32'd131876: dataIn1 = 32'd2019
; 
32'd131877: dataIn1 = 32'd3336
; 
32'd131878: dataIn1 = 32'd3337
; 
32'd131879: dataIn1 = 32'd3340
; 
32'd131880: dataIn1 = 32'd3341
; 
32'd131881: dataIn1 = 32'd4504
; 
32'd131882: dataIn1 = 32'd4505
; 
32'd131883: dataIn1 = 32'd2020
; 
32'd131884: dataIn1 = 32'd3342
; 
32'd131885: dataIn1 = 32'd3343
; 
32'd131886: dataIn1 = 32'd3345
; 
32'd131887: dataIn1 = 32'd3346
; 
32'd131888: dataIn1 = 32'd4499
; 
32'd131889: dataIn1 = 32'd4500
; 
32'd131890: dataIn1 = 32'd2021
; 
32'd131891: dataIn1 = 32'd3349
; 
32'd131892: dataIn1 = 32'd3350
; 
32'd131893: dataIn1 = 32'd3352
; 
32'd131894: dataIn1 = 32'd3353
; 
32'd131895: dataIn1 = 32'd4523
; 
32'd131896: dataIn1 = 32'd4524
; 
32'd131897: dataIn1 = 32'd2022
; 
32'd131898: dataIn1 = 32'd3357
; 
32'd131899: dataIn1 = 32'd3358
; 
32'd131900: dataIn1 = 32'd3361
; 
32'd131901: dataIn1 = 32'd3362
; 
32'd131902: dataIn1 = 32'd4527
; 
32'd131903: dataIn1 = 32'd4528
; 
32'd131904: dataIn1 = 32'd2023
; 
32'd131905: dataIn1 = 32'd3363
; 
32'd131906: dataIn1 = 32'd3365
; 
32'd131907: dataIn1 = 32'd3366
; 
32'd131908: dataIn1 = 32'd3369
; 
32'd131909: dataIn1 = 32'd4574
; 
32'd131910: dataIn1 = 32'd4576
; 
32'd131911: dataIn1 = 32'd2024
; 
32'd131912: dataIn1 = 32'd3370
; 
32'd131913: dataIn1 = 32'd3371
; 
32'd131914: dataIn1 = 32'd3373
; 
32'd131915: dataIn1 = 32'd3374
; 
32'd131916: dataIn1 = 32'd4571
; 
32'd131917: dataIn1 = 32'd4572
; 
32'd131918: dataIn1 = 32'd2025
; 
32'd131919: dataIn1 = 32'd3378
; 
32'd131920: dataIn1 = 32'd3379
; 
32'd131921: dataIn1 = 32'd3382
; 
32'd131922: dataIn1 = 32'd3383
; 
32'd131923: dataIn1 = 32'd4551
; 
32'd131924: dataIn1 = 32'd4552
; 
32'd131925: dataIn1 = 32'd2026
; 
32'd131926: dataIn1 = 32'd3384
; 
32'd131927: dataIn1 = 32'd3386
; 
32'd131928: dataIn1 = 32'd3387
; 
32'd131929: dataIn1 = 32'd3390
; 
32'd131930: dataIn1 = 32'd4547
; 
32'd131931: dataIn1 = 32'd4549
; 
32'd131932: dataIn1 = 32'd2027
; 
32'd131933: dataIn1 = 32'd3392
; 
32'd131934: dataIn1 = 32'd3393
; 
32'd131935: dataIn1 = 32'd3396
; 
32'd131936: dataIn1 = 32'd3397
; 
32'd131937: dataIn1 = 32'd4600
; 
32'd131938: dataIn1 = 32'd4601
; 
32'd131939: dataIn1 = 32'd2028
; 
32'd131940: dataIn1 = 32'd3398
; 
32'd131941: dataIn1 = 32'd3399
; 
32'd131942: dataIn1 = 32'd3401
; 
32'd131943: dataIn1 = 32'd3402
; 
32'd131944: dataIn1 = 32'd4595
; 
32'd131945: dataIn1 = 32'd4596
; 
32'd131946: dataIn1 = 32'd195
; 
32'd131947: dataIn1 = 32'd962
; 
32'd131948: dataIn1 = 32'd964
; 
32'd131949: dataIn1 = 32'd1034
; 
32'd131950: dataIn1 = 32'd1830
; 
32'd131951: dataIn1 = 32'd1834
; 
32'd131952: dataIn1 = 32'd2029
; 
32'd131953: dataIn1 = 32'd195
; 
32'd131954: dataIn1 = 32'd961
; 
32'd131955: dataIn1 = 32'd962
; 
32'd131956: dataIn1 = 32'd1035
; 
32'd131957: dataIn1 = 32'd1829
; 
32'd131958: dataIn1 = 32'd1832
; 
32'd131959: dataIn1 = 32'd2030
; 
32'd131960: dataIn1 = 32'd122
; 
32'd131961: dataIn1 = 32'd961
; 
32'd131962: dataIn1 = 32'd965
; 
32'd131963: dataIn1 = 32'd1035
; 
32'd131964: dataIn1 = 32'd1831
; 
32'd131965: dataIn1 = 32'd1839
; 
32'd131966: dataIn1 = 32'd2031
; 
32'd131967: dataIn1 = 32'd123
; 
32'd131968: dataIn1 = 32'd963
; 
32'd131969: dataIn1 = 32'd964
; 
32'd131970: dataIn1 = 32'd1034
; 
32'd131971: dataIn1 = 32'd1833
; 
32'd131972: dataIn1 = 32'd1835
; 
32'd131973: dataIn1 = 32'd2032
; 
32'd131974: dataIn1 = 32'd122
; 
32'd131975: dataIn1 = 32'd965
; 
32'd131976: dataIn1 = 32'd966
; 
32'd131977: dataIn1 = 32'd1838
; 
32'd131978: dataIn1 = 32'd1840
; 
32'd131979: dataIn1 = 32'd2033
; 
32'd131980: dataIn1 = 32'd966
; 
32'd131981: dataIn1 = 32'd968
; 
32'd131982: dataIn1 = 32'd1036
; 
32'd131983: dataIn1 = 32'd1837
; 
32'd131984: dataIn1 = 32'd1841
; 
32'd131985: dataIn1 = 32'd2034
; 
32'd131986: dataIn1 = 32'd199
; 
32'd131987: dataIn1 = 32'd967
; 
32'd131988: dataIn1 = 32'd968
; 
32'd131989: dataIn1 = 32'd1842
; 
32'd131990: dataIn1 = 32'd1844
; 
32'd131991: dataIn1 = 32'd2035
; 
32'd131992: dataIn1 = 32'd967
; 
32'd131993: dataIn1 = 32'd971
; 
32'd131994: dataIn1 = 32'd1037
; 
32'd131995: dataIn1 = 32'd1843
; 
32'd131996: dataIn1 = 32'd1852
; 
32'd131997: dataIn1 = 32'd2036
; 
32'd131998: dataIn1 = 32'd970
; 
32'd131999: dataIn1 = 32'd972
; 
32'd132000: dataIn1 = 32'd1038
; 
32'd132001: dataIn1 = 32'd1846
; 
32'd132002: dataIn1 = 32'd1850
; 
32'd132003: dataIn1 = 32'd2037
; 
32'd132004: dataIn1 = 32'd202
; 
32'd132005: dataIn1 = 32'd969
; 
32'd132006: dataIn1 = 32'd970
; 
32'd132007: dataIn1 = 32'd1845
; 
32'd132008: dataIn1 = 32'd1848
; 
32'd132009: dataIn1 = 32'd2038
; 
32'd132010: dataIn1 = 32'd969
; 
32'd132011: dataIn1 = 32'd2039
; 
32'd132012: dataIn1 = 32'd2534
; 
32'd132013: dataIn1 = 32'd3405
; 
32'd132014: dataIn1 = 32'd3406
; 
32'd132015: dataIn1 = 32'd3408
; 
32'd132016: dataIn1 = 32'd5306
; 
32'd132017: dataIn1 = 32'd125
; 
32'd132018: dataIn1 = 32'd971
; 
32'd132019: dataIn1 = 32'd972
; 
32'd132020: dataIn1 = 32'd1849
; 
32'd132021: dataIn1 = 32'd1851
; 
32'd132022: dataIn1 = 32'd2040
; 
32'd132023: dataIn1 = 32'd390
; 
32'd132024: dataIn1 = 32'd393
; 
32'd132025: dataIn1 = 32'd745
; 
32'd132026: dataIn1 = 32'd750
; 
32'd132027: dataIn1 = 32'd1856
; 
32'd132028: dataIn1 = 32'd2041
; 
32'd132029: dataIn1 = 32'd2042
; 
32'd132030: dataIn1 = 32'd3415
; 
32'd132031: dataIn1 = 32'd3470
; 
32'd132032: dataIn1 = 32'd266
; 
32'd132033: dataIn1 = 32'd393
; 
32'd132034: dataIn1 = 32'd750
; 
32'd132035: dataIn1 = 32'd959
; 
32'd132036: dataIn1 = 32'd1859
; 
32'd132037: dataIn1 = 32'd2041
; 
32'd132038: dataIn1 = 32'd2042
; 
32'd132039: dataIn1 = 32'd973
; 
32'd132040: dataIn1 = 32'd975
; 
32'd132041: dataIn1 = 32'd1861
; 
32'd132042: dataIn1 = 32'd1863
; 
32'd132043: dataIn1 = 32'd2043
; 
32'd132044: dataIn1 = 32'd2526
; 
32'd132045: dataIn1 = 32'd2528
; 
32'd132046: dataIn1 = 32'd975
; 
32'd132047: dataIn1 = 32'd978
; 
32'd132048: dataIn1 = 32'd1860
; 
32'd132049: dataIn1 = 32'd1864
; 
32'd132050: dataIn1 = 32'd2044
; 
32'd132051: dataIn1 = 32'd2536
; 
32'd132052: dataIn1 = 32'd2537
; 
32'd132053: dataIn1 = 32'd401
; 
32'd132054: dataIn1 = 32'd767
; 
32'd132055: dataIn1 = 32'd973
; 
32'd132056: dataIn1 = 32'd1862
; 
32'd132057: dataIn1 = 32'd2045
; 
32'd132058: dataIn1 = 32'd2523
; 
32'd132059: dataIn1 = 32'd2524
; 
32'd132060: dataIn1 = 32'd977
; 
32'd132061: dataIn1 = 32'd978
; 
32'd132062: dataIn1 = 32'd1865
; 
32'd132063: dataIn1 = 32'd1867
; 
32'd132064: dataIn1 = 32'd2046
; 
32'd132065: dataIn1 = 32'd2529
; 
32'd132066: dataIn1 = 32'd2530
; 
32'd132067: dataIn1 = 32'd977
; 
32'd132068: dataIn1 = 32'd982
; 
32'd132069: dataIn1 = 32'd1866
; 
32'd132070: dataIn1 = 32'd1876
; 
32'd132071: dataIn1 = 32'd2047
; 
32'd132072: dataIn1 = 32'd2540
; 
32'd132073: dataIn1 = 32'd2541
; 
32'd132074: dataIn1 = 32'd4615
; 
32'd132075: dataIn1 = 32'd2048
; 
32'd132076: dataIn1 = 32'd3417
; 
32'd132077: dataIn1 = 32'd3418
; 
32'd132078: dataIn1 = 32'd4624
; 
32'd132079: dataIn1 = 32'd4625
; 
32'd132080: dataIn1 = 32'd4629
; 
32'd132081: dataIn1 = 32'd10261
; 
32'd132082: dataIn1 = 32'd979
; 
32'd132083: dataIn1 = 32'd980
; 
32'd132084: dataIn1 = 32'd1868
; 
32'd132085: dataIn1 = 32'd1871
; 
32'd132086: dataIn1 = 32'd2049
; 
32'd132087: dataIn1 = 32'd3039
; 
32'd132088: dataIn1 = 32'd5428
; 
32'd132089: dataIn1 = 32'd5511
; 
32'd132090: dataIn1 = 32'd979
; 
32'd132091: dataIn1 = 32'd984
; 
32'd132092: dataIn1 = 32'd1043
; 
32'd132093: dataIn1 = 32'd1870
; 
32'd132094: dataIn1 = 32'd1879
; 
32'd132095: dataIn1 = 32'd2050
; 
32'd132096: dataIn1 = 32'd982
; 
32'd132097: dataIn1 = 32'd983
; 
32'd132098: dataIn1 = 32'd1873
; 
32'd132099: dataIn1 = 32'd1875
; 
32'd132100: dataIn1 = 32'd2051
; 
32'd132101: dataIn1 = 32'd2531
; 
32'd132102: dataIn1 = 32'd2532
; 
32'd132103: dataIn1 = 32'd4606
; 
32'd132104: dataIn1 = 32'd4634
; 
32'd132105: dataIn1 = 32'd132
; 
32'd132106: dataIn1 = 32'd984
; 
32'd132107: dataIn1 = 32'd985
; 
32'd132108: dataIn1 = 32'd1878
; 
32'd132109: dataIn1 = 32'd1880
; 
32'd132110: dataIn1 = 32'd2052
; 
32'd132111: dataIn1 = 32'd985
; 
32'd132112: dataIn1 = 32'd987
; 
32'd132113: dataIn1 = 32'd1044
; 
32'd132114: dataIn1 = 32'd1877
; 
32'd132115: dataIn1 = 32'd1881
; 
32'd132116: dataIn1 = 32'd2053
; 
32'd132117: dataIn1 = 32'd215
; 
32'd132118: dataIn1 = 32'd986
; 
32'd132119: dataIn1 = 32'd987
; 
32'd132120: dataIn1 = 32'd1882
; 
32'd132121: dataIn1 = 32'd1884
; 
32'd132122: dataIn1 = 32'd2054
; 
32'd132123: dataIn1 = 32'd986
; 
32'd132124: dataIn1 = 32'd990
; 
32'd132125: dataIn1 = 32'd1045
; 
32'd132126: dataIn1 = 32'd1883
; 
32'd132127: dataIn1 = 32'd1892
; 
32'd132128: dataIn1 = 32'd2055
; 
32'd132129: dataIn1 = 32'd989
; 
32'd132130: dataIn1 = 32'd991
; 
32'd132131: dataIn1 = 32'd1046
; 
32'd132132: dataIn1 = 32'd1886
; 
32'd132133: dataIn1 = 32'd1890
; 
32'd132134: dataIn1 = 32'd2056
; 
32'd132135: dataIn1 = 32'd218
; 
32'd132136: dataIn1 = 32'd988
; 
32'd132137: dataIn1 = 32'd989
; 
32'd132138: dataIn1 = 32'd1885
; 
32'd132139: dataIn1 = 32'd1888
; 
32'd132140: dataIn1 = 32'd2057
; 
32'd132141: dataIn1 = 32'd988
; 
32'd132142: dataIn1 = 32'd992
; 
32'd132143: dataIn1 = 32'd1047
; 
32'd132144: dataIn1 = 32'd1887
; 
32'd132145: dataIn1 = 32'd1895
; 
32'd132146: dataIn1 = 32'd2058
; 
32'd132147: dataIn1 = 32'd134
; 
32'd132148: dataIn1 = 32'd990
; 
32'd132149: dataIn1 = 32'd991
; 
32'd132150: dataIn1 = 32'd1889
; 
32'd132151: dataIn1 = 32'd1891
; 
32'd132152: dataIn1 = 32'd2059
; 
32'd132153: dataIn1 = 32'd135
; 
32'd132154: dataIn1 = 32'd992
; 
32'd132155: dataIn1 = 32'd993
; 
32'd132156: dataIn1 = 32'd1894
; 
32'd132157: dataIn1 = 32'd1896
; 
32'd132158: dataIn1 = 32'd2060
; 
32'd132159: dataIn1 = 32'd993
; 
32'd132160: dataIn1 = 32'd995
; 
32'd132161: dataIn1 = 32'd1048
; 
32'd132162: dataIn1 = 32'd1893
; 
32'd132163: dataIn1 = 32'd1897
; 
32'd132164: dataIn1 = 32'd2061
; 
32'd132165: dataIn1 = 32'd221
; 
32'd132166: dataIn1 = 32'd994
; 
32'd132167: dataIn1 = 32'd995
; 
32'd132168: dataIn1 = 32'd1898
; 
32'd132169: dataIn1 = 32'd1900
; 
32'd132170: dataIn1 = 32'd2062
; 
32'd132171: dataIn1 = 32'd994
; 
32'd132172: dataIn1 = 32'd998
; 
32'd132173: dataIn1 = 32'd1049
; 
32'd132174: dataIn1 = 32'd1899
; 
32'd132175: dataIn1 = 32'd1908
; 
32'd132176: dataIn1 = 32'd2063
; 
32'd132177: dataIn1 = 32'd997
; 
32'd132178: dataIn1 = 32'd999
; 
32'd132179: dataIn1 = 32'd1050
; 
32'd132180: dataIn1 = 32'd1902
; 
32'd132181: dataIn1 = 32'd1906
; 
32'd132182: dataIn1 = 32'd2064
; 
32'd132183: dataIn1 = 32'd224
; 
32'd132184: dataIn1 = 32'd996
; 
32'd132185: dataIn1 = 32'd997
; 
32'd132186: dataIn1 = 32'd1901
; 
32'd132187: dataIn1 = 32'd1904
; 
32'd132188: dataIn1 = 32'd2065
; 
32'd132189: dataIn1 = 32'd996
; 
32'd132190: dataIn1 = 32'd1000
; 
32'd132191: dataIn1 = 32'd1051
; 
32'd132192: dataIn1 = 32'd1903
; 
32'd132193: dataIn1 = 32'd1911
; 
32'd132194: dataIn1 = 32'd2066
; 
32'd132195: dataIn1 = 32'd137
; 
32'd132196: dataIn1 = 32'd998
; 
32'd132197: dataIn1 = 32'd999
; 
32'd132198: dataIn1 = 32'd1905
; 
32'd132199: dataIn1 = 32'd1907
; 
32'd132200: dataIn1 = 32'd2067
; 
32'd132201: dataIn1 = 32'd138
; 
32'd132202: dataIn1 = 32'd1000
; 
32'd132203: dataIn1 = 32'd1001
; 
32'd132204: dataIn1 = 32'd1910
; 
32'd132205: dataIn1 = 32'd1912
; 
32'd132206: dataIn1 = 32'd2068
; 
32'd132207: dataIn1 = 32'd1001
; 
32'd132208: dataIn1 = 32'd1003
; 
32'd132209: dataIn1 = 32'd1052
; 
32'd132210: dataIn1 = 32'd1909
; 
32'd132211: dataIn1 = 32'd1913
; 
32'd132212: dataIn1 = 32'd2069
; 
32'd132213: dataIn1 = 32'd227
; 
32'd132214: dataIn1 = 32'd1002
; 
32'd132215: dataIn1 = 32'd1003
; 
32'd132216: dataIn1 = 32'd1914
; 
32'd132217: dataIn1 = 32'd1916
; 
32'd132218: dataIn1 = 32'd2070
; 
32'd132219: dataIn1 = 32'd1002
; 
32'd132220: dataIn1 = 32'd1006
; 
32'd132221: dataIn1 = 32'd1053
; 
32'd132222: dataIn1 = 32'd1915
; 
32'd132223: dataIn1 = 32'd1924
; 
32'd132224: dataIn1 = 32'd2071
; 
32'd132225: dataIn1 = 32'd1005
; 
32'd132226: dataIn1 = 32'd1007
; 
32'd132227: dataIn1 = 32'd1054
; 
32'd132228: dataIn1 = 32'd1918
; 
32'd132229: dataIn1 = 32'd1922
; 
32'd132230: dataIn1 = 32'd2072
; 
32'd132231: dataIn1 = 32'd230
; 
32'd132232: dataIn1 = 32'd1004
; 
32'd132233: dataIn1 = 32'd1005
; 
32'd132234: dataIn1 = 32'd1917
; 
32'd132235: dataIn1 = 32'd1920
; 
32'd132236: dataIn1 = 32'd2073
; 
32'd132237: dataIn1 = 32'd1004
; 
32'd132238: dataIn1 = 32'd1008
; 
32'd132239: dataIn1 = 32'd1055
; 
32'd132240: dataIn1 = 32'd1919
; 
32'd132241: dataIn1 = 32'd1927
; 
32'd132242: dataIn1 = 32'd2074
; 
32'd132243: dataIn1 = 32'd140
; 
32'd132244: dataIn1 = 32'd1006
; 
32'd132245: dataIn1 = 32'd1007
; 
32'd132246: dataIn1 = 32'd1921
; 
32'd132247: dataIn1 = 32'd1923
; 
32'd132248: dataIn1 = 32'd2075
; 
32'd132249: dataIn1 = 32'd141
; 
32'd132250: dataIn1 = 32'd1008
; 
32'd132251: dataIn1 = 32'd1009
; 
32'd132252: dataIn1 = 32'd1926
; 
32'd132253: dataIn1 = 32'd1928
; 
32'd132254: dataIn1 = 32'd2076
; 
32'd132255: dataIn1 = 32'd1009
; 
32'd132256: dataIn1 = 32'd1011
; 
32'd132257: dataIn1 = 32'd1056
; 
32'd132258: dataIn1 = 32'd1925
; 
32'd132259: dataIn1 = 32'd1929
; 
32'd132260: dataIn1 = 32'd2077
; 
32'd132261: dataIn1 = 32'd233
; 
32'd132262: dataIn1 = 32'd1010
; 
32'd132263: dataIn1 = 32'd1011
; 
32'd132264: dataIn1 = 32'd1930
; 
32'd132265: dataIn1 = 32'd1932
; 
32'd132266: dataIn1 = 32'd2078
; 
32'd132267: dataIn1 = 32'd1010
; 
32'd132268: dataIn1 = 32'd1014
; 
32'd132269: dataIn1 = 32'd1057
; 
32'd132270: dataIn1 = 32'd1931
; 
32'd132271: dataIn1 = 32'd1940
; 
32'd132272: dataIn1 = 32'd2079
; 
32'd132273: dataIn1 = 32'd1013
; 
32'd132274: dataIn1 = 32'd1015
; 
32'd132275: dataIn1 = 32'd1058
; 
32'd132276: dataIn1 = 32'd1934
; 
32'd132277: dataIn1 = 32'd1938
; 
32'd132278: dataIn1 = 32'd2080
; 
32'd132279: dataIn1 = 32'd236
; 
32'd132280: dataIn1 = 32'd1012
; 
32'd132281: dataIn1 = 32'd1013
; 
32'd132282: dataIn1 = 32'd1933
; 
32'd132283: dataIn1 = 32'd1936
; 
32'd132284: dataIn1 = 32'd2081
; 
32'd132285: dataIn1 = 32'd1012
; 
32'd132286: dataIn1 = 32'd1016
; 
32'd132287: dataIn1 = 32'd1059
; 
32'd132288: dataIn1 = 32'd1935
; 
32'd132289: dataIn1 = 32'd1943
; 
32'd132290: dataIn1 = 32'd2082
; 
32'd132291: dataIn1 = 32'd143
; 
32'd132292: dataIn1 = 32'd1014
; 
32'd132293: dataIn1 = 32'd1015
; 
32'd132294: dataIn1 = 32'd1937
; 
32'd132295: dataIn1 = 32'd1939
; 
32'd132296: dataIn1 = 32'd2083
; 
32'd132297: dataIn1 = 32'd144
; 
32'd132298: dataIn1 = 32'd1016
; 
32'd132299: dataIn1 = 32'd1017
; 
32'd132300: dataIn1 = 32'd1942
; 
32'd132301: dataIn1 = 32'd1944
; 
32'd132302: dataIn1 = 32'd2084
; 
32'd132303: dataIn1 = 32'd1017
; 
32'd132304: dataIn1 = 32'd1019
; 
32'd132305: dataIn1 = 32'd1060
; 
32'd132306: dataIn1 = 32'd1941
; 
32'd132307: dataIn1 = 32'd1945
; 
32'd132308: dataIn1 = 32'd2085
; 
32'd132309: dataIn1 = 32'd239
; 
32'd132310: dataIn1 = 32'd1018
; 
32'd132311: dataIn1 = 32'd1019
; 
32'd132312: dataIn1 = 32'd1946
; 
32'd132313: dataIn1 = 32'd1948
; 
32'd132314: dataIn1 = 32'd2086
; 
32'd132315: dataIn1 = 32'd1018
; 
32'd132316: dataIn1 = 32'd1022
; 
32'd132317: dataIn1 = 32'd1061
; 
32'd132318: dataIn1 = 32'd1947
; 
32'd132319: dataIn1 = 32'd1956
; 
32'd132320: dataIn1 = 32'd2087
; 
32'd132321: dataIn1 = 32'd1021
; 
32'd132322: dataIn1 = 32'd1023
; 
32'd132323: dataIn1 = 32'd1062
; 
32'd132324: dataIn1 = 32'd1950
; 
32'd132325: dataIn1 = 32'd1954
; 
32'd132326: dataIn1 = 32'd2088
; 
32'd132327: dataIn1 = 32'd242
; 
32'd132328: dataIn1 = 32'd1020
; 
32'd132329: dataIn1 = 32'd1021
; 
32'd132330: dataIn1 = 32'd1949
; 
32'd132331: dataIn1 = 32'd1952
; 
32'd132332: dataIn1 = 32'd2089
; 
32'd132333: dataIn1 = 32'd1020
; 
32'd132334: dataIn1 = 32'd1024
; 
32'd132335: dataIn1 = 32'd1063
; 
32'd132336: dataIn1 = 32'd1951
; 
32'd132337: dataIn1 = 32'd1959
; 
32'd132338: dataIn1 = 32'd2090
; 
32'd132339: dataIn1 = 32'd146
; 
32'd132340: dataIn1 = 32'd1022
; 
32'd132341: dataIn1 = 32'd1023
; 
32'd132342: dataIn1 = 32'd1953
; 
32'd132343: dataIn1 = 32'd1955
; 
32'd132344: dataIn1 = 32'd2091
; 
32'd132345: dataIn1 = 32'd147
; 
32'd132346: dataIn1 = 32'd1024
; 
32'd132347: dataIn1 = 32'd1025
; 
32'd132348: dataIn1 = 32'd1958
; 
32'd132349: dataIn1 = 32'd1960
; 
32'd132350: dataIn1 = 32'd2092
; 
32'd132351: dataIn1 = 32'd1025
; 
32'd132352: dataIn1 = 32'd1027
; 
32'd132353: dataIn1 = 32'd1064
; 
32'd132354: dataIn1 = 32'd1957
; 
32'd132355: dataIn1 = 32'd1961
; 
32'd132356: dataIn1 = 32'd2093
; 
32'd132357: dataIn1 = 32'd245
; 
32'd132358: dataIn1 = 32'd1026
; 
32'd132359: dataIn1 = 32'd1027
; 
32'd132360: dataIn1 = 32'd1962
; 
32'd132361: dataIn1 = 32'd1964
; 
32'd132362: dataIn1 = 32'd2094
; 
32'd132363: dataIn1 = 32'd1026
; 
32'd132364: dataIn1 = 32'd1030
; 
32'd132365: dataIn1 = 32'd1065
; 
32'd132366: dataIn1 = 32'd1963
; 
32'd132367: dataIn1 = 32'd1972
; 
32'd132368: dataIn1 = 32'd2095
; 
32'd132369: dataIn1 = 32'd149
; 
32'd132370: dataIn1 = 32'd1029
; 
32'd132371: dataIn1 = 32'd1031
; 
32'd132372: dataIn1 = 32'd1066
; 
32'd132373: dataIn1 = 32'd1966
; 
32'd132374: dataIn1 = 32'd1970
; 
32'd132375: dataIn1 = 32'd2096
; 
32'd132376: dataIn1 = 32'd248
; 
32'd132377: dataIn1 = 32'd1028
; 
32'd132378: dataIn1 = 32'd1029
; 
32'd132379: dataIn1 = 32'd1066
; 
32'd132380: dataIn1 = 32'd1965
; 
32'd132381: dataIn1 = 32'd1968
; 
32'd132382: dataIn1 = 32'd2097
; 
32'd132383: dataIn1 = 32'd248
; 
32'd132384: dataIn1 = 32'd1028
; 
32'd132385: dataIn1 = 32'd1032
; 
32'd132386: dataIn1 = 32'd1067
; 
32'd132387: dataIn1 = 32'd1967
; 
32'd132388: dataIn1 = 32'd1975
; 
32'd132389: dataIn1 = 32'd2098
; 
32'd132390: dataIn1 = 32'd149
; 
32'd132391: dataIn1 = 32'd1030
; 
32'd132392: dataIn1 = 32'd1031
; 
32'd132393: dataIn1 = 32'd1969
; 
32'd132394: dataIn1 = 32'd1971
; 
32'd132395: dataIn1 = 32'd2099
; 
32'd132396: dataIn1 = 32'd150
; 
32'd132397: dataIn1 = 32'd1032
; 
32'd132398: dataIn1 = 32'd1033
; 
32'd132399: dataIn1 = 32'd1067
; 
32'd132400: dataIn1 = 32'd1974
; 
32'd132401: dataIn1 = 32'd1976
; 
32'd132402: dataIn1 = 32'd2100
; 
32'd132403: dataIn1 = 32'd557
; 
32'd132404: dataIn1 = 32'd2101
; 
32'd132405: dataIn1 = 32'd10247
; 
32'd132406: dataIn1 = 32'd10248
; 
32'd132407: dataIn1 = 32'd11654
; 
32'd132408: dataIn1 = 32'd11655
; 
32'd132409: dataIn1 = 32'd11656
; 
32'd132410: dataIn1 = 32'd2102
; 
32'd132411: dataIn1 = 32'd3457
; 
32'd132412: dataIn1 = 32'd6693
; 
32'd132413: dataIn1 = 32'd6730
; 
32'd132414: dataIn1 = 32'd9311
; 
32'd132415: dataIn1 = 32'd9312
; 
32'd132416: dataIn1 = 32'd9314
; 
32'd132417: dataIn1 = 32'd2103
; 
32'd132418: dataIn1 = 32'd6826
; 
32'd132419: dataIn1 = 32'd6827
; 
32'd132420: dataIn1 = 32'd10286
; 
32'd132421: dataIn1 = 32'd2104
; 
32'd132422: dataIn1 = 32'd2120
; 
32'd132423: dataIn1 = 32'd6694
; 
32'd132424: dataIn1 = 32'd6731
; 
32'd132425: dataIn1 = 32'd9315
; 
32'd132426: dataIn1 = 32'd9317
; 
32'd132427: dataIn1 = 32'd9318
; 
32'd132428: dataIn1 = 32'd2105
; 
32'd132429: dataIn1 = 32'd5647
; 
32'd132430: dataIn1 = 32'd6843
; 
32'd132431: dataIn1 = 32'd9266
; 
32'd132432: dataIn1 = 32'd10290
; 
32'd132433: dataIn1 = 32'd10291
; 
32'd132434: dataIn1 = 32'd28
; 
32'd132435: dataIn1 = 32'd29
; 
32'd132436: dataIn1 = 32'd2106
; 
32'd132437: dataIn1 = 32'd2107
; 
32'd132438: dataIn1 = 32'd2108
; 
32'd132439: dataIn1 = 32'd2140
; 
32'd132440: dataIn1 = 32'd2141
; 
32'd132441: dataIn1 = 32'd18
; 
32'd132442: dataIn1 = 32'd29
; 
32'd132443: dataIn1 = 32'd1139
; 
32'd132444: dataIn1 = 32'd2106
; 
32'd132445: dataIn1 = 32'd2107
; 
32'd132446: dataIn1 = 32'd2108
; 
32'd132447: dataIn1 = 32'd2109
; 
32'd132448: dataIn1 = 32'd5516
; 
32'd132449: dataIn1 = 32'd18
; 
32'd132450: dataIn1 = 32'd28
; 
32'd132451: dataIn1 = 32'd1138
; 
32'd132452: dataIn1 = 32'd2106
; 
32'd132453: dataIn1 = 32'd2107
; 
32'd132454: dataIn1 = 32'd2108
; 
32'd132455: dataIn1 = 32'd2748
; 
32'd132456: dataIn1 = 32'd5517
; 
32'd132457: dataIn1 = 32'd19
; 
32'd132458: dataIn1 = 32'd29
; 
32'd132459: dataIn1 = 32'd1139
; 
32'd132460: dataIn1 = 32'd2107
; 
32'd132461: dataIn1 = 32'd2109
; 
32'd132462: dataIn1 = 32'd2110
; 
32'd132463: dataIn1 = 32'd2111
; 
32'd132464: dataIn1 = 32'd5519
; 
32'd132465: dataIn1 = 32'd29
; 
32'd132466: dataIn1 = 32'd30
; 
32'd132467: dataIn1 = 32'd2109
; 
32'd132468: dataIn1 = 32'd2110
; 
32'd132469: dataIn1 = 32'd2111
; 
32'd132470: dataIn1 = 32'd2143
; 
32'd132471: dataIn1 = 32'd2144
; 
32'd132472: dataIn1 = 32'd19
; 
32'd132473: dataIn1 = 32'd30
; 
32'd132474: dataIn1 = 32'd1140
; 
32'd132475: dataIn1 = 32'd2109
; 
32'd132476: dataIn1 = 32'd2110
; 
32'd132477: dataIn1 = 32'd2111
; 
32'd132478: dataIn1 = 32'd2112
; 
32'd132479: dataIn1 = 32'd5518
; 
32'd132480: dataIn1 = 32'd9676
; 
32'd132481: dataIn1 = 32'd30
; 
32'd132482: dataIn1 = 32'd2111
; 
32'd132483: dataIn1 = 32'd2112
; 
32'd132484: dataIn1 = 32'd9449
; 
32'd132485: dataIn1 = 32'd9450
; 
32'd132486: dataIn1 = 32'd9452
; 
32'd132487: dataIn1 = 32'd9676
; 
32'd132488: dataIn1 = 32'd30
; 
32'd132489: dataIn1 = 32'd2113
; 
32'd132490: dataIn1 = 32'd9450
; 
32'd132491: dataIn1 = 32'd9819
; 
32'd132492: dataIn1 = 32'd9820
; 
32'd132493: dataIn1 = 32'd9832
; 
32'd132494: dataIn1 = 32'd10155
; 
32'd132495: dataIn1 = 32'd2114
; 
32'd132496: dataIn1 = 32'd9811
; 
32'd132497: dataIn1 = 32'd9813
; 
32'd132498: dataIn1 = 32'd9814
; 
32'd132499: dataIn1 = 32'd9821
; 
32'd132500: dataIn1 = 32'd9826
; 
32'd132501: dataIn1 = 32'd10152
; 
32'd132502: dataIn1 = 32'd2115
; 
32'd132503: dataIn1 = 32'd2116
; 
32'd132504: dataIn1 = 32'd2117
; 
32'd132505: dataIn1 = 32'd10152
; 
32'd132506: dataIn1 = 32'd10153
; 
32'd132507: dataIn1 = 32'd10154
; 
32'd132508: dataIn1 = 32'd10225
; 
32'd132509: dataIn1 = 32'd31
; 
32'd132510: dataIn1 = 32'd32
; 
32'd132511: dataIn1 = 32'd2115
; 
32'd132512: dataIn1 = 32'd2116
; 
32'd132513: dataIn1 = 32'd2117
; 
32'd132514: dataIn1 = 32'd2149
; 
32'd132515: dataIn1 = 32'd2150
; 
32'd132516: dataIn1 = 32'd9462
; 
32'd132517: dataIn1 = 32'd10153
; 
32'd132518: dataIn1 = 32'd21
; 
32'd132519: dataIn1 = 32'd32
; 
32'd132520: dataIn1 = 32'd1142
; 
32'd132521: dataIn1 = 32'd2115
; 
32'd132522: dataIn1 = 32'd2116
; 
32'd132523: dataIn1 = 32'd2117
; 
32'd132524: dataIn1 = 32'd2118
; 
32'd132525: dataIn1 = 32'd5522
; 
32'd132526: dataIn1 = 32'd10225
; 
32'd132527: dataIn1 = 32'd22
; 
32'd132528: dataIn1 = 32'd32
; 
32'd132529: dataIn1 = 32'd1142
; 
32'd132530: dataIn1 = 32'd2117
; 
32'd132531: dataIn1 = 32'd2118
; 
32'd132532: dataIn1 = 32'd2119
; 
32'd132533: dataIn1 = 32'd2120
; 
32'd132534: dataIn1 = 32'd5524
; 
32'd132535: dataIn1 = 32'd32
; 
32'd132536: dataIn1 = 32'd33
; 
32'd132537: dataIn1 = 32'd2118
; 
32'd132538: dataIn1 = 32'd2119
; 
32'd132539: dataIn1 = 32'd2120
; 
32'd132540: dataIn1 = 32'd2152
; 
32'd132541: dataIn1 = 32'd2153
; 
32'd132542: dataIn1 = 32'd22
; 
32'd132543: dataIn1 = 32'd33
; 
32'd132544: dataIn1 = 32'd2104
; 
32'd132545: dataIn1 = 32'd2118
; 
32'd132546: dataIn1 = 32'd2119
; 
32'd132547: dataIn1 = 32'd2120
; 
32'd132548: dataIn1 = 32'd2121
; 
32'd132549: dataIn1 = 32'd6731
; 
32'd132550: dataIn1 = 32'd9317
; 
32'd132551: dataIn1 = 32'd23
; 
32'd132552: dataIn1 = 32'd33
; 
32'd132553: dataIn1 = 32'd2120
; 
32'd132554: dataIn1 = 32'd2121
; 
32'd132555: dataIn1 = 32'd9317
; 
32'd132556: dataIn1 = 32'd34
; 
32'd132557: dataIn1 = 32'd35
; 
32'd132558: dataIn1 = 32'd2122
; 
32'd132559: dataIn1 = 32'd2123
; 
32'd132560: dataIn1 = 32'd2124
; 
32'd132561: dataIn1 = 32'd2156
; 
32'd132562: dataIn1 = 32'd2157
; 
32'd132563: dataIn1 = 32'd24
; 
32'd132564: dataIn1 = 32'd35
; 
32'd132565: dataIn1 = 32'd2122
; 
32'd132566: dataIn1 = 32'd2123
; 
32'd132567: dataIn1 = 32'd2124
; 
32'd132568: dataIn1 = 32'd2125
; 
32'd132569: dataIn1 = 32'd2126
; 
32'd132570: dataIn1 = 32'd24
; 
32'd132571: dataIn1 = 32'd34
; 
32'd132572: dataIn1 = 32'd2122
; 
32'd132573: dataIn1 = 32'd2123
; 
32'd132574: dataIn1 = 32'd2124
; 
32'd132575: dataIn1 = 32'd25
; 
32'd132576: dataIn1 = 32'd35
; 
32'd132577: dataIn1 = 32'd2123
; 
32'd132578: dataIn1 = 32'd2125
; 
32'd132579: dataIn1 = 32'd2126
; 
32'd132580: dataIn1 = 32'd2127
; 
32'd132581: dataIn1 = 32'd2128
; 
32'd132582: dataIn1 = 32'd24
; 
32'd132583: dataIn1 = 32'd25
; 
32'd132584: dataIn1 = 32'd2123
; 
32'd132585: dataIn1 = 32'd2125
; 
32'd132586: dataIn1 = 32'd2126
; 
32'd132587: dataIn1 = 32'd3434
; 
32'd132588: dataIn1 = 32'd3457
; 
32'd132589: dataIn1 = 32'd35
; 
32'd132590: dataIn1 = 32'd36
; 
32'd132591: dataIn1 = 32'd2125
; 
32'd132592: dataIn1 = 32'd2127
; 
32'd132593: dataIn1 = 32'd2128
; 
32'd132594: dataIn1 = 32'd2159
; 
32'd132595: dataIn1 = 32'd2160
; 
32'd132596: dataIn1 = 32'd25
; 
32'd132597: dataIn1 = 32'd36
; 
32'd132598: dataIn1 = 32'd2125
; 
32'd132599: dataIn1 = 32'd2127
; 
32'd132600: dataIn1 = 32'd2128
; 
32'd132601: dataIn1 = 32'd2129
; 
32'd132602: dataIn1 = 32'd2130
; 
32'd132603: dataIn1 = 32'd26
; 
32'd132604: dataIn1 = 32'd36
; 
32'd132605: dataIn1 = 32'd2128
; 
32'd132606: dataIn1 = 32'd2129
; 
32'd132607: dataIn1 = 32'd2130
; 
32'd132608: dataIn1 = 32'd2131
; 
32'd132609: dataIn1 = 32'd2132
; 
32'd132610: dataIn1 = 32'd25
; 
32'd132611: dataIn1 = 32'd26
; 
32'd132612: dataIn1 = 32'd2128
; 
32'd132613: dataIn1 = 32'd2129
; 
32'd132614: dataIn1 = 32'd2130
; 
32'd132615: dataIn1 = 32'd3433
; 
32'd132616: dataIn1 = 32'd3436
; 
32'd132617: dataIn1 = 32'd36
; 
32'd132618: dataIn1 = 32'd37
; 
32'd132619: dataIn1 = 32'd2129
; 
32'd132620: dataIn1 = 32'd2131
; 
32'd132621: dataIn1 = 32'd2132
; 
32'd132622: dataIn1 = 32'd2162
; 
32'd132623: dataIn1 = 32'd2163
; 
32'd132624: dataIn1 = 32'd26
; 
32'd132625: dataIn1 = 32'd37
; 
32'd132626: dataIn1 = 32'd2129
; 
32'd132627: dataIn1 = 32'd2131
; 
32'd132628: dataIn1 = 32'd2132
; 
32'd132629: dataIn1 = 32'd2133
; 
32'd132630: dataIn1 = 32'd2134
; 
32'd132631: dataIn1 = 32'd27
; 
32'd132632: dataIn1 = 32'd37
; 
32'd132633: dataIn1 = 32'd2132
; 
32'd132634: dataIn1 = 32'd2133
; 
32'd132635: dataIn1 = 32'd2134
; 
32'd132636: dataIn1 = 32'd2135
; 
32'd132637: dataIn1 = 32'd2136
; 
32'd132638: dataIn1 = 32'd26
; 
32'd132639: dataIn1 = 32'd27
; 
32'd132640: dataIn1 = 32'd2132
; 
32'd132641: dataIn1 = 32'd2133
; 
32'd132642: dataIn1 = 32'd2134
; 
32'd132643: dataIn1 = 32'd3435
; 
32'd132644: dataIn1 = 32'd3437
; 
32'd132645: dataIn1 = 32'd37
; 
32'd132646: dataIn1 = 32'd38
; 
32'd132647: dataIn1 = 32'd2133
; 
32'd132648: dataIn1 = 32'd2135
; 
32'd132649: dataIn1 = 32'd2136
; 
32'd132650: dataIn1 = 32'd2165
; 
32'd132651: dataIn1 = 32'd2166
; 
32'd132652: dataIn1 = 32'd27
; 
32'd132653: dataIn1 = 32'd38
; 
32'd132654: dataIn1 = 32'd2133
; 
32'd132655: dataIn1 = 32'd2135
; 
32'd132656: dataIn1 = 32'd2136
; 
32'd132657: dataIn1 = 32'd2137
; 
32'd132658: dataIn1 = 32'd2138
; 
32'd132659: dataIn1 = 32'd28
; 
32'd132660: dataIn1 = 32'd38
; 
32'd132661: dataIn1 = 32'd2136
; 
32'd132662: dataIn1 = 32'd2137
; 
32'd132663: dataIn1 = 32'd2138
; 
32'd132664: dataIn1 = 32'd2139
; 
32'd132665: dataIn1 = 32'd2140
; 
32'd132666: dataIn1 = 32'd27
; 
32'd132667: dataIn1 = 32'd28
; 
32'd132668: dataIn1 = 32'd2136
; 
32'd132669: dataIn1 = 32'd2137
; 
32'd132670: dataIn1 = 32'd2138
; 
32'd132671: dataIn1 = 32'd2748
; 
32'd132672: dataIn1 = 32'd3419
; 
32'd132673: dataIn1 = 32'd38
; 
32'd132674: dataIn1 = 32'd39
; 
32'd132675: dataIn1 = 32'd2137
; 
32'd132676: dataIn1 = 32'd2139
; 
32'd132677: dataIn1 = 32'd2140
; 
32'd132678: dataIn1 = 32'd2168
; 
32'd132679: dataIn1 = 32'd2169
; 
32'd132680: dataIn1 = 32'd28
; 
32'd132681: dataIn1 = 32'd39
; 
32'd132682: dataIn1 = 32'd2106
; 
32'd132683: dataIn1 = 32'd2137
; 
32'd132684: dataIn1 = 32'd2139
; 
32'd132685: dataIn1 = 32'd2140
; 
32'd132686: dataIn1 = 32'd2141
; 
32'd132687: dataIn1 = 32'd29
; 
32'd132688: dataIn1 = 32'd39
; 
32'd132689: dataIn1 = 32'd2106
; 
32'd132690: dataIn1 = 32'd2140
; 
32'd132691: dataIn1 = 32'd2141
; 
32'd132692: dataIn1 = 32'd2142
; 
32'd132693: dataIn1 = 32'd2143
; 
32'd132694: dataIn1 = 32'd39
; 
32'd132695: dataIn1 = 32'd40
; 
32'd132696: dataIn1 = 32'd2141
; 
32'd132697: dataIn1 = 32'd2142
; 
32'd132698: dataIn1 = 32'd2143
; 
32'd132699: dataIn1 = 32'd2171
; 
32'd132700: dataIn1 = 32'd2172
; 
32'd132701: dataIn1 = 32'd29
; 
32'd132702: dataIn1 = 32'd40
; 
32'd132703: dataIn1 = 32'd2110
; 
32'd132704: dataIn1 = 32'd2141
; 
32'd132705: dataIn1 = 32'd2142
; 
32'd132706: dataIn1 = 32'd2143
; 
32'd132707: dataIn1 = 32'd2144
; 
32'd132708: dataIn1 = 32'd30
; 
32'd132709: dataIn1 = 32'd40
; 
32'd132710: dataIn1 = 32'd2110
; 
32'd132711: dataIn1 = 32'd2143
; 
32'd132712: dataIn1 = 32'd2144
; 
32'd132713: dataIn1 = 32'd2145
; 
32'd132714: dataIn1 = 32'd2146
; 
32'd132715: dataIn1 = 32'd40
; 
32'd132716: dataIn1 = 32'd41
; 
32'd132717: dataIn1 = 32'd2144
; 
32'd132718: dataIn1 = 32'd2145
; 
32'd132719: dataIn1 = 32'd2146
; 
32'd132720: dataIn1 = 32'd2174
; 
32'd132721: dataIn1 = 32'd2175
; 
32'd132722: dataIn1 = 32'd9781
; 
32'd132723: dataIn1 = 32'd10157
; 
32'd132724: dataIn1 = 32'd30
; 
32'd132725: dataIn1 = 32'd2144
; 
32'd132726: dataIn1 = 32'd2145
; 
32'd132727: dataIn1 = 32'd2146
; 
32'd132728: dataIn1 = 32'd10155
; 
32'd132729: dataIn1 = 32'd10156
; 
32'd132730: dataIn1 = 32'd10157
; 
32'd132731: dataIn1 = 32'd2147
; 
32'd132732: dataIn1 = 32'd9830
; 
32'd132733: dataIn1 = 32'd9831
; 
32'd132734: dataIn1 = 32'd9833
; 
32'd132735: dataIn1 = 32'd9834
; 
32'd132736: dataIn1 = 32'd9842
; 
32'd132737: dataIn1 = 32'd10156
; 
32'd132738: dataIn1 = 32'd2148
; 
32'd132739: dataIn1 = 32'd9461
; 
32'd132740: dataIn1 = 32'd9466
; 
32'd132741: dataIn1 = 32'd9477
; 
32'd132742: dataIn1 = 32'd9840
; 
32'd132743: dataIn1 = 32'd9841
; 
32'd132744: dataIn1 = 32'd9848
; 
32'd132745: dataIn1 = 32'd2116
; 
32'd132746: dataIn1 = 32'd2149
; 
32'd132747: dataIn1 = 32'd2150
; 
32'd132748: dataIn1 = 32'd9459
; 
32'd132749: dataIn1 = 32'd9461
; 
32'd132750: dataIn1 = 32'd9462
; 
32'd132751: dataIn1 = 32'd9769
; 
32'd132752: dataIn1 = 32'd32
; 
32'd132753: dataIn1 = 32'd42
; 
32'd132754: dataIn1 = 32'd2116
; 
32'd132755: dataIn1 = 32'd2149
; 
32'd132756: dataIn1 = 32'd2150
; 
32'd132757: dataIn1 = 32'd2151
; 
32'd132758: dataIn1 = 32'd2152
; 
32'd132759: dataIn1 = 32'd3603
; 
32'd132760: dataIn1 = 32'd9769
; 
32'd132761: dataIn1 = 32'd2150
; 
32'd132762: dataIn1 = 32'd2151
; 
32'd132763: dataIn1 = 32'd2152
; 
32'd132764: dataIn1 = 32'd3600
; 
32'd132765: dataIn1 = 32'd3602
; 
32'd132766: dataIn1 = 32'd3603
; 
32'd132767: dataIn1 = 32'd3605
; 
32'd132768: dataIn1 = 32'd32
; 
32'd132769: dataIn1 = 32'd43
; 
32'd132770: dataIn1 = 32'd2119
; 
32'd132771: dataIn1 = 32'd2150
; 
32'd132772: dataIn1 = 32'd2151
; 
32'd132773: dataIn1 = 32'd2152
; 
32'd132774: dataIn1 = 32'd2153
; 
32'd132775: dataIn1 = 32'd3605
; 
32'd132776: dataIn1 = 32'd33
; 
32'd132777: dataIn1 = 32'd43
; 
32'd132778: dataIn1 = 32'd2119
; 
32'd132779: dataIn1 = 32'd2152
; 
32'd132780: dataIn1 = 32'd2153
; 
32'd132781: dataIn1 = 32'd2154
; 
32'd132782: dataIn1 = 32'd2155
; 
32'd132783: dataIn1 = 32'd43
; 
32'd132784: dataIn1 = 32'd44
; 
32'd132785: dataIn1 = 32'd2153
; 
32'd132786: dataIn1 = 32'd2154
; 
32'd132787: dataIn1 = 32'd2155
; 
32'd132788: dataIn1 = 32'd2183
; 
32'd132789: dataIn1 = 32'd2184
; 
32'd132790: dataIn1 = 32'd5308
; 
32'd132791: dataIn1 = 32'd33
; 
32'd132792: dataIn1 = 32'd44
; 
32'd132793: dataIn1 = 32'd2153
; 
32'd132794: dataIn1 = 32'd2154
; 
32'd132795: dataIn1 = 32'd2155
; 
32'd132796: dataIn1 = 32'd35
; 
32'd132797: dataIn1 = 32'd45
; 
32'd132798: dataIn1 = 32'd2122
; 
32'd132799: dataIn1 = 32'd2156
; 
32'd132800: dataIn1 = 32'd2157
; 
32'd132801: dataIn1 = 32'd2158
; 
32'd132802: dataIn1 = 32'd2159
; 
32'd132803: dataIn1 = 32'd34
; 
32'd132804: dataIn1 = 32'd45
; 
32'd132805: dataIn1 = 32'd2122
; 
32'd132806: dataIn1 = 32'd2156
; 
32'd132807: dataIn1 = 32'd2157
; 
32'd132808: dataIn1 = 32'd45
; 
32'd132809: dataIn1 = 32'd46
; 
32'd132810: dataIn1 = 32'd2156
; 
32'd132811: dataIn1 = 32'd2158
; 
32'd132812: dataIn1 = 32'd2159
; 
32'd132813: dataIn1 = 32'd2186
; 
32'd132814: dataIn1 = 32'd2188
; 
32'd132815: dataIn1 = 32'd35
; 
32'd132816: dataIn1 = 32'd46
; 
32'd132817: dataIn1 = 32'd2127
; 
32'd132818: dataIn1 = 32'd2156
; 
32'd132819: dataIn1 = 32'd2158
; 
32'd132820: dataIn1 = 32'd2159
; 
32'd132821: dataIn1 = 32'd2160
; 
32'd132822: dataIn1 = 32'd36
; 
32'd132823: dataIn1 = 32'd46
; 
32'd132824: dataIn1 = 32'd2127
; 
32'd132825: dataIn1 = 32'd2159
; 
32'd132826: dataIn1 = 32'd2160
; 
32'd132827: dataIn1 = 32'd2161
; 
32'd132828: dataIn1 = 32'd2162
; 
32'd132829: dataIn1 = 32'd46
; 
32'd132830: dataIn1 = 32'd47
; 
32'd132831: dataIn1 = 32'd2160
; 
32'd132832: dataIn1 = 32'd2161
; 
32'd132833: dataIn1 = 32'd2162
; 
32'd132834: dataIn1 = 32'd2190
; 
32'd132835: dataIn1 = 32'd2191
; 
32'd132836: dataIn1 = 32'd36
; 
32'd132837: dataIn1 = 32'd47
; 
32'd132838: dataIn1 = 32'd2131
; 
32'd132839: dataIn1 = 32'd2160
; 
32'd132840: dataIn1 = 32'd2161
; 
32'd132841: dataIn1 = 32'd2162
; 
32'd132842: dataIn1 = 32'd2163
; 
32'd132843: dataIn1 = 32'd37
; 
32'd132844: dataIn1 = 32'd47
; 
32'd132845: dataIn1 = 32'd2131
; 
32'd132846: dataIn1 = 32'd2162
; 
32'd132847: dataIn1 = 32'd2163
; 
32'd132848: dataIn1 = 32'd2164
; 
32'd132849: dataIn1 = 32'd2165
; 
32'd132850: dataIn1 = 32'd47
; 
32'd132851: dataIn1 = 32'd48
; 
32'd132852: dataIn1 = 32'd2163
; 
32'd132853: dataIn1 = 32'd2164
; 
32'd132854: dataIn1 = 32'd2165
; 
32'd132855: dataIn1 = 32'd2193
; 
32'd132856: dataIn1 = 32'd2194
; 
32'd132857: dataIn1 = 32'd37
; 
32'd132858: dataIn1 = 32'd48
; 
32'd132859: dataIn1 = 32'd2135
; 
32'd132860: dataIn1 = 32'd2163
; 
32'd132861: dataIn1 = 32'd2164
; 
32'd132862: dataIn1 = 32'd2165
; 
32'd132863: dataIn1 = 32'd2166
; 
32'd132864: dataIn1 = 32'd38
; 
32'd132865: dataIn1 = 32'd48
; 
32'd132866: dataIn1 = 32'd2135
; 
32'd132867: dataIn1 = 32'd2165
; 
32'd132868: dataIn1 = 32'd2166
; 
32'd132869: dataIn1 = 32'd2167
; 
32'd132870: dataIn1 = 32'd2168
; 
32'd132871: dataIn1 = 32'd48
; 
32'd132872: dataIn1 = 32'd49
; 
32'd132873: dataIn1 = 32'd2166
; 
32'd132874: dataIn1 = 32'd2167
; 
32'd132875: dataIn1 = 32'd2168
; 
32'd132876: dataIn1 = 32'd2196
; 
32'd132877: dataIn1 = 32'd2197
; 
32'd132878: dataIn1 = 32'd38
; 
32'd132879: dataIn1 = 32'd49
; 
32'd132880: dataIn1 = 32'd2139
; 
32'd132881: dataIn1 = 32'd2166
; 
32'd132882: dataIn1 = 32'd2167
; 
32'd132883: dataIn1 = 32'd2168
; 
32'd132884: dataIn1 = 32'd2169
; 
32'd132885: dataIn1 = 32'd39
; 
32'd132886: dataIn1 = 32'd49
; 
32'd132887: dataIn1 = 32'd2139
; 
32'd132888: dataIn1 = 32'd2168
; 
32'd132889: dataIn1 = 32'd2169
; 
32'd132890: dataIn1 = 32'd2170
; 
32'd132891: dataIn1 = 32'd2171
; 
32'd132892: dataIn1 = 32'd49
; 
32'd132893: dataIn1 = 32'd50
; 
32'd132894: dataIn1 = 32'd2169
; 
32'd132895: dataIn1 = 32'd2170
; 
32'd132896: dataIn1 = 32'd2171
; 
32'd132897: dataIn1 = 32'd2199
; 
32'd132898: dataIn1 = 32'd2200
; 
32'd132899: dataIn1 = 32'd39
; 
32'd132900: dataIn1 = 32'd50
; 
32'd132901: dataIn1 = 32'd2142
; 
32'd132902: dataIn1 = 32'd2169
; 
32'd132903: dataIn1 = 32'd2170
; 
32'd132904: dataIn1 = 32'd2171
; 
32'd132905: dataIn1 = 32'd2172
; 
32'd132906: dataIn1 = 32'd40
; 
32'd132907: dataIn1 = 32'd50
; 
32'd132908: dataIn1 = 32'd2142
; 
32'd132909: dataIn1 = 32'd2171
; 
32'd132910: dataIn1 = 32'd2172
; 
32'd132911: dataIn1 = 32'd2173
; 
32'd132912: dataIn1 = 32'd2174
; 
32'd132913: dataIn1 = 32'd50
; 
32'd132914: dataIn1 = 32'd51
; 
32'd132915: dataIn1 = 32'd2172
; 
32'd132916: dataIn1 = 32'd2173
; 
32'd132917: dataIn1 = 32'd2174
; 
32'd132918: dataIn1 = 32'd2202
; 
32'd132919: dataIn1 = 32'd2203
; 
32'd132920: dataIn1 = 32'd3618
; 
32'd132921: dataIn1 = 32'd3623
; 
32'd132922: dataIn1 = 32'd40
; 
32'd132923: dataIn1 = 32'd51
; 
32'd132924: dataIn1 = 32'd2145
; 
32'd132925: dataIn1 = 32'd2172
; 
32'd132926: dataIn1 = 32'd2173
; 
32'd132927: dataIn1 = 32'd2174
; 
32'd132928: dataIn1 = 32'd2175
; 
32'd132929: dataIn1 = 32'd9780
; 
32'd132930: dataIn1 = 32'd2145
; 
32'd132931: dataIn1 = 32'd2174
; 
32'd132932: dataIn1 = 32'd2175
; 
32'd132933: dataIn1 = 32'd9770
; 
32'd132934: dataIn1 = 32'd9771
; 
32'd132935: dataIn1 = 32'd9780
; 
32'd132936: dataIn1 = 32'd9781
; 
32'd132937: dataIn1 = 32'd2176
; 
32'd132938: dataIn1 = 32'd3631
; 
32'd132939: dataIn1 = 32'd9471
; 
32'd132940: dataIn1 = 32'd9472
; 
32'd132941: dataIn1 = 32'd9492
; 
32'd132942: dataIn1 = 32'd9493
; 
32'd132943: dataIn1 = 32'd9771
; 
32'd132944: dataIn1 = 32'd9907
; 
32'd132945: dataIn1 = 32'd2177
; 
32'd132946: dataIn1 = 32'd9843
; 
32'd132947: dataIn1 = 32'd9849
; 
32'd132948: dataIn1 = 32'd9862
; 
32'd132949: dataIn1 = 32'd9863
; 
32'd132950: dataIn1 = 32'd9865
; 
32'd132951: dataIn1 = 32'd10161
; 
32'd132952: dataIn1 = 32'd2178
; 
32'd132953: dataIn1 = 32'd3590
; 
32'd132954: dataIn1 = 32'd3591
; 
32'd132955: dataIn1 = 32'd3592
; 
32'd132956: dataIn1 = 32'd3593
; 
32'd132957: dataIn1 = 32'd3595
; 
32'd132958: dataIn1 = 32'd9466
; 
32'd132959: dataIn1 = 32'd2179
; 
32'd132960: dataIn1 = 32'd3593
; 
32'd132961: dataIn1 = 32'd3594
; 
32'd132962: dataIn1 = 32'd3597
; 
32'd132963: dataIn1 = 32'd3599
; 
32'd132964: dataIn1 = 32'd3641
; 
32'd132965: dataIn1 = 32'd3643
; 
32'd132966: dataIn1 = 32'd2180
; 
32'd132967: dataIn1 = 32'd3592
; 
32'd132968: dataIn1 = 32'd3594
; 
32'd132969: dataIn1 = 32'd3596
; 
32'd132970: dataIn1 = 32'd3598
; 
32'd132971: dataIn1 = 32'd3600
; 
32'd132972: dataIn1 = 32'd3601
; 
32'd132973: dataIn1 = 32'd2181
; 
32'd132974: dataIn1 = 32'd3601
; 
32'd132975: dataIn1 = 32'd3602
; 
32'd132976: dataIn1 = 32'd3604
; 
32'd132977: dataIn1 = 32'd3606
; 
32'd132978: dataIn1 = 32'd3607
; 
32'd132979: dataIn1 = 32'd3608
; 
32'd132980: dataIn1 = 32'd54
; 
32'd132981: dataIn1 = 32'd2182
; 
32'd132982: dataIn1 = 32'd3608
; 
32'd132983: dataIn1 = 32'd3609
; 
32'd132984: dataIn1 = 32'd3610
; 
32'd132985: dataIn1 = 32'd3653
; 
32'd132986: dataIn1 = 32'd5309
; 
32'd132987: dataIn1 = 32'd54
; 
32'd132988: dataIn1 = 32'd2154
; 
32'd132989: dataIn1 = 32'd2183
; 
32'd132990: dataIn1 = 32'd2184
; 
32'd132991: dataIn1 = 32'd3607
; 
32'd132992: dataIn1 = 32'd3609
; 
32'd132993: dataIn1 = 32'd5308
; 
32'd132994: dataIn1 = 32'd44
; 
32'd132995: dataIn1 = 32'd54
; 
32'd132996: dataIn1 = 32'd2154
; 
32'd132997: dataIn1 = 32'd2183
; 
32'd132998: dataIn1 = 32'd2184
; 
32'd132999: dataIn1 = 32'd55
; 
32'd133000: dataIn1 = 32'd56
; 
32'd133001: dataIn1 = 32'd2185
; 
32'd133002: dataIn1 = 32'd2186
; 
32'd133003: dataIn1 = 32'd2187
; 
32'd133004: dataIn1 = 32'd2215
; 
32'd133005: dataIn1 = 32'd3657
; 
32'd133006: dataIn1 = 32'd45
; 
32'd133007: dataIn1 = 32'd56
; 
32'd133008: dataIn1 = 32'd2158
; 
32'd133009: dataIn1 = 32'd2185
; 
32'd133010: dataIn1 = 32'd2186
; 
32'd133011: dataIn1 = 32'd2187
; 
32'd133012: dataIn1 = 32'd2188
; 
32'd133013: dataIn1 = 32'd45
; 
32'd133014: dataIn1 = 32'd55
; 
32'd133015: dataIn1 = 32'd2185
; 
32'd133016: dataIn1 = 32'd2186
; 
32'd133017: dataIn1 = 32'd2187
; 
32'd133018: dataIn1 = 32'd46
; 
32'd133019: dataIn1 = 32'd56
; 
32'd133020: dataIn1 = 32'd2158
; 
32'd133021: dataIn1 = 32'd2186
; 
32'd133022: dataIn1 = 32'd2188
; 
32'd133023: dataIn1 = 32'd2189
; 
32'd133024: dataIn1 = 32'd2190
; 
32'd133025: dataIn1 = 32'd56
; 
32'd133026: dataIn1 = 32'd57
; 
32'd133027: dataIn1 = 32'd2188
; 
32'd133028: dataIn1 = 32'd2189
; 
32'd133029: dataIn1 = 32'd2190
; 
32'd133030: dataIn1 = 32'd2218
; 
32'd133031: dataIn1 = 32'd2219
; 
32'd133032: dataIn1 = 32'd9783
; 
32'd133033: dataIn1 = 32'd46
; 
32'd133034: dataIn1 = 32'd57
; 
32'd133035: dataIn1 = 32'd2161
; 
32'd133036: dataIn1 = 32'd2188
; 
32'd133037: dataIn1 = 32'd2189
; 
32'd133038: dataIn1 = 32'd2190
; 
32'd133039: dataIn1 = 32'd2191
; 
32'd133040: dataIn1 = 32'd47
; 
32'd133041: dataIn1 = 32'd57
; 
32'd133042: dataIn1 = 32'd2161
; 
32'd133043: dataIn1 = 32'd2190
; 
32'd133044: dataIn1 = 32'd2191
; 
32'd133045: dataIn1 = 32'd2192
; 
32'd133046: dataIn1 = 32'd2193
; 
32'd133047: dataIn1 = 32'd57
; 
32'd133048: dataIn1 = 32'd58
; 
32'd133049: dataIn1 = 32'd2191
; 
32'd133050: dataIn1 = 32'd2192
; 
32'd133051: dataIn1 = 32'd2193
; 
32'd133052: dataIn1 = 32'd2221
; 
32'd133053: dataIn1 = 32'd2222
; 
32'd133054: dataIn1 = 32'd3662
; 
32'd133055: dataIn1 = 32'd47
; 
32'd133056: dataIn1 = 32'd58
; 
32'd133057: dataIn1 = 32'd2164
; 
32'd133058: dataIn1 = 32'd2191
; 
32'd133059: dataIn1 = 32'd2192
; 
32'd133060: dataIn1 = 32'd2193
; 
32'd133061: dataIn1 = 32'd2194
; 
32'd133062: dataIn1 = 32'd48
; 
32'd133063: dataIn1 = 32'd58
; 
32'd133064: dataIn1 = 32'd2164
; 
32'd133065: dataIn1 = 32'd2193
; 
32'd133066: dataIn1 = 32'd2194
; 
32'd133067: dataIn1 = 32'd2195
; 
32'd133068: dataIn1 = 32'd2196
; 
32'd133069: dataIn1 = 32'd58
; 
32'd133070: dataIn1 = 32'd59
; 
32'd133071: dataIn1 = 32'd2194
; 
32'd133072: dataIn1 = 32'd2195
; 
32'd133073: dataIn1 = 32'd2196
; 
32'd133074: dataIn1 = 32'd2224
; 
32'd133075: dataIn1 = 32'd2225
; 
32'd133076: dataIn1 = 32'd3670
; 
32'd133077: dataIn1 = 32'd3675
; 
32'd133078: dataIn1 = 32'd48
; 
32'd133079: dataIn1 = 32'd59
; 
32'd133080: dataIn1 = 32'd2167
; 
32'd133081: dataIn1 = 32'd2194
; 
32'd133082: dataIn1 = 32'd2195
; 
32'd133083: dataIn1 = 32'd2196
; 
32'd133084: dataIn1 = 32'd2197
; 
32'd133085: dataIn1 = 32'd49
; 
32'd133086: dataIn1 = 32'd59
; 
32'd133087: dataIn1 = 32'd2167
; 
32'd133088: dataIn1 = 32'd2196
; 
32'd133089: dataIn1 = 32'd2197
; 
32'd133090: dataIn1 = 32'd2198
; 
32'd133091: dataIn1 = 32'd2199
; 
32'd133092: dataIn1 = 32'd3683
; 
32'd133093: dataIn1 = 32'd2197
; 
32'd133094: dataIn1 = 32'd2198
; 
32'd133095: dataIn1 = 32'd2199
; 
32'd133096: dataIn1 = 32'd3680
; 
32'd133097: dataIn1 = 32'd3682
; 
32'd133098: dataIn1 = 32'd3683
; 
32'd133099: dataIn1 = 32'd3685
; 
32'd133100: dataIn1 = 32'd49
; 
32'd133101: dataIn1 = 32'd60
; 
32'd133102: dataIn1 = 32'd2170
; 
32'd133103: dataIn1 = 32'd2197
; 
32'd133104: dataIn1 = 32'd2198
; 
32'd133105: dataIn1 = 32'd2199
; 
32'd133106: dataIn1 = 32'd2200
; 
32'd133107: dataIn1 = 32'd3614
; 
32'd133108: dataIn1 = 32'd3685
; 
32'd133109: dataIn1 = 32'd50
; 
32'd133110: dataIn1 = 32'd2170
; 
32'd133111: dataIn1 = 32'd2199
; 
32'd133112: dataIn1 = 32'd2200
; 
32'd133113: dataIn1 = 32'd3611
; 
32'd133114: dataIn1 = 32'd3612
; 
32'd133115: dataIn1 = 32'd3614
; 
32'd133116: dataIn1 = 32'd2201
; 
32'd133117: dataIn1 = 32'd3612
; 
32'd133118: dataIn1 = 32'd3613
; 
32'd133119: dataIn1 = 32'd3615
; 
32'd133120: dataIn1 = 32'd3617
; 
32'd133121: dataIn1 = 32'd3694
; 
32'd133122: dataIn1 = 32'd3696
; 
32'd133123: dataIn1 = 32'd9538
; 
32'd133124: dataIn1 = 32'd9546
; 
32'd133125: dataIn1 = 32'd50
; 
32'd133126: dataIn1 = 32'd2173
; 
32'd133127: dataIn1 = 32'd2202
; 
32'd133128: dataIn1 = 32'd3611
; 
32'd133129: dataIn1 = 32'd3613
; 
32'd133130: dataIn1 = 32'd3616
; 
32'd133131: dataIn1 = 32'd3618
; 
32'd133132: dataIn1 = 32'd2173
; 
32'd133133: dataIn1 = 32'd2203
; 
32'd133134: dataIn1 = 32'd3618
; 
32'd133135: dataIn1 = 32'd3619
; 
32'd133136: dataIn1 = 32'd3620
; 
32'd133137: dataIn1 = 32'd3621
; 
32'd133138: dataIn1 = 32'd3623
; 
32'd133139: dataIn1 = 32'd9480
; 
32'd133140: dataIn1 = 32'd10165
; 
32'd133141: dataIn1 = 32'd2204
; 
32'd133142: dataIn1 = 32'd3708
; 
32'd133143: dataIn1 = 32'd9481
; 
32'd133144: dataIn1 = 32'd9482
; 
32'd133145: dataIn1 = 32'd9486
; 
32'd133146: dataIn1 = 32'd9557
; 
32'd133147: dataIn1 = 32'd9870
; 
32'd133148: dataIn1 = 32'd9878
; 
32'd133149: dataIn1 = 32'd10163
; 
32'd133150: dataIn1 = 32'd2205
; 
32'd133151: dataIn1 = 32'd9484
; 
32'd133152: dataIn1 = 32'd9887
; 
32'd133153: dataIn1 = 32'd9888
; 
32'd133154: dataIn1 = 32'd9903
; 
32'd133155: dataIn1 = 32'd9904
; 
32'd133156: dataIn1 = 32'd10169
; 
32'd133157: dataIn1 = 32'd2206
; 
32'd133158: dataIn1 = 32'd3632
; 
32'd133159: dataIn1 = 32'd3634
; 
32'd133160: dataIn1 = 32'd3635
; 
32'd133161: dataIn1 = 32'd10167
; 
32'd133162: dataIn1 = 32'd10168
; 
32'd133163: dataIn1 = 32'd10228
; 
32'd133164: dataIn1 = 32'd2207
; 
32'd133165: dataIn1 = 32'd3635
; 
32'd133166: dataIn1 = 32'd3636
; 
32'd133167: dataIn1 = 32'd3638
; 
32'd133168: dataIn1 = 32'd3640
; 
32'd133169: dataIn1 = 32'd3718
; 
32'd133170: dataIn1 = 32'd3720
; 
32'd133171: dataIn1 = 32'd2208
; 
32'd133172: dataIn1 = 32'd3634
; 
32'd133173: dataIn1 = 32'd3636
; 
32'd133174: dataIn1 = 32'd3637
; 
32'd133175: dataIn1 = 32'd3639
; 
32'd133176: dataIn1 = 32'd3641
; 
32'd133177: dataIn1 = 32'd3642
; 
32'd133178: dataIn1 = 32'd2209
; 
32'd133179: dataIn1 = 32'd3642
; 
32'd133180: dataIn1 = 32'd3643
; 
32'd133181: dataIn1 = 32'd3644
; 
32'd133182: dataIn1 = 32'd3645
; 
32'd133183: dataIn1 = 32'd3646
; 
32'd133184: dataIn1 = 32'd3647
; 
32'd133185: dataIn1 = 32'd2210
; 
32'd133186: dataIn1 = 32'd3647
; 
32'd133187: dataIn1 = 32'd3648
; 
32'd133188: dataIn1 = 32'd3650
; 
32'd133189: dataIn1 = 32'd3652
; 
32'd133190: dataIn1 = 32'd3728
; 
32'd133191: dataIn1 = 32'd3730
; 
32'd133192: dataIn1 = 32'd2211
; 
32'd133193: dataIn1 = 32'd3646
; 
32'd133194: dataIn1 = 32'd3648
; 
32'd133195: dataIn1 = 32'd3649
; 
32'd133196: dataIn1 = 32'd3651
; 
32'd133197: dataIn1 = 32'd3653
; 
32'd133198: dataIn1 = 32'd3654
; 
32'd133199: dataIn1 = 32'd54
; 
32'd133200: dataIn1 = 32'd2212
; 
32'd133201: dataIn1 = 32'd2213
; 
32'd133202: dataIn1 = 32'd2214
; 
32'd133203: dataIn1 = 32'd3654
; 
32'd133204: dataIn1 = 32'd3655
; 
32'd133205: dataIn1 = 32'd5309
; 
32'd133206: dataIn1 = 32'd64
; 
32'd133207: dataIn1 = 32'd65
; 
32'd133208: dataIn1 = 32'd2212
; 
32'd133209: dataIn1 = 32'd2213
; 
32'd133210: dataIn1 = 32'd2214
; 
32'd133211: dataIn1 = 32'd3655
; 
32'd133212: dataIn1 = 32'd5312
; 
32'd133213: dataIn1 = 32'd5455
; 
32'd133214: dataIn1 = 32'd54
; 
32'd133215: dataIn1 = 32'd65
; 
32'd133216: dataIn1 = 32'd2212
; 
32'd133217: dataIn1 = 32'd2213
; 
32'd133218: dataIn1 = 32'd2214
; 
32'd133219: dataIn1 = 32'd56
; 
32'd133220: dataIn1 = 32'd2185
; 
32'd133221: dataIn1 = 32'd2215
; 
32'd133222: dataIn1 = 32'd3657
; 
32'd133223: dataIn1 = 32'd3658
; 
32'd133224: dataIn1 = 32'd5310
; 
32'd133225: dataIn1 = 32'd9782
; 
32'd133226: dataIn1 = 32'd55
; 
32'd133227: dataIn1 = 32'd2216
; 
32'd133228: dataIn1 = 32'd3656
; 
32'd133229: dataIn1 = 32'd3657
; 
32'd133230: dataIn1 = 32'd2217
; 
32'd133231: dataIn1 = 32'd5310
; 
32'd133232: dataIn1 = 32'd9568
; 
32'd133233: dataIn1 = 32'd10039
; 
32'd133234: dataIn1 = 32'd10040
; 
32'd133235: dataIn1 = 32'd10057
; 
32'd133236: dataIn1 = 32'd10204
; 
32'd133237: dataIn1 = 32'd56
; 
32'd133238: dataIn1 = 32'd2189
; 
32'd133239: dataIn1 = 32'd2218
; 
32'd133240: dataIn1 = 32'd9772
; 
32'd133241: dataIn1 = 32'd9773
; 
32'd133242: dataIn1 = 32'd9782
; 
32'd133243: dataIn1 = 32'd9783
; 
32'd133244: dataIn1 = 32'd10238
; 
32'd133245: dataIn1 = 32'd57
; 
32'd133246: dataIn1 = 32'd2189
; 
32'd133247: dataIn1 = 32'd2219
; 
32'd133248: dataIn1 = 32'd9774
; 
32'd133249: dataIn1 = 32'd9775
; 
32'd133250: dataIn1 = 32'd9783
; 
32'd133251: dataIn1 = 32'd9784
; 
32'd133252: dataIn1 = 32'd10240
; 
32'd133253: dataIn1 = 32'd2220
; 
32'd133254: dataIn1 = 32'd10066
; 
32'd133255: dataIn1 = 32'd10068
; 
32'd133256: dataIn1 = 32'd10080
; 
32'd133257: dataIn1 = 32'd10089
; 
32'd133258: dataIn1 = 32'd10210
; 
32'd133259: dataIn1 = 32'd10212
; 
32'd133260: dataIn1 = 32'd57
; 
32'd133261: dataIn1 = 32'd2192
; 
32'd133262: dataIn1 = 32'd2221
; 
32'd133263: dataIn1 = 32'd3659
; 
32'd133264: dataIn1 = 32'd3661
; 
32'd133265: dataIn1 = 32'd3662
; 
32'd133266: dataIn1 = 32'd9784
; 
32'd133267: dataIn1 = 32'd10242
; 
32'd133268: dataIn1 = 32'd58
; 
32'd133269: dataIn1 = 32'd2192
; 
32'd133270: dataIn1 = 32'd2222
; 
32'd133271: dataIn1 = 32'd3662
; 
32'd133272: dataIn1 = 32'd3663
; 
32'd133273: dataIn1 = 32'd3664
; 
32'd133274: dataIn1 = 32'd3665
; 
32'd133275: dataIn1 = 32'd10244
; 
32'd133276: dataIn1 = 32'd2223
; 
32'd133277: dataIn1 = 32'd9501
; 
32'd133278: dataIn1 = 32'd10098
; 
32'd133279: dataIn1 = 32'd10100
; 
32'd133280: dataIn1 = 32'd10112
; 
32'd133281: dataIn1 = 32'd10118
; 
32'd133282: dataIn1 = 32'd10218
; 
32'd133283: dataIn1 = 32'd58
; 
32'd133284: dataIn1 = 32'd2195
; 
32'd133285: dataIn1 = 32'd2224
; 
32'd133286: dataIn1 = 32'd3664
; 
32'd133287: dataIn1 = 32'd3666
; 
32'd133288: dataIn1 = 32'd3668
; 
32'd133289: dataIn1 = 32'd3670
; 
32'd133290: dataIn1 = 32'd9499
; 
32'd133291: dataIn1 = 32'd2195
; 
32'd133292: dataIn1 = 32'd2225
; 
32'd133293: dataIn1 = 32'd3670
; 
32'd133294: dataIn1 = 32'd3671
; 
32'd133295: dataIn1 = 32'd3672
; 
32'd133296: dataIn1 = 32'd3673
; 
32'd133297: dataIn1 = 32'd3675
; 
32'd133298: dataIn1 = 32'd9512
; 
32'd133299: dataIn1 = 32'd10176
; 
32'd133300: dataIn1 = 32'd2226
; 
32'd133301: dataIn1 = 32'd3782
; 
32'd133302: dataIn1 = 32'd9518
; 
32'd133303: dataIn1 = 32'd9927
; 
32'd133304: dataIn1 = 32'd9928
; 
32'd133305: dataIn1 = 32'd9937
; 
32'd133306: dataIn1 = 32'd10178
; 
32'd133307: dataIn1 = 32'd2227
; 
32'd133308: dataIn1 = 32'd3676
; 
32'd133309: dataIn1 = 32'd3680
; 
32'd133310: dataIn1 = 32'd10181
; 
32'd133311: dataIn1 = 32'd10182
; 
32'd133312: dataIn1 = 32'd10231
; 
32'd133313: dataIn1 = 32'd10233
; 
32'd133314: dataIn1 = 32'd2228
; 
32'd133315: dataIn1 = 32'd3682
; 
32'd133316: dataIn1 = 32'd3686
; 
32'd133317: dataIn1 = 32'd9524
; 
32'd133318: dataIn1 = 32'd9525
; 
32'd133319: dataIn1 = 32'd9532
; 
32'd133320: dataIn1 = 32'd9533
; 
32'd133321: dataIn1 = 32'd9981
; 
32'd133322: dataIn1 = 32'd2229
; 
32'd133323: dataIn1 = 32'd3693
; 
32'd133324: dataIn1 = 32'd3792
; 
32'd133325: dataIn1 = 32'd3794
; 
32'd133326: dataIn1 = 32'd10185
; 
32'd133327: dataIn1 = 32'd10186
; 
32'd133328: dataIn1 = 32'd10234
; 
32'd133329: dataIn1 = 32'd2230
; 
32'd133330: dataIn1 = 32'd9975
; 
32'd133331: dataIn1 = 32'd9976
; 
32'd133332: dataIn1 = 32'd9984
; 
32'd133333: dataIn1 = 32'd9999
; 
32'd133334: dataIn1 = 32'd10000
; 
32'd133335: dataIn1 = 32'd10187
; 
32'd133336: dataIn1 = 32'd2231
; 
32'd133337: dataIn1 = 32'd3700
; 
32'd133338: dataIn1 = 32'd9540
; 
32'd133339: dataIn1 = 32'd9541
; 
32'd133340: dataIn1 = 32'd9548
; 
32'd133341: dataIn1 = 32'd9989
; 
32'd133342: dataIn1 = 32'd10005
; 
32'd133343: dataIn1 = 32'd10191
; 
32'd133344: dataIn1 = 32'd10193
; 
32'd133345: dataIn1 = 32'd2232
; 
32'd133346: dataIn1 = 32'd3700
; 
32'd133347: dataIn1 = 32'd3701
; 
32'd133348: dataIn1 = 32'd3703
; 
32'd133349: dataIn1 = 32'd3705
; 
32'd133350: dataIn1 = 32'd3804
; 
32'd133351: dataIn1 = 32'd3806
; 
32'd133352: dataIn1 = 32'd2233
; 
32'd133353: dataIn1 = 32'd3699
; 
32'd133354: dataIn1 = 32'd3701
; 
32'd133355: dataIn1 = 32'd3702
; 
32'd133356: dataIn1 = 32'd3704
; 
32'd133357: dataIn1 = 32'd3706
; 
32'd133358: dataIn1 = 32'd3707
; 
32'd133359: dataIn1 = 32'd9555
; 
32'd133360: dataIn1 = 32'd10195
; 
32'd133361: dataIn1 = 32'd2234
; 
32'd133362: dataIn1 = 32'd3707
; 
32'd133363: dataIn1 = 32'd3708
; 
32'd133364: dataIn1 = 32'd3709
; 
32'd133365: dataIn1 = 32'd3710
; 
32'd133366: dataIn1 = 32'd3711
; 
32'd133367: dataIn1 = 32'd3712
; 
32'd133368: dataIn1 = 32'd2235
; 
32'd133369: dataIn1 = 32'd3712
; 
32'd133370: dataIn1 = 32'd3713
; 
32'd133371: dataIn1 = 32'd3715
; 
32'd133372: dataIn1 = 32'd3717
; 
32'd133373: dataIn1 = 32'd3816
; 
32'd133374: dataIn1 = 32'd3818
; 
32'd133375: dataIn1 = 32'd2236
; 
32'd133376: dataIn1 = 32'd3711
; 
32'd133377: dataIn1 = 32'd3713
; 
32'd133378: dataIn1 = 32'd3714
; 
32'd133379: dataIn1 = 32'd3716
; 
32'd133380: dataIn1 = 32'd3718
; 
32'd133381: dataIn1 = 32'd3719
; 
32'd133382: dataIn1 = 32'd2237
; 
32'd133383: dataIn1 = 32'd3719
; 
32'd133384: dataIn1 = 32'd3720
; 
32'd133385: dataIn1 = 32'd3721
; 
32'd133386: dataIn1 = 32'd3722
; 
32'd133387: dataIn1 = 32'd3723
; 
32'd133388: dataIn1 = 32'd3724
; 
32'd133389: dataIn1 = 32'd74
; 
32'd133390: dataIn1 = 32'd2238
; 
32'd133391: dataIn1 = 32'd2264
; 
32'd133392: dataIn1 = 32'd2265
; 
32'd133393: dataIn1 = 32'd3724
; 
32'd133394: dataIn1 = 32'd3725
; 
32'd133395: dataIn1 = 32'd3727
; 
32'd133396: dataIn1 = 32'd74
; 
32'd133397: dataIn1 = 32'd2239
; 
32'd133398: dataIn1 = 32'd3723
; 
32'd133399: dataIn1 = 32'd3725
; 
32'd133400: dataIn1 = 32'd3726
; 
32'd133401: dataIn1 = 32'd3728
; 
32'd133402: dataIn1 = 32'd3729
; 
32'd133403: dataIn1 = 32'd74
; 
32'd133404: dataIn1 = 32'd2240
; 
32'd133405: dataIn1 = 32'd3729
; 
32'd133406: dataIn1 = 32'd3730
; 
32'd133407: dataIn1 = 32'd3731
; 
32'd133408: dataIn1 = 32'd5311
; 
32'd133409: dataIn1 = 32'd5312
; 
32'd133410: dataIn1 = 32'd2241
; 
32'd133411: dataIn1 = 32'd3733
; 
32'd133412: dataIn1 = 32'd3734
; 
32'd133413: dataIn1 = 32'd3738
; 
32'd133414: dataIn1 = 32'd3740
; 
32'd133415: dataIn1 = 32'd3821
; 
32'd133416: dataIn1 = 32'd3823
; 
32'd133417: dataIn1 = 32'd2242
; 
32'd133418: dataIn1 = 32'd3734
; 
32'd133419: dataIn1 = 32'd3739
; 
32'd133420: dataIn1 = 32'd10201
; 
32'd133421: dataIn1 = 32'd10202
; 
32'd133422: dataIn1 = 32'd10236
; 
32'd133423: dataIn1 = 32'd10237
; 
32'd133424: dataIn1 = 32'd2243
; 
32'd133425: dataIn1 = 32'd3732
; 
32'd133426: dataIn1 = 32'd3733
; 
32'd133427: dataIn1 = 32'd3737
; 
32'd133428: dataIn1 = 32'd10198
; 
32'd133429: dataIn1 = 32'd10287
; 
32'd133430: dataIn1 = 32'd2244
; 
32'd133431: dataIn1 = 32'd3742
; 
32'd133432: dataIn1 = 32'd3743
; 
32'd133433: dataIn1 = 32'd3745
; 
32'd133434: dataIn1 = 32'd3747
; 
32'd133435: dataIn1 = 32'd3748
; 
32'd133436: dataIn1 = 32'd3749
; 
32'd133437: dataIn1 = 32'd9569
; 
32'd133438: dataIn1 = 32'd10199
; 
32'd133439: dataIn1 = 32'd2245
; 
32'd133440: dataIn1 = 32'd3749
; 
32'd133441: dataIn1 = 32'd3750
; 
32'd133442: dataIn1 = 32'd3752
; 
32'd133443: dataIn1 = 32'd3754
; 
32'd133444: dataIn1 = 32'd3831
; 
32'd133445: dataIn1 = 32'd3833
; 
32'd133446: dataIn1 = 32'd2246
; 
32'd133447: dataIn1 = 32'd3748
; 
32'd133448: dataIn1 = 32'd3750
; 
32'd133449: dataIn1 = 32'd3751
; 
32'd133450: dataIn1 = 32'd3753
; 
32'd133451: dataIn1 = 32'd3755
; 
32'd133452: dataIn1 = 32'd3756
; 
32'd133453: dataIn1 = 32'd9582
; 
32'd133454: dataIn1 = 32'd2247
; 
32'd133455: dataIn1 = 32'd3756
; 
32'd133456: dataIn1 = 32'd3757
; 
32'd133457: dataIn1 = 32'd3759
; 
32'd133458: dataIn1 = 32'd3760
; 
32'd133459: dataIn1 = 32'd3761
; 
32'd133460: dataIn1 = 32'd3762
; 
32'd133461: dataIn1 = 32'd9585
; 
32'd133462: dataIn1 = 32'd2248
; 
32'd133463: dataIn1 = 32'd3762
; 
32'd133464: dataIn1 = 32'd3763
; 
32'd133465: dataIn1 = 32'd3765
; 
32'd133466: dataIn1 = 32'd3767
; 
32'd133467: dataIn1 = 32'd3843
; 
32'd133468: dataIn1 = 32'd3845
; 
32'd133469: dataIn1 = 32'd2249
; 
32'd133470: dataIn1 = 32'd3761
; 
32'd133471: dataIn1 = 32'd3763
; 
32'd133472: dataIn1 = 32'd3764
; 
32'd133473: dataIn1 = 32'd3766
; 
32'd133474: dataIn1 = 32'd3768
; 
32'd133475: dataIn1 = 32'd3769
; 
32'd133476: dataIn1 = 32'd9598
; 
32'd133477: dataIn1 = 32'd2250
; 
32'd133478: dataIn1 = 32'd3769
; 
32'd133479: dataIn1 = 32'd3770
; 
32'd133480: dataIn1 = 32'd3771
; 
32'd133481: dataIn1 = 32'd3772
; 
32'd133482: dataIn1 = 32'd3773
; 
32'd133483: dataIn1 = 32'd3774
; 
32'd133484: dataIn1 = 32'd10219
; 
32'd133485: dataIn1 = 32'd2251
; 
32'd133486: dataIn1 = 32'd3774
; 
32'd133487: dataIn1 = 32'd3775
; 
32'd133488: dataIn1 = 32'd3777
; 
32'd133489: dataIn1 = 32'd3779
; 
32'd133490: dataIn1 = 32'd3850
; 
32'd133491: dataIn1 = 32'd3852
; 
32'd133492: dataIn1 = 32'd2252
; 
32'd133493: dataIn1 = 32'd3773
; 
32'd133494: dataIn1 = 32'd3775
; 
32'd133495: dataIn1 = 32'd3776
; 
32'd133496: dataIn1 = 32'd3778
; 
32'd133497: dataIn1 = 32'd3780
; 
32'd133498: dataIn1 = 32'd3781
; 
32'd133499: dataIn1 = 32'd10232
; 
32'd133500: dataIn1 = 32'd2253
; 
32'd133501: dataIn1 = 32'd3781
; 
32'd133502: dataIn1 = 32'd3782
; 
32'd133503: dataIn1 = 32'd3783
; 
32'd133504: dataIn1 = 32'd3784
; 
32'd133505: dataIn1 = 32'd3785
; 
32'd133506: dataIn1 = 32'd3786
; 
32'd133507: dataIn1 = 32'd2254
; 
32'd133508: dataIn1 = 32'd3786
; 
32'd133509: dataIn1 = 32'd3787
; 
32'd133510: dataIn1 = 32'd3789
; 
32'd133511: dataIn1 = 32'd3791
; 
32'd133512: dataIn1 = 32'd3856
; 
32'd133513: dataIn1 = 32'd3858
; 
32'd133514: dataIn1 = 32'd2255
; 
32'd133515: dataIn1 = 32'd3785
; 
32'd133516: dataIn1 = 32'd3787
; 
32'd133517: dataIn1 = 32'd3788
; 
32'd133518: dataIn1 = 32'd3790
; 
32'd133519: dataIn1 = 32'd3792
; 
32'd133520: dataIn1 = 32'd3793
; 
32'd133521: dataIn1 = 32'd2256
; 
32'd133522: dataIn1 = 32'd3793
; 
32'd133523: dataIn1 = 32'd3794
; 
32'd133524: dataIn1 = 32'd3795
; 
32'd133525: dataIn1 = 32'd3796
; 
32'd133526: dataIn1 = 32'd3797
; 
32'd133527: dataIn1 = 32'd3798
; 
32'd133528: dataIn1 = 32'd2257
; 
32'd133529: dataIn1 = 32'd2282
; 
32'd133530: dataIn1 = 32'd3798
; 
32'd133531: dataIn1 = 32'd3799
; 
32'd133532: dataIn1 = 32'd3801
; 
32'd133533: dataIn1 = 32'd3803
; 
32'd133534: dataIn1 = 32'd3862
; 
32'd133535: dataIn1 = 32'd2258
; 
32'd133536: dataIn1 = 32'd3797
; 
32'd133537: dataIn1 = 32'd3799
; 
32'd133538: dataIn1 = 32'd3800
; 
32'd133539: dataIn1 = 32'd3802
; 
32'd133540: dataIn1 = 32'd3804
; 
32'd133541: dataIn1 = 32'd3805
; 
32'd133542: dataIn1 = 32'd2259
; 
32'd133543: dataIn1 = 32'd3805
; 
32'd133544: dataIn1 = 32'd3806
; 
32'd133545: dataIn1 = 32'd3807
; 
32'd133546: dataIn1 = 32'd3808
; 
32'd133547: dataIn1 = 32'd3809
; 
32'd133548: dataIn1 = 32'd3810
; 
32'd133549: dataIn1 = 32'd2260
; 
32'd133550: dataIn1 = 32'd2284
; 
32'd133551: dataIn1 = 32'd2285
; 
32'd133552: dataIn1 = 32'd3810
; 
32'd133553: dataIn1 = 32'd3811
; 
32'd133554: dataIn1 = 32'd3813
; 
32'd133555: dataIn1 = 32'd3815
; 
32'd133556: dataIn1 = 32'd2261
; 
32'd133557: dataIn1 = 32'd3809
; 
32'd133558: dataIn1 = 32'd3811
; 
32'd133559: dataIn1 = 32'd3812
; 
32'd133560: dataIn1 = 32'd3814
; 
32'd133561: dataIn1 = 32'd3816
; 
32'd133562: dataIn1 = 32'd3817
; 
32'd133563: dataIn1 = 32'd2262
; 
32'd133564: dataIn1 = 32'd2263
; 
32'd133565: dataIn1 = 32'd2264
; 
32'd133566: dataIn1 = 32'd3817
; 
32'd133567: dataIn1 = 32'd3818
; 
32'd133568: dataIn1 = 32'd3819
; 
32'd133569: dataIn1 = 32'd3820
; 
32'd133570: dataIn1 = 32'd83
; 
32'd133571: dataIn1 = 32'd84
; 
32'd133572: dataIn1 = 32'd94
; 
32'd133573: dataIn1 = 32'd2262
; 
32'd133574: dataIn1 = 32'd2263
; 
32'd133575: dataIn1 = 32'd2264
; 
32'd133576: dataIn1 = 32'd3819
; 
32'd133577: dataIn1 = 32'd73
; 
32'd133578: dataIn1 = 32'd84
; 
32'd133579: dataIn1 = 32'd2238
; 
32'd133580: dataIn1 = 32'd2262
; 
32'd133581: dataIn1 = 32'd2263
; 
32'd133582: dataIn1 = 32'd2264
; 
32'd133583: dataIn1 = 32'd2265
; 
32'd133584: dataIn1 = 32'd3727
; 
32'd133585: dataIn1 = 32'd3820
; 
32'd133586: dataIn1 = 32'd74
; 
32'd133587: dataIn1 = 32'd84
; 
32'd133588: dataIn1 = 32'd85
; 
32'd133589: dataIn1 = 32'd2238
; 
32'd133590: dataIn1 = 32'd2264
; 
32'd133591: dataIn1 = 32'd2265
; 
32'd133592: dataIn1 = 32'd87
; 
32'd133593: dataIn1 = 32'd2266
; 
32'd133594: dataIn1 = 32'd3822
; 
32'd133595: dataIn1 = 32'd3823
; 
32'd133596: dataIn1 = 32'd3825
; 
32'd133597: dataIn1 = 32'd3826
; 
32'd133598: dataIn1 = 32'd5313
; 
32'd133599: dataIn1 = 32'd87
; 
32'd133600: dataIn1 = 32'd2267
; 
32'd133601: dataIn1 = 32'd3821
; 
32'd133602: dataIn1 = 32'd3822
; 
32'd133603: dataIn1 = 32'd3824
; 
32'd133604: dataIn1 = 32'd87
; 
32'd133605: dataIn1 = 32'd2268
; 
32'd133606: dataIn1 = 32'd3829
; 
32'd133607: dataIn1 = 32'd3830
; 
32'd133608: dataIn1 = 32'd5313
; 
32'd133609: dataIn1 = 32'd5314
; 
32'd133610: dataIn1 = 32'd5315
; 
32'd133611: dataIn1 = 32'd2269
; 
32'd133612: dataIn1 = 32'd3826
; 
32'd133613: dataIn1 = 32'd3827
; 
32'd133614: dataIn1 = 32'd3828
; 
32'd133615: dataIn1 = 32'd3830
; 
32'd133616: dataIn1 = 32'd3831
; 
32'd133617: dataIn1 = 32'd3832
; 
32'd133618: dataIn1 = 32'd2270
; 
32'd133619: dataIn1 = 32'd3832
; 
32'd133620: dataIn1 = 32'd3833
; 
32'd133621: dataIn1 = 32'd3834
; 
32'd133622: dataIn1 = 32'd3835
; 
32'd133623: dataIn1 = 32'd3836
; 
32'd133624: dataIn1 = 32'd3838
; 
32'd133625: dataIn1 = 32'd2271
; 
32'd133626: dataIn1 = 32'd3838
; 
32'd133627: dataIn1 = 32'd3839
; 
32'd133628: dataIn1 = 32'd3841
; 
32'd133629: dataIn1 = 32'd3842
; 
32'd133630: dataIn1 = 32'd5316
; 
32'd133631: dataIn1 = 32'd5317
; 
32'd133632: dataIn1 = 32'd2272
; 
32'd133633: dataIn1 = 32'd3836
; 
32'd133634: dataIn1 = 32'd3837
; 
32'd133635: dataIn1 = 32'd3840
; 
32'd133636: dataIn1 = 32'd3842
; 
32'd133637: dataIn1 = 32'd3843
; 
32'd133638: dataIn1 = 32'd3844
; 
32'd133639: dataIn1 = 32'd2273
; 
32'd133640: dataIn1 = 32'd2274
; 
32'd133641: dataIn1 = 32'd3844
; 
32'd133642: dataIn1 = 32'd3845
; 
32'd133643: dataIn1 = 32'd3846
; 
32'd133644: dataIn1 = 32'd3847
; 
32'd133645: dataIn1 = 32'd3848
; 
32'd133646: dataIn1 = 32'd89
; 
32'd133647: dataIn1 = 32'd90
; 
32'd133648: dataIn1 = 32'd100
; 
32'd133649: dataIn1 = 32'd2273
; 
32'd133650: dataIn1 = 32'd2274
; 
32'd133651: dataIn1 = 32'd2275
; 
32'd133652: dataIn1 = 32'd3846
; 
32'd133653: dataIn1 = 32'd3848
; 
32'd133654: dataIn1 = 32'd90
; 
32'd133655: dataIn1 = 32'd2274
; 
32'd133656: dataIn1 = 32'd2275
; 
32'd133657: dataIn1 = 32'd3848
; 
32'd133658: dataIn1 = 32'd3849
; 
32'd133659: dataIn1 = 32'd3850
; 
32'd133660: dataIn1 = 32'd3851
; 
32'd133661: dataIn1 = 32'd90
; 
32'd133662: dataIn1 = 32'd2276
; 
32'd133663: dataIn1 = 32'd2277
; 
32'd133664: dataIn1 = 32'd3851
; 
32'd133665: dataIn1 = 32'd3852
; 
32'd133666: dataIn1 = 32'd3853
; 
32'd133667: dataIn1 = 32'd3854
; 
32'd133668: dataIn1 = 32'd90
; 
32'd133669: dataIn1 = 32'd91
; 
32'd133670: dataIn1 = 32'd101
; 
32'd133671: dataIn1 = 32'd2276
; 
32'd133672: dataIn1 = 32'd2277
; 
32'd133673: dataIn1 = 32'd2278
; 
32'd133674: dataIn1 = 32'd3854
; 
32'd133675: dataIn1 = 32'd91
; 
32'd133676: dataIn1 = 32'd2277
; 
32'd133677: dataIn1 = 32'd2278
; 
32'd133678: dataIn1 = 32'd3854
; 
32'd133679: dataIn1 = 32'd3855
; 
32'd133680: dataIn1 = 32'd3856
; 
32'd133681: dataIn1 = 32'd3857
; 
32'd133682: dataIn1 = 32'd91
; 
32'd133683: dataIn1 = 32'd2279
; 
32'd133684: dataIn1 = 32'd2280
; 
32'd133685: dataIn1 = 32'd3857
; 
32'd133686: dataIn1 = 32'd3858
; 
32'd133687: dataIn1 = 32'd3859
; 
32'd133688: dataIn1 = 32'd3860
; 
32'd133689: dataIn1 = 32'd91
; 
32'd133690: dataIn1 = 32'd92
; 
32'd133691: dataIn1 = 32'd102
; 
32'd133692: dataIn1 = 32'd2279
; 
32'd133693: dataIn1 = 32'd2280
; 
32'd133694: dataIn1 = 32'd2281
; 
32'd133695: dataIn1 = 32'd3860
; 
32'd133696: dataIn1 = 32'd92
; 
32'd133697: dataIn1 = 32'd2280
; 
32'd133698: dataIn1 = 32'd2281
; 
32'd133699: dataIn1 = 32'd2282
; 
32'd133700: dataIn1 = 32'd3860
; 
32'd133701: dataIn1 = 32'd3861
; 
32'd133702: dataIn1 = 32'd3862
; 
32'd133703: dataIn1 = 32'd82
; 
32'd133704: dataIn1 = 32'd92
; 
32'd133705: dataIn1 = 32'd2257
; 
32'd133706: dataIn1 = 32'd2281
; 
32'd133707: dataIn1 = 32'd2282
; 
32'd133708: dataIn1 = 32'd2283
; 
32'd133709: dataIn1 = 32'd2284
; 
32'd133710: dataIn1 = 32'd3803
; 
32'd133711: dataIn1 = 32'd3862
; 
32'd133712: dataIn1 = 32'd92
; 
32'd133713: dataIn1 = 32'd93
; 
32'd133714: dataIn1 = 32'd103
; 
32'd133715: dataIn1 = 32'd2282
; 
32'd133716: dataIn1 = 32'd2283
; 
32'd133717: dataIn1 = 32'd2284
; 
32'd133718: dataIn1 = 32'd82
; 
32'd133719: dataIn1 = 32'd93
; 
32'd133720: dataIn1 = 32'd2260
; 
32'd133721: dataIn1 = 32'd2282
; 
32'd133722: dataIn1 = 32'd2283
; 
32'd133723: dataIn1 = 32'd2284
; 
32'd133724: dataIn1 = 32'd2285
; 
32'd133725: dataIn1 = 32'd3813
; 
32'd133726: dataIn1 = 32'd83
; 
32'd133727: dataIn1 = 32'd93
; 
32'd133728: dataIn1 = 32'd94
; 
32'd133729: dataIn1 = 32'd2260
; 
32'd133730: dataIn1 = 32'd2284
; 
32'd133731: dataIn1 = 32'd2285
; 
32'd133732: dataIn1 = 32'd3815
; 
32'd133733: dataIn1 = 32'd392
; 
32'd133734: dataIn1 = 32'd2286
; 
32'd133735: dataIn1 = 32'd2289
; 
32'd133736: dataIn1 = 32'd3863
; 
32'd133737: dataIn1 = 32'd3865
; 
32'd133738: dataIn1 = 32'd3867
; 
32'd133739: dataIn1 = 32'd10272
; 
32'd133740: dataIn1 = 32'd2287
; 
32'd133741: dataIn1 = 32'd3863
; 
32'd133742: dataIn1 = 32'd3864
; 
32'd133743: dataIn1 = 32'd4607
; 
32'd133744: dataIn1 = 32'd4608
; 
32'd133745: dataIn1 = 32'd4611
; 
32'd133746: dataIn1 = 32'd10263
; 
32'd133747: dataIn1 = 32'd2288
; 
32'd133748: dataIn1 = 32'd2289
; 
32'd133749: dataIn1 = 32'd3866
; 
32'd133750: dataIn1 = 32'd3867
; 
32'd133751: dataIn1 = 32'd5689
; 
32'd133752: dataIn1 = 32'd5690
; 
32'd133753: dataIn1 = 32'd5692
; 
32'd133754: dataIn1 = 32'd392
; 
32'd133755: dataIn1 = 32'd400
; 
32'd133756: dataIn1 = 32'd761
; 
32'd133757: dataIn1 = 32'd2286
; 
32'd133758: dataIn1 = 32'd2288
; 
32'd133759: dataIn1 = 32'd2289
; 
32'd133760: dataIn1 = 32'd2489
; 
32'd133761: dataIn1 = 32'd3867
; 
32'd133762: dataIn1 = 32'd5692
; 
32'd133763: dataIn1 = 32'd206
; 
32'd133764: dataIn1 = 32'd403
; 
32'd133765: dataIn1 = 32'd763
; 
32'd133766: dataIn1 = 32'd2290
; 
32'd133767: dataIn1 = 32'd2291
; 
32'd133768: dataIn1 = 32'd2292
; 
32'd133769: dataIn1 = 32'd2293
; 
32'd133770: dataIn1 = 32'd206
; 
32'd133771: dataIn1 = 32'd401
; 
32'd133772: dataIn1 = 32'd763
; 
32'd133773: dataIn1 = 32'd2290
; 
32'd133774: dataIn1 = 32'd2291
; 
32'd133775: dataIn1 = 32'd2524
; 
32'd133776: dataIn1 = 32'd2527
; 
32'd133777: dataIn1 = 32'd403
; 
32'd133778: dataIn1 = 32'd404
; 
32'd133779: dataIn1 = 32'd769
; 
32'd133780: dataIn1 = 32'd2290
; 
32'd133781: dataIn1 = 32'd2292
; 
32'd133782: dataIn1 = 32'd2293
; 
32'd133783: dataIn1 = 32'd2490
; 
32'd133784: dataIn1 = 32'd206
; 
32'd133785: dataIn1 = 32'd404
; 
32'd133786: dataIn1 = 32'd2290
; 
32'd133787: dataIn1 = 32'd2292
; 
32'd133788: dataIn1 = 32'd2293
; 
32'd133789: dataIn1 = 32'd3905
; 
32'd133790: dataIn1 = 32'd3922
; 
32'd133791: dataIn1 = 32'd5756
; 
32'd133792: dataIn1 = 32'd443
; 
32'd133793: dataIn1 = 32'd2294
; 
32'd133794: dataIn1 = 32'd3869
; 
32'd133795: dataIn1 = 32'd3870
; 
32'd133796: dataIn1 = 32'd3928
; 
32'd133797: dataIn1 = 32'd3929
; 
32'd133798: dataIn1 = 32'd3933
; 
32'd133799: dataIn1 = 32'd443
; 
32'd133800: dataIn1 = 32'd2295
; 
32'd133801: dataIn1 = 32'd3421
; 
32'd133802: dataIn1 = 32'd3449
; 
32'd133803: dataIn1 = 32'd3868
; 
32'd133804: dataIn1 = 32'd3870
; 
32'd133805: dataIn1 = 32'd5304
; 
32'd133806: dataIn1 = 32'd2296
; 
32'd133807: dataIn1 = 32'd3872
; 
32'd133808: dataIn1 = 32'd3873
; 
32'd133809: dataIn1 = 32'd3877
; 
32'd133810: dataIn1 = 32'd3879
; 
32'd133811: dataIn1 = 32'd3881
; 
32'd133812: dataIn1 = 32'd3882
; 
32'd133813: dataIn1 = 32'd5649
; 
32'd133814: dataIn1 = 32'd2297
; 
32'd133815: dataIn1 = 32'd5652
; 
32'd133816: dataIn1 = 32'd5653
; 
32'd133817: dataIn1 = 32'd5659
; 
32'd133818: dataIn1 = 32'd5664
; 
32'd133819: dataIn1 = 32'd5668
; 
32'd133820: dataIn1 = 32'd5670
; 
32'd133821: dataIn1 = 32'd2298
; 
32'd133822: dataIn1 = 32'd5654
; 
32'd133823: dataIn1 = 32'd5655
; 
32'd133824: dataIn1 = 32'd5660
; 
32'd133825: dataIn1 = 32'd5661
; 
32'd133826: dataIn1 = 32'd5684
; 
32'd133827: dataIn1 = 32'd5685
; 
32'd133828: dataIn1 = 32'd2299
; 
32'd133829: dataIn1 = 32'd3880
; 
32'd133830: dataIn1 = 32'd3882
; 
32'd133831: dataIn1 = 32'd3886
; 
32'd133832: dataIn1 = 32'd5780
; 
32'd133833: dataIn1 = 32'd5781
; 
32'd133834: dataIn1 = 32'd5788
; 
32'd133835: dataIn1 = 32'd2300
; 
32'd133836: dataIn1 = 32'd3880
; 
32'd133837: dataIn1 = 32'd3881
; 
32'd133838: dataIn1 = 32'd3883
; 
32'd133839: dataIn1 = 32'd3885
; 
32'd133840: dataIn1 = 32'd4827
; 
32'd133841: dataIn1 = 32'd4828
; 
32'd133842: dataIn1 = 32'd5943
; 
32'd133843: dataIn1 = 32'd2301
; 
32'd133844: dataIn1 = 32'd3888
; 
32'd133845: dataIn1 = 32'd3892
; 
32'd133846: dataIn1 = 32'd5675
; 
32'd133847: dataIn1 = 32'd5676
; 
32'd133848: dataIn1 = 32'd5799
; 
32'd133849: dataIn1 = 32'd5800
; 
32'd133850: dataIn1 = 32'd2302
; 
32'd133851: dataIn1 = 32'd3898
; 
32'd133852: dataIn1 = 32'd5318
; 
32'd133853: dataIn1 = 32'd5680
; 
32'd133854: dataIn1 = 32'd5681
; 
32'd133855: dataIn1 = 32'd5691
; 
32'd133856: dataIn1 = 32'd5950
; 
32'd133857: dataIn1 = 32'd2303
; 
32'd133858: dataIn1 = 32'd5696
; 
32'd133859: dataIn1 = 32'd5697
; 
32'd133860: dataIn1 = 32'd5705
; 
32'd133861: dataIn1 = 32'd5708
; 
32'd133862: dataIn1 = 32'd5712
; 
32'd133863: dataIn1 = 32'd5713
; 
32'd133864: dataIn1 = 32'd2304
; 
32'd133865: dataIn1 = 32'd3900
; 
32'd133866: dataIn1 = 32'd3902
; 
32'd133867: dataIn1 = 32'd3904
; 
32'd133868: dataIn1 = 32'd3907
; 
32'd133869: dataIn1 = 32'd3914
; 
32'd133870: dataIn1 = 32'd3916
; 
32'd133871: dataIn1 = 32'd5694
; 
32'd133872: dataIn1 = 32'd5728
; 
32'd133873: dataIn1 = 32'd2305
; 
32'd133874: dataIn1 = 32'd5698
; 
32'd133875: dataIn1 = 32'd5699
; 
32'd133876: dataIn1 = 32'd5700
; 
32'd133877: dataIn1 = 32'd5706
; 
32'd133878: dataIn1 = 32'd5750
; 
32'd133879: dataIn1 = 32'd5751
; 
32'd133880: dataIn1 = 32'd2306
; 
32'd133881: dataIn1 = 32'd3913
; 
32'd133882: dataIn1 = 32'd4881
; 
32'd133883: dataIn1 = 32'd5714
; 
32'd133884: dataIn1 = 32'd5715
; 
32'd133885: dataIn1 = 32'd5723
; 
32'd133886: dataIn1 = 32'd6064
; 
32'd133887: dataIn1 = 32'd2307
; 
32'd133888: dataIn1 = 32'd5730
; 
32'd133889: dataIn1 = 32'd5731
; 
32'd133890: dataIn1 = 32'd5739
; 
32'd133891: dataIn1 = 32'd5744
; 
32'd133892: dataIn1 = 32'd6049
; 
32'd133893: dataIn1 = 32'd6050
; 
32'd133894: dataIn1 = 32'd2308
; 
32'd133895: dataIn1 = 32'd5732
; 
32'd133896: dataIn1 = 32'd5733
; 
32'd133897: dataIn1 = 32'd5734
; 
32'd133898: dataIn1 = 32'd5742
; 
32'd133899: dataIn1 = 32'd5810
; 
32'd133900: dataIn1 = 32'd5811
; 
32'd133901: dataIn1 = 32'd2309
; 
32'd133902: dataIn1 = 32'd3925
; 
32'd133903: dataIn1 = 32'd5748
; 
32'd133904: dataIn1 = 32'd5749
; 
32'd133905: dataIn1 = 32'd5755
; 
32'd133906: dataIn1 = 32'd5801
; 
32'd133907: dataIn1 = 32'd5802
; 
32'd133908: dataIn1 = 32'd443
; 
32'd133909: dataIn1 = 32'd2310
; 
32'd133910: dataIn1 = 32'd3927
; 
32'd133911: dataIn1 = 32'd3929
; 
32'd133912: dataIn1 = 32'd3931
; 
32'd133913: dataIn1 = 32'd5319
; 
32'd133914: dataIn1 = 32'd5320
; 
32'd133915: dataIn1 = 32'd2311
; 
32'd133916: dataIn1 = 32'd3927
; 
32'd133917: dataIn1 = 32'd3928
; 
32'd133918: dataIn1 = 32'd3930
; 
32'd133919: dataIn1 = 32'd3932
; 
32'd133920: dataIn1 = 32'd3956
; 
32'd133921: dataIn1 = 32'd3957
; 
32'd133922: dataIn1 = 32'd2312
; 
32'd133923: dataIn1 = 32'd5760
; 
32'd133924: dataIn1 = 32'd5761
; 
32'd133925: dataIn1 = 32'd5769
; 
32'd133926: dataIn1 = 32'd5774
; 
32'd133927: dataIn1 = 32'd5778
; 
32'd133928: dataIn1 = 32'd5779
; 
32'd133929: dataIn1 = 32'd2313
; 
32'd133930: dataIn1 = 32'd3934
; 
32'd133931: dataIn1 = 32'd3936
; 
32'd133932: dataIn1 = 32'd3938
; 
32'd133933: dataIn1 = 32'd3941
; 
32'd133934: dataIn1 = 32'd3948
; 
32'd133935: dataIn1 = 32'd3950
; 
32'd133936: dataIn1 = 32'd5758
; 
32'd133937: dataIn1 = 32'd5797
; 
32'd133938: dataIn1 = 32'd2314
; 
32'd133939: dataIn1 = 32'd5762
; 
32'd133940: dataIn1 = 32'd5763
; 
32'd133941: dataIn1 = 32'd5764
; 
32'd133942: dataIn1 = 32'd5772
; 
32'd133943: dataIn1 = 32'd5812
; 
32'd133944: dataIn1 = 32'd5813
; 
32'd133945: dataIn1 = 32'd2315
; 
32'd133946: dataIn1 = 32'd5782
; 
32'd133947: dataIn1 = 32'd5783
; 
32'd133948: dataIn1 = 32'd5789
; 
32'd133949: dataIn1 = 32'd5794
; 
32'd133950: dataIn1 = 32'd7024
; 
32'd133951: dataIn1 = 32'd7025
; 
32'd133952: dataIn1 = 32'd2316
; 
32'd133953: dataIn1 = 32'd5808
; 
32'd133954: dataIn1 = 32'd5809
; 
32'd133955: dataIn1 = 32'd5820
; 
32'd133956: dataIn1 = 32'd5825
; 
32'd133957: dataIn1 = 32'd7040
; 
32'd133958: dataIn1 = 32'd7041
; 
32'd133959: dataIn1 = 32'd2317
; 
32'd133960: dataIn1 = 32'd3957
; 
32'd133961: dataIn1 = 32'd3958
; 
32'd133962: dataIn1 = 32'd3960
; 
32'd133963: dataIn1 = 32'd3962
; 
32'd133964: dataIn1 = 32'd3996
; 
32'd133965: dataIn1 = 32'd3997
; 
32'd133966: dataIn1 = 32'd2318
; 
32'd133967: dataIn1 = 32'd3956
; 
32'd133968: dataIn1 = 32'd3958
; 
32'd133969: dataIn1 = 32'd3959
; 
32'd133970: dataIn1 = 32'd3961
; 
32'd133971: dataIn1 = 32'd5321
; 
32'd133972: dataIn1 = 32'd5322
; 
32'd133973: dataIn1 = 32'd2319
; 
32'd133974: dataIn1 = 32'd6863
; 
32'd133975: dataIn1 = 32'd6864
; 
32'd133976: dataIn1 = 32'd6886
; 
32'd133977: dataIn1 = 32'd6903
; 
32'd133978: dataIn1 = 32'd6919
; 
32'd133979: dataIn1 = 32'd6920
; 
32'd133980: dataIn1 = 32'd2320
; 
32'd133981: dataIn1 = 32'd3967
; 
32'd133982: dataIn1 = 32'd3977
; 
32'd133983: dataIn1 = 32'd3979
; 
32'd133984: dataIn1 = 32'd9270
; 
32'd133985: dataIn1 = 32'd9271
; 
32'd133986: dataIn1 = 32'd9319
; 
32'd133987: dataIn1 = 32'd2321
; 
32'd133988: dataIn1 = 32'd5834
; 
32'd133989: dataIn1 = 32'd6872
; 
32'd133990: dataIn1 = 32'd6873
; 
32'd133991: dataIn1 = 32'd6899
; 
32'd133992: dataIn1 = 32'd7015
; 
32'd133993: dataIn1 = 32'd7016
; 
32'd133994: dataIn1 = 32'd2322
; 
32'd133995: dataIn1 = 32'd6927
; 
32'd133996: dataIn1 = 32'd6928
; 
32'd133997: dataIn1 = 32'd6949
; 
32'd133998: dataIn1 = 32'd6988
; 
32'd133999: dataIn1 = 32'd8891
; 
32'd134000: dataIn1 = 32'd8892
; 
32'd134001: dataIn1 = 32'd15
; 
32'd134002: dataIn1 = 32'd2323
; 
32'd134003: dataIn1 = 32'd2737
; 
32'd134004: dataIn1 = 32'd3978
; 
32'd134005: dataIn1 = 32'd3979
; 
32'd134006: dataIn1 = 32'd3980
; 
32'd134007: dataIn1 = 32'd6742
; 
32'd134008: dataIn1 = 32'd15
; 
32'd134009: dataIn1 = 32'd2324
; 
32'd134010: dataIn1 = 32'd2741
; 
32'd134011: dataIn1 = 32'd3977
; 
32'd134012: dataIn1 = 32'd3978
; 
32'd134013: dataIn1 = 32'd5323
; 
32'd134014: dataIn1 = 32'd6691
; 
32'd134015: dataIn1 = 32'd2325
; 
32'd134016: dataIn1 = 32'd5271
; 
32'd134017: dataIn1 = 32'd5876
; 
32'd134018: dataIn1 = 32'd5877
; 
32'd134019: dataIn1 = 32'd5887
; 
32'd134020: dataIn1 = 32'd6598
; 
32'd134021: dataIn1 = 32'd7006
; 
32'd134022: dataIn1 = 32'd7048
; 
32'd134023: dataIn1 = 32'd9272
; 
32'd134024: dataIn1 = 32'd2326
; 
32'd134025: dataIn1 = 32'd3987
; 
32'd134026: dataIn1 = 32'd3988
; 
32'd134027: dataIn1 = 32'd3992
; 
32'd134028: dataIn1 = 32'd3994
; 
32'd134029: dataIn1 = 32'd5324
; 
32'd134030: dataIn1 = 32'd5325
; 
32'd134031: dataIn1 = 32'd2327
; 
32'd134032: dataIn1 = 32'd3986
; 
32'd134033: dataIn1 = 32'd3988
; 
32'd134034: dataIn1 = 32'd3990
; 
32'd134035: dataIn1 = 32'd3993
; 
32'd134036: dataIn1 = 32'd3995
; 
32'd134037: dataIn1 = 32'd3997
; 
32'd134038: dataIn1 = 32'd2328
; 
32'd134039: dataIn1 = 32'd3986
; 
32'd134040: dataIn1 = 32'd3987
; 
32'd134041: dataIn1 = 32'd3989
; 
32'd134042: dataIn1 = 32'd3991
; 
32'd134043: dataIn1 = 32'd3998
; 
32'd134044: dataIn1 = 32'd3999
; 
32'd134045: dataIn1 = 32'd2329
; 
32'd134046: dataIn1 = 32'd3999
; 
32'd134047: dataIn1 = 32'd4000
; 
32'd134048: dataIn1 = 32'd4001
; 
32'd134049: dataIn1 = 32'd4003
; 
32'd134050: dataIn1 = 32'd4004
; 
32'd134051: dataIn1 = 32'd4009
; 
32'd134052: dataIn1 = 32'd2330
; 
32'd134053: dataIn1 = 32'd4002
; 
32'd134054: dataIn1 = 32'd4004
; 
32'd134055: dataIn1 = 32'd4006
; 
32'd134056: dataIn1 = 32'd4008
; 
32'd134057: dataIn1 = 32'd4023
; 
32'd134058: dataIn1 = 32'd4025
; 
32'd134059: dataIn1 = 32'd2331
; 
32'd134060: dataIn1 = 32'd4002
; 
32'd134061: dataIn1 = 32'd4003
; 
32'd134062: dataIn1 = 32'd4005
; 
32'd134063: dataIn1 = 32'd4007
; 
32'd134064: dataIn1 = 32'd5326
; 
32'd134065: dataIn1 = 32'd5327
; 
32'd134066: dataIn1 = 32'd2332
; 
32'd134067: dataIn1 = 32'd4011
; 
32'd134068: dataIn1 = 32'd4012
; 
32'd134069: dataIn1 = 32'd4016
; 
32'd134070: dataIn1 = 32'd4018
; 
32'd134071: dataIn1 = 32'd4020
; 
32'd134072: dataIn1 = 32'd4021
; 
32'd134073: dataIn1 = 32'd2333
; 
32'd134074: dataIn1 = 32'd4010
; 
32'd134075: dataIn1 = 32'd4012
; 
32'd134076: dataIn1 = 32'd4014
; 
32'd134077: dataIn1 = 32'd4017
; 
32'd134078: dataIn1 = 32'd5328
; 
32'd134079: dataIn1 = 32'd5329
; 
32'd134080: dataIn1 = 32'd2334
; 
32'd134081: dataIn1 = 32'd4010
; 
32'd134082: dataIn1 = 32'd4011
; 
32'd134083: dataIn1 = 32'd4013
; 
32'd134084: dataIn1 = 32'd4015
; 
32'd134085: dataIn1 = 32'd4023
; 
32'd134086: dataIn1 = 32'd4024
; 
32'd134087: dataIn1 = 32'd2335
; 
32'd134088: dataIn1 = 32'd4019
; 
32'd134089: dataIn1 = 32'd4021
; 
32'd134090: dataIn1 = 32'd4022
; 
32'd134091: dataIn1 = 32'd4026
; 
32'd134092: dataIn1 = 32'd4027
; 
32'd134093: dataIn1 = 32'd4029
; 
32'd134094: dataIn1 = 32'd2336
; 
32'd134095: dataIn1 = 32'd4027
; 
32'd134096: dataIn1 = 32'd4028
; 
32'd134097: dataIn1 = 32'd4031
; 
32'd134098: dataIn1 = 32'd4033
; 
32'd134099: dataIn1 = 32'd5330
; 
32'd134100: dataIn1 = 32'd5331
; 
32'd134101: dataIn1 = 32'd2337
; 
32'd134102: dataIn1 = 32'd4026
; 
32'd134103: dataIn1 = 32'd4028
; 
32'd134104: dataIn1 = 32'd4030
; 
32'd134105: dataIn1 = 32'd4032
; 
32'd134106: dataIn1 = 32'd4043
; 
32'd134107: dataIn1 = 32'd4045
; 
32'd134108: dataIn1 = 32'd2338
; 
32'd134109: dataIn1 = 32'd4035
; 
32'd134110: dataIn1 = 32'd4036
; 
32'd134111: dataIn1 = 32'd4040
; 
32'd134112: dataIn1 = 32'd4042
; 
32'd134113: dataIn1 = 32'd4044
; 
32'd134114: dataIn1 = 32'd4045
; 
32'd134115: dataIn1 = 32'd2339
; 
32'd134116: dataIn1 = 32'd4034
; 
32'd134117: dataIn1 = 32'd4036
; 
32'd134118: dataIn1 = 32'd4038
; 
32'd134119: dataIn1 = 32'd4041
; 
32'd134120: dataIn1 = 32'd5332
; 
32'd134121: dataIn1 = 32'd5333
; 
32'd134122: dataIn1 = 32'd2340
; 
32'd134123: dataIn1 = 32'd4034
; 
32'd134124: dataIn1 = 32'd4035
; 
32'd134125: dataIn1 = 32'd4037
; 
32'd134126: dataIn1 = 32'd4039
; 
32'd134127: dataIn1 = 32'd4046
; 
32'd134128: dataIn1 = 32'd4047
; 
32'd134129: dataIn1 = 32'd2341
; 
32'd134130: dataIn1 = 32'd4046
; 
32'd134131: dataIn1 = 32'd4048
; 
32'd134132: dataIn1 = 32'd4049
; 
32'd134133: dataIn1 = 32'd4050
; 
32'd134134: dataIn1 = 32'd4052
; 
32'd134135: dataIn1 = 32'd4056
; 
32'd134136: dataIn1 = 32'd2342
; 
32'd134137: dataIn1 = 32'd4051
; 
32'd134138: dataIn1 = 32'd4052
; 
32'd134139: dataIn1 = 32'd4055
; 
32'd134140: dataIn1 = 32'd4057
; 
32'd134141: dataIn1 = 32'd4067
; 
32'd134142: dataIn1 = 32'd4068
; 
32'd134143: dataIn1 = 32'd2343
; 
32'd134144: dataIn1 = 32'd4050
; 
32'd134145: dataIn1 = 32'd4051
; 
32'd134146: dataIn1 = 32'd4053
; 
32'd134147: dataIn1 = 32'd4054
; 
32'd134148: dataIn1 = 32'd5334
; 
32'd134149: dataIn1 = 32'd5335
; 
32'd134150: dataIn1 = 32'd2344
; 
32'd134151: dataIn1 = 32'd4059
; 
32'd134152: dataIn1 = 32'd4060
; 
32'd134153: dataIn1 = 32'd4064
; 
32'd134154: dataIn1 = 32'd4066
; 
32'd134155: dataIn1 = 32'd4068
; 
32'd134156: dataIn1 = 32'd4069
; 
32'd134157: dataIn1 = 32'd2345
; 
32'd134158: dataIn1 = 32'd4058
; 
32'd134159: dataIn1 = 32'd4060
; 
32'd134160: dataIn1 = 32'd4062
; 
32'd134161: dataIn1 = 32'd4065
; 
32'd134162: dataIn1 = 32'd4070
; 
32'd134163: dataIn1 = 32'd4072
; 
32'd134164: dataIn1 = 32'd2346
; 
32'd134165: dataIn1 = 32'd4058
; 
32'd134166: dataIn1 = 32'd4059
; 
32'd134167: dataIn1 = 32'd4061
; 
32'd134168: dataIn1 = 32'd4063
; 
32'd134169: dataIn1 = 32'd5336
; 
32'd134170: dataIn1 = 32'd5337
; 
32'd134171: dataIn1 = 32'd2347
; 
32'd134172: dataIn1 = 32'd4070
; 
32'd134173: dataIn1 = 32'd4071
; 
32'd134174: dataIn1 = 32'd4073
; 
32'd134175: dataIn1 = 32'd4074
; 
32'd134176: dataIn1 = 32'd4075
; 
32'd134177: dataIn1 = 32'd4078
; 
32'd134178: dataIn1 = 32'd2348
; 
32'd134179: dataIn1 = 32'd4075
; 
32'd134180: dataIn1 = 32'd4076
; 
32'd134181: dataIn1 = 32'd4079
; 
32'd134182: dataIn1 = 32'd4081
; 
32'd134183: dataIn1 = 32'd4092
; 
32'd134184: dataIn1 = 32'd4093
; 
32'd134185: dataIn1 = 32'd2349
; 
32'd134186: dataIn1 = 32'd4074
; 
32'd134187: dataIn1 = 32'd4076
; 
32'd134188: dataIn1 = 32'd4077
; 
32'd134189: dataIn1 = 32'd4080
; 
32'd134190: dataIn1 = 32'd5338
; 
32'd134191: dataIn1 = 32'd5339
; 
32'd134192: dataIn1 = 32'd2350
; 
32'd134193: dataIn1 = 32'd4083
; 
32'd134194: dataIn1 = 32'd4084
; 
32'd134195: dataIn1 = 32'd4088
; 
32'd134196: dataIn1 = 32'd4090
; 
32'd134197: dataIn1 = 32'd5340
; 
32'd134198: dataIn1 = 32'd5341
; 
32'd134199: dataIn1 = 32'd2351
; 
32'd134200: dataIn1 = 32'd4082
; 
32'd134201: dataIn1 = 32'd4084
; 
32'd134202: dataIn1 = 32'd4086
; 
32'd134203: dataIn1 = 32'd4089
; 
32'd134204: dataIn1 = 32'd4091
; 
32'd134205: dataIn1 = 32'd4093
; 
32'd134206: dataIn1 = 32'd2352
; 
32'd134207: dataIn1 = 32'd4082
; 
32'd134208: dataIn1 = 32'd4083
; 
32'd134209: dataIn1 = 32'd4085
; 
32'd134210: dataIn1 = 32'd4087
; 
32'd134211: dataIn1 = 32'd4094
; 
32'd134212: dataIn1 = 32'd4095
; 
32'd134213: dataIn1 = 32'd2353
; 
32'd134214: dataIn1 = 32'd4095
; 
32'd134215: dataIn1 = 32'd4096
; 
32'd134216: dataIn1 = 32'd4097
; 
32'd134217: dataIn1 = 32'd4099
; 
32'd134218: dataIn1 = 32'd4100
; 
32'd134219: dataIn1 = 32'd4105
; 
32'd134220: dataIn1 = 32'd2354
; 
32'd134221: dataIn1 = 32'd4098
; 
32'd134222: dataIn1 = 32'd4100
; 
32'd134223: dataIn1 = 32'd4102
; 
32'd134224: dataIn1 = 32'd4104
; 
32'd134225: dataIn1 = 32'd4119
; 
32'd134226: dataIn1 = 32'd4121
; 
32'd134227: dataIn1 = 32'd2355
; 
32'd134228: dataIn1 = 32'd4098
; 
32'd134229: dataIn1 = 32'd4099
; 
32'd134230: dataIn1 = 32'd4101
; 
32'd134231: dataIn1 = 32'd4103
; 
32'd134232: dataIn1 = 32'd5342
; 
32'd134233: dataIn1 = 32'd5343
; 
32'd134234: dataIn1 = 32'd2356
; 
32'd134235: dataIn1 = 32'd4107
; 
32'd134236: dataIn1 = 32'd4108
; 
32'd134237: dataIn1 = 32'd4112
; 
32'd134238: dataIn1 = 32'd4114
; 
32'd134239: dataIn1 = 32'd4116
; 
32'd134240: dataIn1 = 32'd4117
; 
32'd134241: dataIn1 = 32'd2357
; 
32'd134242: dataIn1 = 32'd4106
; 
32'd134243: dataIn1 = 32'd4108
; 
32'd134244: dataIn1 = 32'd4110
; 
32'd134245: dataIn1 = 32'd4113
; 
32'd134246: dataIn1 = 32'd5344
; 
32'd134247: dataIn1 = 32'd5345
; 
32'd134248: dataIn1 = 32'd2358
; 
32'd134249: dataIn1 = 32'd4106
; 
32'd134250: dataIn1 = 32'd4107
; 
32'd134251: dataIn1 = 32'd4109
; 
32'd134252: dataIn1 = 32'd4111
; 
32'd134253: dataIn1 = 32'd4119
; 
32'd134254: dataIn1 = 32'd4120
; 
32'd134255: dataIn1 = 32'd2359
; 
32'd134256: dataIn1 = 32'd4115
; 
32'd134257: dataIn1 = 32'd4117
; 
32'd134258: dataIn1 = 32'd4118
; 
32'd134259: dataIn1 = 32'd4122
; 
32'd134260: dataIn1 = 32'd4123
; 
32'd134261: dataIn1 = 32'd4125
; 
32'd134262: dataIn1 = 32'd2360
; 
32'd134263: dataIn1 = 32'd4123
; 
32'd134264: dataIn1 = 32'd4124
; 
32'd134265: dataIn1 = 32'd4127
; 
32'd134266: dataIn1 = 32'd4129
; 
32'd134267: dataIn1 = 32'd5346
; 
32'd134268: dataIn1 = 32'd5347
; 
32'd134269: dataIn1 = 32'd2361
; 
32'd134270: dataIn1 = 32'd4122
; 
32'd134271: dataIn1 = 32'd4124
; 
32'd134272: dataIn1 = 32'd4126
; 
32'd134273: dataIn1 = 32'd4128
; 
32'd134274: dataIn1 = 32'd4139
; 
32'd134275: dataIn1 = 32'd4141
; 
32'd134276: dataIn1 = 32'd2362
; 
32'd134277: dataIn1 = 32'd4131
; 
32'd134278: dataIn1 = 32'd4132
; 
32'd134279: dataIn1 = 32'd4136
; 
32'd134280: dataIn1 = 32'd4138
; 
32'd134281: dataIn1 = 32'd4140
; 
32'd134282: dataIn1 = 32'd4141
; 
32'd134283: dataIn1 = 32'd2363
; 
32'd134284: dataIn1 = 32'd4130
; 
32'd134285: dataIn1 = 32'd4132
; 
32'd134286: dataIn1 = 32'd4134
; 
32'd134287: dataIn1 = 32'd4137
; 
32'd134288: dataIn1 = 32'd5348
; 
32'd134289: dataIn1 = 32'd5349
; 
32'd134290: dataIn1 = 32'd2364
; 
32'd134291: dataIn1 = 32'd4130
; 
32'd134292: dataIn1 = 32'd4131
; 
32'd134293: dataIn1 = 32'd4133
; 
32'd134294: dataIn1 = 32'd4135
; 
32'd134295: dataIn1 = 32'd4142
; 
32'd134296: dataIn1 = 32'd4143
; 
32'd134297: dataIn1 = 32'd2365
; 
32'd134298: dataIn1 = 32'd4142
; 
32'd134299: dataIn1 = 32'd4144
; 
32'd134300: dataIn1 = 32'd4145
; 
32'd134301: dataIn1 = 32'd4146
; 
32'd134302: dataIn1 = 32'd4148
; 
32'd134303: dataIn1 = 32'd4152
; 
32'd134304: dataIn1 = 32'd2366
; 
32'd134305: dataIn1 = 32'd4147
; 
32'd134306: dataIn1 = 32'd4148
; 
32'd134307: dataIn1 = 32'd4151
; 
32'd134308: dataIn1 = 32'd4153
; 
32'd134309: dataIn1 = 32'd4163
; 
32'd134310: dataIn1 = 32'd4164
; 
32'd134311: dataIn1 = 32'd2367
; 
32'd134312: dataIn1 = 32'd4146
; 
32'd134313: dataIn1 = 32'd4147
; 
32'd134314: dataIn1 = 32'd4149
; 
32'd134315: dataIn1 = 32'd4150
; 
32'd134316: dataIn1 = 32'd5350
; 
32'd134317: dataIn1 = 32'd5351
; 
32'd134318: dataIn1 = 32'd2368
; 
32'd134319: dataIn1 = 32'd4155
; 
32'd134320: dataIn1 = 32'd4156
; 
32'd134321: dataIn1 = 32'd4160
; 
32'd134322: dataIn1 = 32'd4162
; 
32'd134323: dataIn1 = 32'd4164
; 
32'd134324: dataIn1 = 32'd4165
; 
32'd134325: dataIn1 = 32'd2369
; 
32'd134326: dataIn1 = 32'd4154
; 
32'd134327: dataIn1 = 32'd4156
; 
32'd134328: dataIn1 = 32'd4158
; 
32'd134329: dataIn1 = 32'd4161
; 
32'd134330: dataIn1 = 32'd4166
; 
32'd134331: dataIn1 = 32'd4168
; 
32'd134332: dataIn1 = 32'd2370
; 
32'd134333: dataIn1 = 32'd4154
; 
32'd134334: dataIn1 = 32'd4155
; 
32'd134335: dataIn1 = 32'd4157
; 
32'd134336: dataIn1 = 32'd4159
; 
32'd134337: dataIn1 = 32'd5352
; 
32'd134338: dataIn1 = 32'd5353
; 
32'd134339: dataIn1 = 32'd2371
; 
32'd134340: dataIn1 = 32'd4166
; 
32'd134341: dataIn1 = 32'd4167
; 
32'd134342: dataIn1 = 32'd4169
; 
32'd134343: dataIn1 = 32'd4170
; 
32'd134344: dataIn1 = 32'd4171
; 
32'd134345: dataIn1 = 32'd4174
; 
32'd134346: dataIn1 = 32'd2372
; 
32'd134347: dataIn1 = 32'd4171
; 
32'd134348: dataIn1 = 32'd4172
; 
32'd134349: dataIn1 = 32'd4175
; 
32'd134350: dataIn1 = 32'd4177
; 
32'd134351: dataIn1 = 32'd4188
; 
32'd134352: dataIn1 = 32'd4189
; 
32'd134353: dataIn1 = 32'd2373
; 
32'd134354: dataIn1 = 32'd4170
; 
32'd134355: dataIn1 = 32'd4172
; 
32'd134356: dataIn1 = 32'd4173
; 
32'd134357: dataIn1 = 32'd4176
; 
32'd134358: dataIn1 = 32'd5354
; 
32'd134359: dataIn1 = 32'd5355
; 
32'd134360: dataIn1 = 32'd2374
; 
32'd134361: dataIn1 = 32'd4179
; 
32'd134362: dataIn1 = 32'd4180
; 
32'd134363: dataIn1 = 32'd4184
; 
32'd134364: dataIn1 = 32'd4186
; 
32'd134365: dataIn1 = 32'd5356
; 
32'd134366: dataIn1 = 32'd5357
; 
32'd134367: dataIn1 = 32'd2375
; 
32'd134368: dataIn1 = 32'd4178
; 
32'd134369: dataIn1 = 32'd4180
; 
32'd134370: dataIn1 = 32'd4182
; 
32'd134371: dataIn1 = 32'd4185
; 
32'd134372: dataIn1 = 32'd4187
; 
32'd134373: dataIn1 = 32'd4189
; 
32'd134374: dataIn1 = 32'd2376
; 
32'd134375: dataIn1 = 32'd4178
; 
32'd134376: dataIn1 = 32'd4179
; 
32'd134377: dataIn1 = 32'd4181
; 
32'd134378: dataIn1 = 32'd4183
; 
32'd134379: dataIn1 = 32'd4190
; 
32'd134380: dataIn1 = 32'd4191
; 
32'd134381: dataIn1 = 32'd2377
; 
32'd134382: dataIn1 = 32'd4191
; 
32'd134383: dataIn1 = 32'd4192
; 
32'd134384: dataIn1 = 32'd4193
; 
32'd134385: dataIn1 = 32'd4195
; 
32'd134386: dataIn1 = 32'd4196
; 
32'd134387: dataIn1 = 32'd4201
; 
32'd134388: dataIn1 = 32'd2378
; 
32'd134389: dataIn1 = 32'd4194
; 
32'd134390: dataIn1 = 32'd4196
; 
32'd134391: dataIn1 = 32'd4198
; 
32'd134392: dataIn1 = 32'd4200
; 
32'd134393: dataIn1 = 32'd4215
; 
32'd134394: dataIn1 = 32'd4217
; 
32'd134395: dataIn1 = 32'd2379
; 
32'd134396: dataIn1 = 32'd4194
; 
32'd134397: dataIn1 = 32'd4195
; 
32'd134398: dataIn1 = 32'd4197
; 
32'd134399: dataIn1 = 32'd4199
; 
32'd134400: dataIn1 = 32'd5358
; 
32'd134401: dataIn1 = 32'd5359
; 
32'd134402: dataIn1 = 32'd2380
; 
32'd134403: dataIn1 = 32'd4203
; 
32'd134404: dataIn1 = 32'd4204
; 
32'd134405: dataIn1 = 32'd4208
; 
32'd134406: dataIn1 = 32'd4210
; 
32'd134407: dataIn1 = 32'd4212
; 
32'd134408: dataIn1 = 32'd4213
; 
32'd134409: dataIn1 = 32'd2381
; 
32'd134410: dataIn1 = 32'd4202
; 
32'd134411: dataIn1 = 32'd4204
; 
32'd134412: dataIn1 = 32'd4206
; 
32'd134413: dataIn1 = 32'd4209
; 
32'd134414: dataIn1 = 32'd5360
; 
32'd134415: dataIn1 = 32'd5361
; 
32'd134416: dataIn1 = 32'd2382
; 
32'd134417: dataIn1 = 32'd4202
; 
32'd134418: dataIn1 = 32'd4203
; 
32'd134419: dataIn1 = 32'd4205
; 
32'd134420: dataIn1 = 32'd4207
; 
32'd134421: dataIn1 = 32'd4215
; 
32'd134422: dataIn1 = 32'd4216
; 
32'd134423: dataIn1 = 32'd2383
; 
32'd134424: dataIn1 = 32'd4211
; 
32'd134425: dataIn1 = 32'd4213
; 
32'd134426: dataIn1 = 32'd4214
; 
32'd134427: dataIn1 = 32'd4218
; 
32'd134428: dataIn1 = 32'd4219
; 
32'd134429: dataIn1 = 32'd4221
; 
32'd134430: dataIn1 = 32'd2384
; 
32'd134431: dataIn1 = 32'd4219
; 
32'd134432: dataIn1 = 32'd4220
; 
32'd134433: dataIn1 = 32'd4223
; 
32'd134434: dataIn1 = 32'd4225
; 
32'd134435: dataIn1 = 32'd5362
; 
32'd134436: dataIn1 = 32'd5363
; 
32'd134437: dataIn1 = 32'd2385
; 
32'd134438: dataIn1 = 32'd4218
; 
32'd134439: dataIn1 = 32'd4220
; 
32'd134440: dataIn1 = 32'd4222
; 
32'd134441: dataIn1 = 32'd4224
; 
32'd134442: dataIn1 = 32'd4235
; 
32'd134443: dataIn1 = 32'd4237
; 
32'd134444: dataIn1 = 32'd2386
; 
32'd134445: dataIn1 = 32'd4227
; 
32'd134446: dataIn1 = 32'd4228
; 
32'd134447: dataIn1 = 32'd4232
; 
32'd134448: dataIn1 = 32'd4234
; 
32'd134449: dataIn1 = 32'd4236
; 
32'd134450: dataIn1 = 32'd4237
; 
32'd134451: dataIn1 = 32'd2387
; 
32'd134452: dataIn1 = 32'd4226
; 
32'd134453: dataIn1 = 32'd4228
; 
32'd134454: dataIn1 = 32'd4230
; 
32'd134455: dataIn1 = 32'd4233
; 
32'd134456: dataIn1 = 32'd5364
; 
32'd134457: dataIn1 = 32'd5365
; 
32'd134458: dataIn1 = 32'd2388
; 
32'd134459: dataIn1 = 32'd4226
; 
32'd134460: dataIn1 = 32'd4227
; 
32'd134461: dataIn1 = 32'd4229
; 
32'd134462: dataIn1 = 32'd4231
; 
32'd134463: dataIn1 = 32'd4238
; 
32'd134464: dataIn1 = 32'd4239
; 
32'd134465: dataIn1 = 32'd2389
; 
32'd134466: dataIn1 = 32'd4238
; 
32'd134467: dataIn1 = 32'd4240
; 
32'd134468: dataIn1 = 32'd4241
; 
32'd134469: dataIn1 = 32'd4242
; 
32'd134470: dataIn1 = 32'd4244
; 
32'd134471: dataIn1 = 32'd4248
; 
32'd134472: dataIn1 = 32'd2390
; 
32'd134473: dataIn1 = 32'd4243
; 
32'd134474: dataIn1 = 32'd4244
; 
32'd134475: dataIn1 = 32'd4247
; 
32'd134476: dataIn1 = 32'd4249
; 
32'd134477: dataIn1 = 32'd4259
; 
32'd134478: dataIn1 = 32'd4260
; 
32'd134479: dataIn1 = 32'd2391
; 
32'd134480: dataIn1 = 32'd4242
; 
32'd134481: dataIn1 = 32'd4243
; 
32'd134482: dataIn1 = 32'd4245
; 
32'd134483: dataIn1 = 32'd4246
; 
32'd134484: dataIn1 = 32'd5366
; 
32'd134485: dataIn1 = 32'd5367
; 
32'd134486: dataIn1 = 32'd2392
; 
32'd134487: dataIn1 = 32'd4251
; 
32'd134488: dataIn1 = 32'd4252
; 
32'd134489: dataIn1 = 32'd4256
; 
32'd134490: dataIn1 = 32'd4258
; 
32'd134491: dataIn1 = 32'd4260
; 
32'd134492: dataIn1 = 32'd4261
; 
32'd134493: dataIn1 = 32'd2393
; 
32'd134494: dataIn1 = 32'd4250
; 
32'd134495: dataIn1 = 32'd4252
; 
32'd134496: dataIn1 = 32'd4254
; 
32'd134497: dataIn1 = 32'd4257
; 
32'd134498: dataIn1 = 32'd4262
; 
32'd134499: dataIn1 = 32'd4264
; 
32'd134500: dataIn1 = 32'd2394
; 
32'd134501: dataIn1 = 32'd4250
; 
32'd134502: dataIn1 = 32'd4251
; 
32'd134503: dataIn1 = 32'd4253
; 
32'd134504: dataIn1 = 32'd4255
; 
32'd134505: dataIn1 = 32'd5368
; 
32'd134506: dataIn1 = 32'd5369
; 
32'd134507: dataIn1 = 32'd2395
; 
32'd134508: dataIn1 = 32'd4262
; 
32'd134509: dataIn1 = 32'd4263
; 
32'd134510: dataIn1 = 32'd4265
; 
32'd134511: dataIn1 = 32'd4266
; 
32'd134512: dataIn1 = 32'd4267
; 
32'd134513: dataIn1 = 32'd4270
; 
32'd134514: dataIn1 = 32'd2396
; 
32'd134515: dataIn1 = 32'd4267
; 
32'd134516: dataIn1 = 32'd4268
; 
32'd134517: dataIn1 = 32'd4271
; 
32'd134518: dataIn1 = 32'd4273
; 
32'd134519: dataIn1 = 32'd4284
; 
32'd134520: dataIn1 = 32'd4285
; 
32'd134521: dataIn1 = 32'd2397
; 
32'd134522: dataIn1 = 32'd4266
; 
32'd134523: dataIn1 = 32'd4268
; 
32'd134524: dataIn1 = 32'd4269
; 
32'd134525: dataIn1 = 32'd4272
; 
32'd134526: dataIn1 = 32'd5370
; 
32'd134527: dataIn1 = 32'd5371
; 
32'd134528: dataIn1 = 32'd2398
; 
32'd134529: dataIn1 = 32'd4275
; 
32'd134530: dataIn1 = 32'd4276
; 
32'd134531: dataIn1 = 32'd4280
; 
32'd134532: dataIn1 = 32'd4282
; 
32'd134533: dataIn1 = 32'd5372
; 
32'd134534: dataIn1 = 32'd5373
; 
32'd134535: dataIn1 = 32'd2399
; 
32'd134536: dataIn1 = 32'd4274
; 
32'd134537: dataIn1 = 32'd4276
; 
32'd134538: dataIn1 = 32'd4278
; 
32'd134539: dataIn1 = 32'd4281
; 
32'd134540: dataIn1 = 32'd4283
; 
32'd134541: dataIn1 = 32'd4285
; 
32'd134542: dataIn1 = 32'd2400
; 
32'd134543: dataIn1 = 32'd4274
; 
32'd134544: dataIn1 = 32'd4275
; 
32'd134545: dataIn1 = 32'd4277
; 
32'd134546: dataIn1 = 32'd4279
; 
32'd134547: dataIn1 = 32'd4286
; 
32'd134548: dataIn1 = 32'd4287
; 
32'd134549: dataIn1 = 32'd2401
; 
32'd134550: dataIn1 = 32'd4287
; 
32'd134551: dataIn1 = 32'd4288
; 
32'd134552: dataIn1 = 32'd4289
; 
32'd134553: dataIn1 = 32'd4291
; 
32'd134554: dataIn1 = 32'd4292
; 
32'd134555: dataIn1 = 32'd4297
; 
32'd134556: dataIn1 = 32'd2402
; 
32'd134557: dataIn1 = 32'd4290
; 
32'd134558: dataIn1 = 32'd4292
; 
32'd134559: dataIn1 = 32'd4294
; 
32'd134560: dataIn1 = 32'd4296
; 
32'd134561: dataIn1 = 32'd4311
; 
32'd134562: dataIn1 = 32'd4313
; 
32'd134563: dataIn1 = 32'd2403
; 
32'd134564: dataIn1 = 32'd4290
; 
32'd134565: dataIn1 = 32'd4291
; 
32'd134566: dataIn1 = 32'd4293
; 
32'd134567: dataIn1 = 32'd4295
; 
32'd134568: dataIn1 = 32'd5374
; 
32'd134569: dataIn1 = 32'd5375
; 
32'd134570: dataIn1 = 32'd2404
; 
32'd134571: dataIn1 = 32'd4299
; 
32'd134572: dataIn1 = 32'd4300
; 
32'd134573: dataIn1 = 32'd4304
; 
32'd134574: dataIn1 = 32'd4306
; 
32'd134575: dataIn1 = 32'd4308
; 
32'd134576: dataIn1 = 32'd4309
; 
32'd134577: dataIn1 = 32'd2405
; 
32'd134578: dataIn1 = 32'd4298
; 
32'd134579: dataIn1 = 32'd4300
; 
32'd134580: dataIn1 = 32'd4302
; 
32'd134581: dataIn1 = 32'd4305
; 
32'd134582: dataIn1 = 32'd5376
; 
32'd134583: dataIn1 = 32'd5377
; 
32'd134584: dataIn1 = 32'd2406
; 
32'd134585: dataIn1 = 32'd4298
; 
32'd134586: dataIn1 = 32'd4299
; 
32'd134587: dataIn1 = 32'd4301
; 
32'd134588: dataIn1 = 32'd4303
; 
32'd134589: dataIn1 = 32'd4311
; 
32'd134590: dataIn1 = 32'd4312
; 
32'd134591: dataIn1 = 32'd2407
; 
32'd134592: dataIn1 = 32'd4307
; 
32'd134593: dataIn1 = 32'd4309
; 
32'd134594: dataIn1 = 32'd4310
; 
32'd134595: dataIn1 = 32'd4314
; 
32'd134596: dataIn1 = 32'd4315
; 
32'd134597: dataIn1 = 32'd4317
; 
32'd134598: dataIn1 = 32'd2408
; 
32'd134599: dataIn1 = 32'd4315
; 
32'd134600: dataIn1 = 32'd4316
; 
32'd134601: dataIn1 = 32'd4319
; 
32'd134602: dataIn1 = 32'd4321
; 
32'd134603: dataIn1 = 32'd5378
; 
32'd134604: dataIn1 = 32'd5379
; 
32'd134605: dataIn1 = 32'd2409
; 
32'd134606: dataIn1 = 32'd4314
; 
32'd134607: dataIn1 = 32'd4316
; 
32'd134608: dataIn1 = 32'd4318
; 
32'd134609: dataIn1 = 32'd4320
; 
32'd134610: dataIn1 = 32'd4331
; 
32'd134611: dataIn1 = 32'd4333
; 
32'd134612: dataIn1 = 32'd2410
; 
32'd134613: dataIn1 = 32'd4323
; 
32'd134614: dataIn1 = 32'd4324
; 
32'd134615: dataIn1 = 32'd4328
; 
32'd134616: dataIn1 = 32'd4330
; 
32'd134617: dataIn1 = 32'd4332
; 
32'd134618: dataIn1 = 32'd4333
; 
32'd134619: dataIn1 = 32'd2411
; 
32'd134620: dataIn1 = 32'd4322
; 
32'd134621: dataIn1 = 32'd4324
; 
32'd134622: dataIn1 = 32'd4326
; 
32'd134623: dataIn1 = 32'd4329
; 
32'd134624: dataIn1 = 32'd5380
; 
32'd134625: dataIn1 = 32'd5381
; 
32'd134626: dataIn1 = 32'd2412
; 
32'd134627: dataIn1 = 32'd4322
; 
32'd134628: dataIn1 = 32'd4323
; 
32'd134629: dataIn1 = 32'd4325
; 
32'd134630: dataIn1 = 32'd4327
; 
32'd134631: dataIn1 = 32'd4334
; 
32'd134632: dataIn1 = 32'd4335
; 
32'd134633: dataIn1 = 32'd2413
; 
32'd134634: dataIn1 = 32'd4334
; 
32'd134635: dataIn1 = 32'd4336
; 
32'd134636: dataIn1 = 32'd4337
; 
32'd134637: dataIn1 = 32'd4338
; 
32'd134638: dataIn1 = 32'd4340
; 
32'd134639: dataIn1 = 32'd4344
; 
32'd134640: dataIn1 = 32'd2414
; 
32'd134641: dataIn1 = 32'd4339
; 
32'd134642: dataIn1 = 32'd4340
; 
32'd134643: dataIn1 = 32'd4343
; 
32'd134644: dataIn1 = 32'd4345
; 
32'd134645: dataIn1 = 32'd4355
; 
32'd134646: dataIn1 = 32'd4356
; 
32'd134647: dataIn1 = 32'd2415
; 
32'd134648: dataIn1 = 32'd4338
; 
32'd134649: dataIn1 = 32'd4339
; 
32'd134650: dataIn1 = 32'd4341
; 
32'd134651: dataIn1 = 32'd4342
; 
32'd134652: dataIn1 = 32'd5382
; 
32'd134653: dataIn1 = 32'd5383
; 
32'd134654: dataIn1 = 32'd2416
; 
32'd134655: dataIn1 = 32'd4347
; 
32'd134656: dataIn1 = 32'd4348
; 
32'd134657: dataIn1 = 32'd4352
; 
32'd134658: dataIn1 = 32'd4354
; 
32'd134659: dataIn1 = 32'd4356
; 
32'd134660: dataIn1 = 32'd4357
; 
32'd134661: dataIn1 = 32'd2417
; 
32'd134662: dataIn1 = 32'd4346
; 
32'd134663: dataIn1 = 32'd4348
; 
32'd134664: dataIn1 = 32'd4350
; 
32'd134665: dataIn1 = 32'd4353
; 
32'd134666: dataIn1 = 32'd4358
; 
32'd134667: dataIn1 = 32'd4360
; 
32'd134668: dataIn1 = 32'd2418
; 
32'd134669: dataIn1 = 32'd4346
; 
32'd134670: dataIn1 = 32'd4347
; 
32'd134671: dataIn1 = 32'd4349
; 
32'd134672: dataIn1 = 32'd4351
; 
32'd134673: dataIn1 = 32'd5384
; 
32'd134674: dataIn1 = 32'd5385
; 
32'd134675: dataIn1 = 32'd2419
; 
32'd134676: dataIn1 = 32'd4358
; 
32'd134677: dataIn1 = 32'd4359
; 
32'd134678: dataIn1 = 32'd4361
; 
32'd134679: dataIn1 = 32'd4362
; 
32'd134680: dataIn1 = 32'd4363
; 
32'd134681: dataIn1 = 32'd4366
; 
32'd134682: dataIn1 = 32'd2420
; 
32'd134683: dataIn1 = 32'd4363
; 
32'd134684: dataIn1 = 32'd4364
; 
32'd134685: dataIn1 = 32'd4367
; 
32'd134686: dataIn1 = 32'd4369
; 
32'd134687: dataIn1 = 32'd4380
; 
32'd134688: dataIn1 = 32'd4381
; 
32'd134689: dataIn1 = 32'd2421
; 
32'd134690: dataIn1 = 32'd4362
; 
32'd134691: dataIn1 = 32'd4364
; 
32'd134692: dataIn1 = 32'd4365
; 
32'd134693: dataIn1 = 32'd4368
; 
32'd134694: dataIn1 = 32'd5386
; 
32'd134695: dataIn1 = 32'd5387
; 
32'd134696: dataIn1 = 32'd2422
; 
32'd134697: dataIn1 = 32'd4371
; 
32'd134698: dataIn1 = 32'd4372
; 
32'd134699: dataIn1 = 32'd4376
; 
32'd134700: dataIn1 = 32'd4378
; 
32'd134701: dataIn1 = 32'd5388
; 
32'd134702: dataIn1 = 32'd5389
; 
32'd134703: dataIn1 = 32'd2423
; 
32'd134704: dataIn1 = 32'd4370
; 
32'd134705: dataIn1 = 32'd4372
; 
32'd134706: dataIn1 = 32'd4374
; 
32'd134707: dataIn1 = 32'd4377
; 
32'd134708: dataIn1 = 32'd4379
; 
32'd134709: dataIn1 = 32'd4381
; 
32'd134710: dataIn1 = 32'd2424
; 
32'd134711: dataIn1 = 32'd4370
; 
32'd134712: dataIn1 = 32'd4371
; 
32'd134713: dataIn1 = 32'd4373
; 
32'd134714: dataIn1 = 32'd4375
; 
32'd134715: dataIn1 = 32'd4382
; 
32'd134716: dataIn1 = 32'd4383
; 
32'd134717: dataIn1 = 32'd2425
; 
32'd134718: dataIn1 = 32'd4383
; 
32'd134719: dataIn1 = 32'd4384
; 
32'd134720: dataIn1 = 32'd4385
; 
32'd134721: dataIn1 = 32'd4387
; 
32'd134722: dataIn1 = 32'd4388
; 
32'd134723: dataIn1 = 32'd4393
; 
32'd134724: dataIn1 = 32'd2426
; 
32'd134725: dataIn1 = 32'd4386
; 
32'd134726: dataIn1 = 32'd4388
; 
32'd134727: dataIn1 = 32'd4390
; 
32'd134728: dataIn1 = 32'd4392
; 
32'd134729: dataIn1 = 32'd4407
; 
32'd134730: dataIn1 = 32'd4409
; 
32'd134731: dataIn1 = 32'd2427
; 
32'd134732: dataIn1 = 32'd4386
; 
32'd134733: dataIn1 = 32'd4387
; 
32'd134734: dataIn1 = 32'd4389
; 
32'd134735: dataIn1 = 32'd4391
; 
32'd134736: dataIn1 = 32'd5390
; 
32'd134737: dataIn1 = 32'd5391
; 
32'd134738: dataIn1 = 32'd2428
; 
32'd134739: dataIn1 = 32'd4395
; 
32'd134740: dataIn1 = 32'd4396
; 
32'd134741: dataIn1 = 32'd4400
; 
32'd134742: dataIn1 = 32'd4402
; 
32'd134743: dataIn1 = 32'd4404
; 
32'd134744: dataIn1 = 32'd4405
; 
32'd134745: dataIn1 = 32'd2429
; 
32'd134746: dataIn1 = 32'd4394
; 
32'd134747: dataIn1 = 32'd4396
; 
32'd134748: dataIn1 = 32'd4398
; 
32'd134749: dataIn1 = 32'd4401
; 
32'd134750: dataIn1 = 32'd5392
; 
32'd134751: dataIn1 = 32'd5393
; 
32'd134752: dataIn1 = 32'd2430
; 
32'd134753: dataIn1 = 32'd4394
; 
32'd134754: dataIn1 = 32'd4395
; 
32'd134755: dataIn1 = 32'd4397
; 
32'd134756: dataIn1 = 32'd4399
; 
32'd134757: dataIn1 = 32'd4407
; 
32'd134758: dataIn1 = 32'd4408
; 
32'd134759: dataIn1 = 32'd2431
; 
32'd134760: dataIn1 = 32'd4403
; 
32'd134761: dataIn1 = 32'd4405
; 
32'd134762: dataIn1 = 32'd4406
; 
32'd134763: dataIn1 = 32'd4410
; 
32'd134764: dataIn1 = 32'd4411
; 
32'd134765: dataIn1 = 32'd4413
; 
32'd134766: dataIn1 = 32'd2432
; 
32'd134767: dataIn1 = 32'd4411
; 
32'd134768: dataIn1 = 32'd4412
; 
32'd134769: dataIn1 = 32'd4415
; 
32'd134770: dataIn1 = 32'd4417
; 
32'd134771: dataIn1 = 32'd5394
; 
32'd134772: dataIn1 = 32'd5395
; 
32'd134773: dataIn1 = 32'd2433
; 
32'd134774: dataIn1 = 32'd4410
; 
32'd134775: dataIn1 = 32'd4412
; 
32'd134776: dataIn1 = 32'd4414
; 
32'd134777: dataIn1 = 32'd4416
; 
32'd134778: dataIn1 = 32'd4427
; 
32'd134779: dataIn1 = 32'd4429
; 
32'd134780: dataIn1 = 32'd2434
; 
32'd134781: dataIn1 = 32'd4419
; 
32'd134782: dataIn1 = 32'd4420
; 
32'd134783: dataIn1 = 32'd4424
; 
32'd134784: dataIn1 = 32'd4426
; 
32'd134785: dataIn1 = 32'd4428
; 
32'd134786: dataIn1 = 32'd4429
; 
32'd134787: dataIn1 = 32'd2435
; 
32'd134788: dataIn1 = 32'd4418
; 
32'd134789: dataIn1 = 32'd4420
; 
32'd134790: dataIn1 = 32'd4422
; 
32'd134791: dataIn1 = 32'd4425
; 
32'd134792: dataIn1 = 32'd5396
; 
32'd134793: dataIn1 = 32'd5397
; 
32'd134794: dataIn1 = 32'd2436
; 
32'd134795: dataIn1 = 32'd4418
; 
32'd134796: dataIn1 = 32'd4419
; 
32'd134797: dataIn1 = 32'd4421
; 
32'd134798: dataIn1 = 32'd4423
; 
32'd134799: dataIn1 = 32'd4430
; 
32'd134800: dataIn1 = 32'd4431
; 
32'd134801: dataIn1 = 32'd2437
; 
32'd134802: dataIn1 = 32'd4430
; 
32'd134803: dataIn1 = 32'd4432
; 
32'd134804: dataIn1 = 32'd4433
; 
32'd134805: dataIn1 = 32'd4434
; 
32'd134806: dataIn1 = 32'd4436
; 
32'd134807: dataIn1 = 32'd4440
; 
32'd134808: dataIn1 = 32'd2438
; 
32'd134809: dataIn1 = 32'd4435
; 
32'd134810: dataIn1 = 32'd4436
; 
32'd134811: dataIn1 = 32'd4439
; 
32'd134812: dataIn1 = 32'd4441
; 
32'd134813: dataIn1 = 32'd4451
; 
32'd134814: dataIn1 = 32'd4452
; 
32'd134815: dataIn1 = 32'd2439
; 
32'd134816: dataIn1 = 32'd4434
; 
32'd134817: dataIn1 = 32'd4435
; 
32'd134818: dataIn1 = 32'd4437
; 
32'd134819: dataIn1 = 32'd4438
; 
32'd134820: dataIn1 = 32'd5398
; 
32'd134821: dataIn1 = 32'd5399
; 
32'd134822: dataIn1 = 32'd2440
; 
32'd134823: dataIn1 = 32'd4443
; 
32'd134824: dataIn1 = 32'd4444
; 
32'd134825: dataIn1 = 32'd4448
; 
32'd134826: dataIn1 = 32'd4450
; 
32'd134827: dataIn1 = 32'd4452
; 
32'd134828: dataIn1 = 32'd4453
; 
32'd134829: dataIn1 = 32'd2441
; 
32'd134830: dataIn1 = 32'd4442
; 
32'd134831: dataIn1 = 32'd4444
; 
32'd134832: dataIn1 = 32'd4446
; 
32'd134833: dataIn1 = 32'd4449
; 
32'd134834: dataIn1 = 32'd4454
; 
32'd134835: dataIn1 = 32'd4456
; 
32'd134836: dataIn1 = 32'd2442
; 
32'd134837: dataIn1 = 32'd4442
; 
32'd134838: dataIn1 = 32'd4443
; 
32'd134839: dataIn1 = 32'd4445
; 
32'd134840: dataIn1 = 32'd4447
; 
32'd134841: dataIn1 = 32'd5400
; 
32'd134842: dataIn1 = 32'd5401
; 
32'd134843: dataIn1 = 32'd2443
; 
32'd134844: dataIn1 = 32'd4454
; 
32'd134845: dataIn1 = 32'd4455
; 
32'd134846: dataIn1 = 32'd4457
; 
32'd134847: dataIn1 = 32'd4458
; 
32'd134848: dataIn1 = 32'd4459
; 
32'd134849: dataIn1 = 32'd4462
; 
32'd134850: dataIn1 = 32'd2444
; 
32'd134851: dataIn1 = 32'd4459
; 
32'd134852: dataIn1 = 32'd4460
; 
32'd134853: dataIn1 = 32'd4463
; 
32'd134854: dataIn1 = 32'd4465
; 
32'd134855: dataIn1 = 32'd4476
; 
32'd134856: dataIn1 = 32'd4477
; 
32'd134857: dataIn1 = 32'd2445
; 
32'd134858: dataIn1 = 32'd4458
; 
32'd134859: dataIn1 = 32'd4460
; 
32'd134860: dataIn1 = 32'd4461
; 
32'd134861: dataIn1 = 32'd4464
; 
32'd134862: dataIn1 = 32'd5402
; 
32'd134863: dataIn1 = 32'd5403
; 
32'd134864: dataIn1 = 32'd2446
; 
32'd134865: dataIn1 = 32'd4467
; 
32'd134866: dataIn1 = 32'd4468
; 
32'd134867: dataIn1 = 32'd4472
; 
32'd134868: dataIn1 = 32'd4474
; 
32'd134869: dataIn1 = 32'd5404
; 
32'd134870: dataIn1 = 32'd5405
; 
32'd134871: dataIn1 = 32'd2447
; 
32'd134872: dataIn1 = 32'd4466
; 
32'd134873: dataIn1 = 32'd4468
; 
32'd134874: dataIn1 = 32'd4470
; 
32'd134875: dataIn1 = 32'd4473
; 
32'd134876: dataIn1 = 32'd4475
; 
32'd134877: dataIn1 = 32'd4477
; 
32'd134878: dataIn1 = 32'd2448
; 
32'd134879: dataIn1 = 32'd4466
; 
32'd134880: dataIn1 = 32'd4467
; 
32'd134881: dataIn1 = 32'd4469
; 
32'd134882: dataIn1 = 32'd4471
; 
32'd134883: dataIn1 = 32'd4478
; 
32'd134884: dataIn1 = 32'd4479
; 
32'd134885: dataIn1 = 32'd2449
; 
32'd134886: dataIn1 = 32'd4479
; 
32'd134887: dataIn1 = 32'd4480
; 
32'd134888: dataIn1 = 32'd4481
; 
32'd134889: dataIn1 = 32'd4483
; 
32'd134890: dataIn1 = 32'd4484
; 
32'd134891: dataIn1 = 32'd4489
; 
32'd134892: dataIn1 = 32'd2450
; 
32'd134893: dataIn1 = 32'd4482
; 
32'd134894: dataIn1 = 32'd4484
; 
32'd134895: dataIn1 = 32'd4486
; 
32'd134896: dataIn1 = 32'd4488
; 
32'd134897: dataIn1 = 32'd4503
; 
32'd134898: dataIn1 = 32'd4505
; 
32'd134899: dataIn1 = 32'd2451
; 
32'd134900: dataIn1 = 32'd4482
; 
32'd134901: dataIn1 = 32'd4483
; 
32'd134902: dataIn1 = 32'd4485
; 
32'd134903: dataIn1 = 32'd4487
; 
32'd134904: dataIn1 = 32'd5406
; 
32'd134905: dataIn1 = 32'd5407
; 
32'd134906: dataIn1 = 32'd2452
; 
32'd134907: dataIn1 = 32'd4491
; 
32'd134908: dataIn1 = 32'd4492
; 
32'd134909: dataIn1 = 32'd4496
; 
32'd134910: dataIn1 = 32'd4498
; 
32'd134911: dataIn1 = 32'd4500
; 
32'd134912: dataIn1 = 32'd4501
; 
32'd134913: dataIn1 = 32'd2453
; 
32'd134914: dataIn1 = 32'd4490
; 
32'd134915: dataIn1 = 32'd4492
; 
32'd134916: dataIn1 = 32'd4494
; 
32'd134917: dataIn1 = 32'd4497
; 
32'd134918: dataIn1 = 32'd5408
; 
32'd134919: dataIn1 = 32'd5409
; 
32'd134920: dataIn1 = 32'd2454
; 
32'd134921: dataIn1 = 32'd4490
; 
32'd134922: dataIn1 = 32'd4491
; 
32'd134923: dataIn1 = 32'd4493
; 
32'd134924: dataIn1 = 32'd4495
; 
32'd134925: dataIn1 = 32'd4503
; 
32'd134926: dataIn1 = 32'd4504
; 
32'd134927: dataIn1 = 32'd2455
; 
32'd134928: dataIn1 = 32'd4499
; 
32'd134929: dataIn1 = 32'd4501
; 
32'd134930: dataIn1 = 32'd4502
; 
32'd134931: dataIn1 = 32'd4506
; 
32'd134932: dataIn1 = 32'd4507
; 
32'd134933: dataIn1 = 32'd4509
; 
32'd134934: dataIn1 = 32'd2456
; 
32'd134935: dataIn1 = 32'd4507
; 
32'd134936: dataIn1 = 32'd4508
; 
32'd134937: dataIn1 = 32'd4511
; 
32'd134938: dataIn1 = 32'd4513
; 
32'd134939: dataIn1 = 32'd5410
; 
32'd134940: dataIn1 = 32'd5411
; 
32'd134941: dataIn1 = 32'd2457
; 
32'd134942: dataIn1 = 32'd4506
; 
32'd134943: dataIn1 = 32'd4508
; 
32'd134944: dataIn1 = 32'd4510
; 
32'd134945: dataIn1 = 32'd4512
; 
32'd134946: dataIn1 = 32'd4523
; 
32'd134947: dataIn1 = 32'd4525
; 
32'd134948: dataIn1 = 32'd2458
; 
32'd134949: dataIn1 = 32'd4515
; 
32'd134950: dataIn1 = 32'd4516
; 
32'd134951: dataIn1 = 32'd4520
; 
32'd134952: dataIn1 = 32'd4522
; 
32'd134953: dataIn1 = 32'd4524
; 
32'd134954: dataIn1 = 32'd4525
; 
32'd134955: dataIn1 = 32'd2459
; 
32'd134956: dataIn1 = 32'd4514
; 
32'd134957: dataIn1 = 32'd4516
; 
32'd134958: dataIn1 = 32'd4518
; 
32'd134959: dataIn1 = 32'd4521
; 
32'd134960: dataIn1 = 32'd5412
; 
32'd134961: dataIn1 = 32'd5413
; 
32'd134962: dataIn1 = 32'd2460
; 
32'd134963: dataIn1 = 32'd4514
; 
32'd134964: dataIn1 = 32'd4515
; 
32'd134965: dataIn1 = 32'd4517
; 
32'd134966: dataIn1 = 32'd4519
; 
32'd134967: dataIn1 = 32'd4526
; 
32'd134968: dataIn1 = 32'd4527
; 
32'd134969: dataIn1 = 32'd2461
; 
32'd134970: dataIn1 = 32'd4526
; 
32'd134971: dataIn1 = 32'd4528
; 
32'd134972: dataIn1 = 32'd4529
; 
32'd134973: dataIn1 = 32'd4530
; 
32'd134974: dataIn1 = 32'd4532
; 
32'd134975: dataIn1 = 32'd4536
; 
32'd134976: dataIn1 = 32'd2462
; 
32'd134977: dataIn1 = 32'd4531
; 
32'd134978: dataIn1 = 32'd4532
; 
32'd134979: dataIn1 = 32'd4535
; 
32'd134980: dataIn1 = 32'd4537
; 
32'd134981: dataIn1 = 32'd4547
; 
32'd134982: dataIn1 = 32'd4548
; 
32'd134983: dataIn1 = 32'd2463
; 
32'd134984: dataIn1 = 32'd4530
; 
32'd134985: dataIn1 = 32'd4531
; 
32'd134986: dataIn1 = 32'd4533
; 
32'd134987: dataIn1 = 32'd4534
; 
32'd134988: dataIn1 = 32'd5414
; 
32'd134989: dataIn1 = 32'd5415
; 
32'd134990: dataIn1 = 32'd2464
; 
32'd134991: dataIn1 = 32'd4539
; 
32'd134992: dataIn1 = 32'd4540
; 
32'd134993: dataIn1 = 32'd4544
; 
32'd134994: dataIn1 = 32'd4546
; 
32'd134995: dataIn1 = 32'd4548
; 
32'd134996: dataIn1 = 32'd4549
; 
32'd134997: dataIn1 = 32'd2465
; 
32'd134998: dataIn1 = 32'd4538
; 
32'd134999: dataIn1 = 32'd4540
; 
32'd135000: dataIn1 = 32'd4542
; 
32'd135001: dataIn1 = 32'd4545
; 
32'd135002: dataIn1 = 32'd4550
; 
32'd135003: dataIn1 = 32'd4552
; 
32'd135004: dataIn1 = 32'd2466
; 
32'd135005: dataIn1 = 32'd4538
; 
32'd135006: dataIn1 = 32'd4539
; 
32'd135007: dataIn1 = 32'd4541
; 
32'd135008: dataIn1 = 32'd4543
; 
32'd135009: dataIn1 = 32'd5416
; 
32'd135010: dataIn1 = 32'd2467
; 
32'd135011: dataIn1 = 32'd4550
; 
32'd135012: dataIn1 = 32'd4551
; 
32'd135013: dataIn1 = 32'd4553
; 
32'd135014: dataIn1 = 32'd4554
; 
32'd135015: dataIn1 = 32'd4555
; 
32'd135016: dataIn1 = 32'd4558
; 
32'd135017: dataIn1 = 32'd2468
; 
32'd135018: dataIn1 = 32'd4555
; 
32'd135019: dataIn1 = 32'd4556
; 
32'd135020: dataIn1 = 32'd4559
; 
32'd135021: dataIn1 = 32'd4561
; 
32'd135022: dataIn1 = 32'd4572
; 
32'd135023: dataIn1 = 32'd4573
; 
32'd135024: dataIn1 = 32'd2469
; 
32'd135025: dataIn1 = 32'd4554
; 
32'd135026: dataIn1 = 32'd4556
; 
32'd135027: dataIn1 = 32'd4557
; 
32'd135028: dataIn1 = 32'd4560
; 
32'd135029: dataIn1 = 32'd5419
; 
32'd135030: dataIn1 = 32'd2470
; 
32'd135031: dataIn1 = 32'd4563
; 
32'd135032: dataIn1 = 32'd4564
; 
32'd135033: dataIn1 = 32'd4568
; 
32'd135034: dataIn1 = 32'd4570
; 
32'd135035: dataIn1 = 32'd5420
; 
32'd135036: dataIn1 = 32'd2471
; 
32'd135037: dataIn1 = 32'd4562
; 
32'd135038: dataIn1 = 32'd4564
; 
32'd135039: dataIn1 = 32'd4566
; 
32'd135040: dataIn1 = 32'd4569
; 
32'd135041: dataIn1 = 32'd4571
; 
32'd135042: dataIn1 = 32'd4573
; 
32'd135043: dataIn1 = 32'd2472
; 
32'd135044: dataIn1 = 32'd4562
; 
32'd135045: dataIn1 = 32'd4563
; 
32'd135046: dataIn1 = 32'd4565
; 
32'd135047: dataIn1 = 32'd4567
; 
32'd135048: dataIn1 = 32'd4574
; 
32'd135049: dataIn1 = 32'd4575
; 
32'd135050: dataIn1 = 32'd2473
; 
32'd135051: dataIn1 = 32'd4575
; 
32'd135052: dataIn1 = 32'd4576
; 
32'd135053: dataIn1 = 32'd4577
; 
32'd135054: dataIn1 = 32'd4579
; 
32'd135055: dataIn1 = 32'd4580
; 
32'd135056: dataIn1 = 32'd4585
; 
32'd135057: dataIn1 = 32'd2474
; 
32'd135058: dataIn1 = 32'd4578
; 
32'd135059: dataIn1 = 32'd4580
; 
32'd135060: dataIn1 = 32'd4582
; 
32'd135061: dataIn1 = 32'd4584
; 
32'd135062: dataIn1 = 32'd4599
; 
32'd135063: dataIn1 = 32'd4601
; 
32'd135064: dataIn1 = 32'd2475
; 
32'd135065: dataIn1 = 32'd4578
; 
32'd135066: dataIn1 = 32'd4579
; 
32'd135067: dataIn1 = 32'd4581
; 
32'd135068: dataIn1 = 32'd4583
; 
32'd135069: dataIn1 = 32'd5422
; 
32'd135070: dataIn1 = 32'd2476
; 
32'd135071: dataIn1 = 32'd4587
; 
32'd135072: dataIn1 = 32'd4588
; 
32'd135073: dataIn1 = 32'd4592
; 
32'd135074: dataIn1 = 32'd4594
; 
32'd135075: dataIn1 = 32'd4596
; 
32'd135076: dataIn1 = 32'd4597
; 
32'd135077: dataIn1 = 32'd2477
; 
32'd135078: dataIn1 = 32'd4586
; 
32'd135079: dataIn1 = 32'd4588
; 
32'd135080: dataIn1 = 32'd4590
; 
32'd135081: dataIn1 = 32'd4593
; 
32'd135082: dataIn1 = 32'd5425
; 
32'd135083: dataIn1 = 32'd2478
; 
32'd135084: dataIn1 = 32'd4586
; 
32'd135085: dataIn1 = 32'd4587
; 
32'd135086: dataIn1 = 32'd4589
; 
32'd135087: dataIn1 = 32'd4591
; 
32'd135088: dataIn1 = 32'd4599
; 
32'd135089: dataIn1 = 32'd4600
; 
32'd135090: dataIn1 = 32'd2479
; 
32'd135091: dataIn1 = 32'd4595
; 
32'd135092: dataIn1 = 32'd4597
; 
32'd135093: dataIn1 = 32'd4598
; 
32'd135094: dataIn1 = 32'd5305
; 
32'd135095: dataIn1 = 32'd265
; 
32'd135096: dataIn1 = 32'd548
; 
32'd135097: dataIn1 = 32'd1260
; 
32'd135098: dataIn1 = 32'd2480
; 
32'd135099: dataIn1 = 32'd2481
; 
32'd135100: dataIn1 = 32'd2482
; 
32'd135101: dataIn1 = 32'd2755
; 
32'd135102: dataIn1 = 32'd265
; 
32'd135103: dataIn1 = 32'd542
; 
32'd135104: dataIn1 = 32'd1244
; 
32'd135105: dataIn1 = 32'd2480
; 
32'd135106: dataIn1 = 32'd2481
; 
32'd135107: dataIn1 = 32'd2482
; 
32'd135108: dataIn1 = 32'd2753
; 
32'd135109: dataIn1 = 32'd542
; 
32'd135110: dataIn1 = 32'd548
; 
32'd135111: dataIn1 = 32'd1262
; 
32'd135112: dataIn1 = 32'd2480
; 
32'd135113: dataIn1 = 32'd2481
; 
32'd135114: dataIn1 = 32'd2482
; 
32'd135115: dataIn1 = 32'd2756
; 
32'd135116: dataIn1 = 32'd584
; 
32'd135117: dataIn1 = 32'd586
; 
32'd135118: dataIn1 = 32'd1300
; 
32'd135119: dataIn1 = 32'd2483
; 
32'd135120: dataIn1 = 32'd2484
; 
32'd135121: dataIn1 = 32'd2485
; 
32'd135122: dataIn1 = 32'd2488
; 
32'd135123: dataIn1 = 32'd285
; 
32'd135124: dataIn1 = 32'd584
; 
32'd135125: dataIn1 = 32'd2483
; 
32'd135126: dataIn1 = 32'd2484
; 
32'd135127: dataIn1 = 32'd2485
; 
32'd135128: dataIn1 = 32'd2757
; 
32'd135129: dataIn1 = 32'd10983
; 
32'd135130: dataIn1 = 32'd10984
; 
32'd135131: dataIn1 = 32'd10985
; 
32'd135132: dataIn1 = 32'd285
; 
32'd135133: dataIn1 = 32'd586
; 
32'd135134: dataIn1 = 32'd2483
; 
32'd135135: dataIn1 = 32'd2484
; 
32'd135136: dataIn1 = 32'd2485
; 
32'd135137: dataIn1 = 32'd3421
; 
32'd135138: dataIn1 = 32'd156
; 
32'd135139: dataIn1 = 32'd586
; 
32'd135140: dataIn1 = 32'd2486
; 
32'd135141: dataIn1 = 32'd2487
; 
32'd135142: dataIn1 = 32'd2488
; 
32'd135143: dataIn1 = 32'd3420
; 
32'd135144: dataIn1 = 32'd156
; 
32'd135145: dataIn1 = 32'd585
; 
32'd135146: dataIn1 = 32'd2486
; 
32'd135147: dataIn1 = 32'd2487
; 
32'd135148: dataIn1 = 32'd2488
; 
32'd135149: dataIn1 = 32'd2521
; 
32'd135150: dataIn1 = 32'd2522
; 
32'd135151: dataIn1 = 32'd585
; 
32'd135152: dataIn1 = 32'd586
; 
32'd135153: dataIn1 = 32'd1300
; 
32'd135154: dataIn1 = 32'd2483
; 
32'd135155: dataIn1 = 32'd2486
; 
32'd135156: dataIn1 = 32'd2487
; 
32'd135157: dataIn1 = 32'd2488
; 
32'd135158: dataIn1 = 32'd396
; 
32'd135159: dataIn1 = 32'd400
; 
32'd135160: dataIn1 = 32'd761
; 
32'd135161: dataIn1 = 32'd2289
; 
32'd135162: dataIn1 = 32'd2489
; 
32'd135163: dataIn1 = 32'd3897
; 
32'd135164: dataIn1 = 32'd4602
; 
32'd135165: dataIn1 = 32'd404
; 
32'd135166: dataIn1 = 32'd405
; 
32'd135167: dataIn1 = 32'd769
; 
32'd135168: dataIn1 = 32'd2292
; 
32'd135169: dataIn1 = 32'd2490
; 
32'd135170: dataIn1 = 32'd3926
; 
32'd135171: dataIn1 = 32'd4603
; 
32'd135172: dataIn1 = 32'd407
; 
32'd135173: dataIn1 = 32'd777
; 
32'd135174: dataIn1 = 32'd1485
; 
32'd135175: dataIn1 = 32'd2491
; 
32'd135176: dataIn1 = 32'd2492
; 
32'd135177: dataIn1 = 32'd2493
; 
32'd135178: dataIn1 = 32'd2499
; 
32'd135179: dataIn1 = 32'd775
; 
32'd135180: dataIn1 = 32'd777
; 
32'd135181: dataIn1 = 32'd1481
; 
32'd135182: dataIn1 = 32'd2491
; 
32'd135183: dataIn1 = 32'd2492
; 
32'd135184: dataIn1 = 32'd2493
; 
32'd135185: dataIn1 = 32'd2496
; 
32'd135186: dataIn1 = 32'd407
; 
32'd135187: dataIn1 = 32'd775
; 
32'd135188: dataIn1 = 32'd2491
; 
32'd135189: dataIn1 = 32'd2492
; 
32'd135190: dataIn1 = 32'd2493
; 
32'd135191: dataIn1 = 32'd3423
; 
32'd135192: dataIn1 = 32'd408
; 
32'd135193: dataIn1 = 32'd776
; 
32'd135194: dataIn1 = 32'd1482
; 
32'd135195: dataIn1 = 32'd2494
; 
32'd135196: dataIn1 = 32'd2495
; 
32'd135197: dataIn1 = 32'd2496
; 
32'd135198: dataIn1 = 32'd2504
; 
32'd135199: dataIn1 = 32'd408
; 
32'd135200: dataIn1 = 32'd775
; 
32'd135201: dataIn1 = 32'd2494
; 
32'd135202: dataIn1 = 32'd2495
; 
32'd135203: dataIn1 = 32'd2496
; 
32'd135204: dataIn1 = 32'd3422
; 
32'd135205: dataIn1 = 32'd775
; 
32'd135206: dataIn1 = 32'd776
; 
32'd135207: dataIn1 = 32'd1481
; 
32'd135208: dataIn1 = 32'd2492
; 
32'd135209: dataIn1 = 32'd2494
; 
32'd135210: dataIn1 = 32'd2495
; 
32'd135211: dataIn1 = 32'd2496
; 
32'd135212: dataIn1 = 32'd407
; 
32'd135213: dataIn1 = 32'd783
; 
32'd135214: dataIn1 = 32'd976
; 
32'd135215: dataIn1 = 32'd2497
; 
32'd135216: dataIn1 = 32'd2498
; 
32'd135217: dataIn1 = 32'd2499
; 
32'd135218: dataIn1 = 32'd780
; 
32'd135219: dataIn1 = 32'd783
; 
32'd135220: dataIn1 = 32'd1490
; 
32'd135221: dataIn1 = 32'd2497
; 
32'd135222: dataIn1 = 32'd2498
; 
32'd135223: dataIn1 = 32'd2499
; 
32'd135224: dataIn1 = 32'd2758
; 
32'd135225: dataIn1 = 32'd407
; 
32'd135226: dataIn1 = 32'd780
; 
32'd135227: dataIn1 = 32'd1485
; 
32'd135228: dataIn1 = 32'd2491
; 
32'd135229: dataIn1 = 32'd2497
; 
32'd135230: dataIn1 = 32'd2498
; 
32'd135231: dataIn1 = 32'd2499
; 
32'd135232: dataIn1 = 32'd784
; 
32'd135233: dataIn1 = 32'd785
; 
32'd135234: dataIn1 = 32'd1491
; 
32'd135235: dataIn1 = 32'd2500
; 
32'd135236: dataIn1 = 32'd2501
; 
32'd135237: dataIn1 = 32'd2502
; 
32'd135238: dataIn1 = 32'd2505
; 
32'd135239: dataIn1 = 32'd409
; 
32'd135240: dataIn1 = 32'd785
; 
32'd135241: dataIn1 = 32'd1493
; 
32'd135242: dataIn1 = 32'd2500
; 
32'd135243: dataIn1 = 32'd2501
; 
32'd135244: dataIn1 = 32'd2502
; 
32'd135245: dataIn1 = 32'd2509
; 
32'd135246: dataIn1 = 32'd409
; 
32'd135247: dataIn1 = 32'd784
; 
32'd135248: dataIn1 = 32'd2500
; 
32'd135249: dataIn1 = 32'd2501
; 
32'd135250: dataIn1 = 32'd2502
; 
32'd135251: dataIn1 = 32'd3425
; 
32'd135252: dataIn1 = 32'd408
; 
32'd135253: dataIn1 = 32'd784
; 
32'd135254: dataIn1 = 32'd2503
; 
32'd135255: dataIn1 = 32'd2504
; 
32'd135256: dataIn1 = 32'd2505
; 
32'd135257: dataIn1 = 32'd3424
; 
32'd135258: dataIn1 = 32'd408
; 
32'd135259: dataIn1 = 32'd778
; 
32'd135260: dataIn1 = 32'd1482
; 
32'd135261: dataIn1 = 32'd2494
; 
32'd135262: dataIn1 = 32'd2503
; 
32'd135263: dataIn1 = 32'd2504
; 
32'd135264: dataIn1 = 32'd2505
; 
32'd135265: dataIn1 = 32'd778
; 
32'd135266: dataIn1 = 32'd784
; 
32'd135267: dataIn1 = 32'd1491
; 
32'd135268: dataIn1 = 32'd2500
; 
32'd135269: dataIn1 = 32'd2503
; 
32'd135270: dataIn1 = 32'd2504
; 
32'd135271: dataIn1 = 32'd2505
; 
32'd135272: dataIn1 = 32'd411
; 
32'd135273: dataIn1 = 32'd788
; 
32'd135274: dataIn1 = 32'd1496
; 
32'd135275: dataIn1 = 32'd2506
; 
32'd135276: dataIn1 = 32'd2507
; 
32'd135277: dataIn1 = 32'd2508
; 
32'd135278: dataIn1 = 32'd2519
; 
32'd135279: dataIn1 = 32'd786
; 
32'd135280: dataIn1 = 32'd788
; 
32'd135281: dataIn1 = 32'd1492
; 
32'd135282: dataIn1 = 32'd2506
; 
32'd135283: dataIn1 = 32'd2507
; 
32'd135284: dataIn1 = 32'd2508
; 
32'd135285: dataIn1 = 32'd2511
; 
32'd135286: dataIn1 = 32'd411
; 
32'd135287: dataIn1 = 32'd786
; 
32'd135288: dataIn1 = 32'd2506
; 
32'd135289: dataIn1 = 32'd2507
; 
32'd135290: dataIn1 = 32'd2508
; 
32'd135291: dataIn1 = 32'd3427
; 
32'd135292: dataIn1 = 32'd409
; 
32'd135293: dataIn1 = 32'd787
; 
32'd135294: dataIn1 = 32'd1493
; 
32'd135295: dataIn1 = 32'd2501
; 
32'd135296: dataIn1 = 32'd2509
; 
32'd135297: dataIn1 = 32'd2510
; 
32'd135298: dataIn1 = 32'd2511
; 
32'd135299: dataIn1 = 32'd409
; 
32'd135300: dataIn1 = 32'd786
; 
32'd135301: dataIn1 = 32'd2509
; 
32'd135302: dataIn1 = 32'd2510
; 
32'd135303: dataIn1 = 32'd2511
; 
32'd135304: dataIn1 = 32'd3426
; 
32'd135305: dataIn1 = 32'd786
; 
32'd135306: dataIn1 = 32'd787
; 
32'd135307: dataIn1 = 32'd1492
; 
32'd135308: dataIn1 = 32'd2507
; 
32'd135309: dataIn1 = 32'd2509
; 
32'd135310: dataIn1 = 32'd2510
; 
32'd135311: dataIn1 = 32'd2511
; 
32'd135312: dataIn1 = 32'd799
; 
32'd135313: dataIn1 = 32'd800
; 
32'd135314: dataIn1 = 32'd1506
; 
32'd135315: dataIn1 = 32'd2512
; 
32'd135316: dataIn1 = 32'd2513
; 
32'd135317: dataIn1 = 32'd2514
; 
32'd135318: dataIn1 = 32'd2759
; 
32'd135319: dataIn1 = 32'd413
; 
32'd135320: dataIn1 = 32'd800
; 
32'd135321: dataIn1 = 32'd2512
; 
32'd135322: dataIn1 = 32'd2513
; 
32'd135323: dataIn1 = 32'd2514
; 
32'd135324: dataIn1 = 32'd10251
; 
32'd135325: dataIn1 = 32'd10264
; 
32'd135326: dataIn1 = 32'd413
; 
32'd135327: dataIn1 = 32'd799
; 
32'd135328: dataIn1 = 32'd1510
; 
32'd135329: dataIn1 = 32'd2512
; 
32'd135330: dataIn1 = 32'd2513
; 
32'd135331: dataIn1 = 32'd2514
; 
32'd135332: dataIn1 = 32'd2516
; 
32'd135333: dataIn1 = 32'd804
; 
32'd135334: dataIn1 = 32'd805
; 
32'd135335: dataIn1 = 32'd1513
; 
32'd135336: dataIn1 = 32'd2515
; 
32'd135337: dataIn1 = 32'd2516
; 
32'd135338: dataIn1 = 32'd2517
; 
32'd135339: dataIn1 = 32'd2520
; 
32'd135340: dataIn1 = 32'd413
; 
32'd135341: dataIn1 = 32'd804
; 
32'd135342: dataIn1 = 32'd1510
; 
32'd135343: dataIn1 = 32'd2514
; 
32'd135344: dataIn1 = 32'd2515
; 
32'd135345: dataIn1 = 32'd2516
; 
32'd135346: dataIn1 = 32'd2517
; 
32'd135347: dataIn1 = 32'd413
; 
32'd135348: dataIn1 = 32'd805
; 
32'd135349: dataIn1 = 32'd2515
; 
32'd135350: dataIn1 = 32'd2516
; 
32'd135351: dataIn1 = 32'd2517
; 
32'd135352: dataIn1 = 32'd3429
; 
32'd135353: dataIn1 = 32'd411
; 
32'd135354: dataIn1 = 32'd805
; 
32'd135355: dataIn1 = 32'd2518
; 
32'd135356: dataIn1 = 32'd2519
; 
32'd135357: dataIn1 = 32'd2520
; 
32'd135358: dataIn1 = 32'd3428
; 
32'd135359: dataIn1 = 32'd411
; 
32'd135360: dataIn1 = 32'd790
; 
32'd135361: dataIn1 = 32'd1496
; 
32'd135362: dataIn1 = 32'd2506
; 
32'd135363: dataIn1 = 32'd2518
; 
32'd135364: dataIn1 = 32'd2519
; 
32'd135365: dataIn1 = 32'd2520
; 
32'd135366: dataIn1 = 32'd790
; 
32'd135367: dataIn1 = 32'd805
; 
32'd135368: dataIn1 = 32'd1513
; 
32'd135369: dataIn1 = 32'd2515
; 
32'd135370: dataIn1 = 32'd2518
; 
32'd135371: dataIn1 = 32'd2519
; 
32'd135372: dataIn1 = 32'd2520
; 
32'd135373: dataIn1 = 32'd156
; 
32'd135374: dataIn1 = 32'd806
; 
32'd135375: dataIn1 = 32'd2487
; 
32'd135376: dataIn1 = 32'd2521
; 
32'd135377: dataIn1 = 32'd2522
; 
32'd135378: dataIn1 = 32'd10252
; 
32'd135379: dataIn1 = 32'd10265
; 
32'd135380: dataIn1 = 32'd585
; 
32'd135381: dataIn1 = 32'd806
; 
32'd135382: dataIn1 = 32'd1518
; 
32'd135383: dataIn1 = 32'd2487
; 
32'd135384: dataIn1 = 32'd2521
; 
32'd135385: dataIn1 = 32'd2522
; 
32'd135386: dataIn1 = 32'd2760
; 
32'd135387: dataIn1 = 32'd973
; 
32'd135388: dataIn1 = 32'd974
; 
32'd135389: dataIn1 = 32'd2045
; 
32'd135390: dataIn1 = 32'd2523
; 
32'd135391: dataIn1 = 32'd2524
; 
32'd135392: dataIn1 = 32'd2525
; 
32'd135393: dataIn1 = 32'd2526
; 
32'd135394: dataIn1 = 32'd5724
; 
32'd135395: dataIn1 = 32'd401
; 
32'd135396: dataIn1 = 32'd974
; 
32'd135397: dataIn1 = 32'd2045
; 
32'd135398: dataIn1 = 32'd2291
; 
32'd135399: dataIn1 = 32'd2523
; 
32'd135400: dataIn1 = 32'd2524
; 
32'd135401: dataIn1 = 32'd2527
; 
32'd135402: dataIn1 = 32'd2523
; 
32'd135403: dataIn1 = 32'd2525
; 
32'd135404: dataIn1 = 32'd2526
; 
32'd135405: dataIn1 = 32'd5718
; 
32'd135406: dataIn1 = 32'd5720
; 
32'd135407: dataIn1 = 32'd5722
; 
32'd135408: dataIn1 = 32'd5724
; 
32'd135409: dataIn1 = 32'd129
; 
32'd135410: dataIn1 = 32'd973
; 
32'd135411: dataIn1 = 32'd2043
; 
32'd135412: dataIn1 = 32'd2523
; 
32'd135413: dataIn1 = 32'd2525
; 
32'd135414: dataIn1 = 32'd2526
; 
32'd135415: dataIn1 = 32'd2528
; 
32'd135416: dataIn1 = 32'd5722
; 
32'd135417: dataIn1 = 32'd206
; 
32'd135418: dataIn1 = 32'd974
; 
32'd135419: dataIn1 = 32'd2291
; 
32'd135420: dataIn1 = 32'd2524
; 
32'd135421: dataIn1 = 32'd2527
; 
32'd135422: dataIn1 = 32'd3906
; 
32'd135423: dataIn1 = 32'd3910
; 
32'd135424: dataIn1 = 32'd5716
; 
32'd135425: dataIn1 = 32'd5725
; 
32'd135426: dataIn1 = 32'd129
; 
32'd135427: dataIn1 = 32'd975
; 
32'd135428: dataIn1 = 32'd2043
; 
32'd135429: dataIn1 = 32'd2526
; 
32'd135430: dataIn1 = 32'd2528
; 
32'd135431: dataIn1 = 32'd2537
; 
32'd135432: dataIn1 = 32'd2539
; 
32'd135433: dataIn1 = 32'd5937
; 
32'd135434: dataIn1 = 32'd209
; 
32'd135435: dataIn1 = 32'd978
; 
32'd135436: dataIn1 = 32'd2046
; 
32'd135437: dataIn1 = 32'd2529
; 
32'd135438: dataIn1 = 32'd2530
; 
32'd135439: dataIn1 = 32'd2536
; 
32'd135440: dataIn1 = 32'd2538
; 
32'd135441: dataIn1 = 32'd5930
; 
32'd135442: dataIn1 = 32'd209
; 
32'd135443: dataIn1 = 32'd977
; 
32'd135444: dataIn1 = 32'd2046
; 
32'd135445: dataIn1 = 32'd2529
; 
32'd135446: dataIn1 = 32'd2530
; 
32'd135447: dataIn1 = 32'd2540
; 
32'd135448: dataIn1 = 32'd2542
; 
32'd135449: dataIn1 = 32'd4617
; 
32'd135450: dataIn1 = 32'd5920
; 
32'd135451: dataIn1 = 32'd2051
; 
32'd135452: dataIn1 = 32'd2531
; 
32'd135453: dataIn1 = 32'd4605
; 
32'd135454: dataIn1 = 32'd4606
; 
32'd135455: dataIn1 = 32'd4631
; 
32'd135456: dataIn1 = 32'd4632
; 
32'd135457: dataIn1 = 32'd4634
; 
32'd135458: dataIn1 = 32'd982
; 
32'd135459: dataIn1 = 32'd2051
; 
32'd135460: dataIn1 = 32'd2532
; 
32'd135461: dataIn1 = 32'd4604
; 
32'd135462: dataIn1 = 32'd4606
; 
32'd135463: dataIn1 = 32'd4618
; 
32'd135464: dataIn1 = 32'd4619
; 
32'd135465: dataIn1 = 32'd1039
; 
32'd135466: dataIn1 = 32'd2533
; 
32'd135467: dataIn1 = 32'd2534
; 
32'd135468: dataIn1 = 32'd4608
; 
32'd135469: dataIn1 = 32'd4609
; 
32'd135470: dataIn1 = 32'd4612
; 
32'd135471: dataIn1 = 32'd5306
; 
32'd135472: dataIn1 = 32'd202
; 
32'd135473: dataIn1 = 32'd969
; 
32'd135474: dataIn1 = 32'd1039
; 
32'd135475: dataIn1 = 32'd2039
; 
32'd135476: dataIn1 = 32'd2533
; 
32'd135477: dataIn1 = 32'd2534
; 
32'd135478: dataIn1 = 32'd5306
; 
32'd135479: dataIn1 = 32'd1039
; 
32'd135480: dataIn1 = 32'd2535
; 
32'd135481: dataIn1 = 32'd4607
; 
32'd135482: dataIn1 = 32'd4609
; 
32'd135483: dataIn1 = 32'd4610
; 
32'd135484: dataIn1 = 32'd4642
; 
32'd135485: dataIn1 = 32'd6698
; 
32'd135486: dataIn1 = 32'd978
; 
32'd135487: dataIn1 = 32'd1040
; 
32'd135488: dataIn1 = 32'd2044
; 
32'd135489: dataIn1 = 32'd2529
; 
32'd135490: dataIn1 = 32'd2536
; 
32'd135491: dataIn1 = 32'd2537
; 
32'd135492: dataIn1 = 32'd2538
; 
32'd135493: dataIn1 = 32'd5931
; 
32'd135494: dataIn1 = 32'd975
; 
32'd135495: dataIn1 = 32'd1040
; 
32'd135496: dataIn1 = 32'd2044
; 
32'd135497: dataIn1 = 32'd2528
; 
32'd135498: dataIn1 = 32'd2536
; 
32'd135499: dataIn1 = 32'd2537
; 
32'd135500: dataIn1 = 32'd2539
; 
32'd135501: dataIn1 = 32'd5935
; 
32'd135502: dataIn1 = 32'd2529
; 
32'd135503: dataIn1 = 32'd2536
; 
32'd135504: dataIn1 = 32'd2538
; 
32'd135505: dataIn1 = 32'd5927
; 
32'd135506: dataIn1 = 32'd5928
; 
32'd135507: dataIn1 = 32'd5930
; 
32'd135508: dataIn1 = 32'd5931
; 
32'd135509: dataIn1 = 32'd2528
; 
32'd135510: dataIn1 = 32'd2537
; 
32'd135511: dataIn1 = 32'd2539
; 
32'd135512: dataIn1 = 32'd5933
; 
32'd135513: dataIn1 = 32'd5934
; 
32'd135514: dataIn1 = 32'd5935
; 
32'd135515: dataIn1 = 32'd5937
; 
32'd135516: dataIn1 = 32'd977
; 
32'd135517: dataIn1 = 32'd2047
; 
32'd135518: dataIn1 = 32'd2530
; 
32'd135519: dataIn1 = 32'd2540
; 
32'd135520: dataIn1 = 32'd4614
; 
32'd135521: dataIn1 = 32'd4615
; 
32'd135522: dataIn1 = 32'd4617
; 
32'd135523: dataIn1 = 32'd982
; 
32'd135524: dataIn1 = 32'd2047
; 
32'd135525: dataIn1 = 32'd2541
; 
32'd135526: dataIn1 = 32'd4613
; 
32'd135527: dataIn1 = 32'd4615
; 
32'd135528: dataIn1 = 32'd4618
; 
32'd135529: dataIn1 = 32'd4620
; 
32'd135530: dataIn1 = 32'd2530
; 
32'd135531: dataIn1 = 32'd2542
; 
32'd135532: dataIn1 = 32'd4616
; 
32'd135533: dataIn1 = 32'd4617
; 
32'd135534: dataIn1 = 32'd5917
; 
32'd135535: dataIn1 = 32'd5919
; 
32'd135536: dataIn1 = 32'd5920
; 
32'd135537: dataIn1 = 32'd2543
; 
32'd135538: dataIn1 = 32'd4619
; 
32'd135539: dataIn1 = 32'd4620
; 
32'd135540: dataIn1 = 32'd4621
; 
32'd135541: dataIn1 = 32'd4622
; 
32'd135542: dataIn1 = 32'd5922
; 
32'd135543: dataIn1 = 32'd5923
; 
32'd135544: dataIn1 = 32'd2544
; 
32'd135545: dataIn1 = 32'd4623
; 
32'd135546: dataIn1 = 32'd4625
; 
32'd135547: dataIn1 = 32'd4627
; 
32'd135548: dataIn1 = 32'd5307
; 
32'd135549: dataIn1 = 32'd5428
; 
32'd135550: dataIn1 = 32'd5429
; 
32'd135551: dataIn1 = 32'd2545
; 
32'd135552: dataIn1 = 32'd4623
; 
32'd135553: dataIn1 = 32'd4624
; 
32'd135554: dataIn1 = 32'd4626
; 
32'd135555: dataIn1 = 32'd4628
; 
32'd135556: dataIn1 = 32'd4630
; 
32'd135557: dataIn1 = 32'd4631
; 
32'd135558: dataIn1 = 32'd2546
; 
32'd135559: dataIn1 = 32'd4630
; 
32'd135560: dataIn1 = 32'd4632
; 
32'd135561: dataIn1 = 32'd4633
; 
32'd135562: dataIn1 = 32'd4635
; 
32'd135563: dataIn1 = 32'd4683
; 
32'd135564: dataIn1 = 32'd6699
; 
32'd135565: dataIn1 = 32'd1069
; 
32'd135566: dataIn1 = 32'd2547
; 
32'd135567: dataIn1 = 32'd2548
; 
32'd135568: dataIn1 = 32'd4637
; 
32'd135569: dataIn1 = 32'd4638
; 
32'd135570: dataIn1 = 32'd4800
; 
32'd135571: dataIn1 = 32'd4801
; 
32'd135572: dataIn1 = 32'd1068
; 
32'd135573: dataIn1 = 32'd1069
; 
32'd135574: dataIn1 = 32'd2547
; 
32'd135575: dataIn1 = 32'd2548
; 
32'd135576: dataIn1 = 32'd3488
; 
32'd135577: dataIn1 = 32'd3492
; 
32'd135578: dataIn1 = 32'd4637
; 
32'd135579: dataIn1 = 32'd1068
; 
32'd135580: dataIn1 = 32'd2549
; 
32'd135581: dataIn1 = 32'd4636
; 
32'd135582: dataIn1 = 32'd4637
; 
32'd135583: dataIn1 = 32'd1070
; 
32'd135584: dataIn1 = 32'd1071
; 
32'd135585: dataIn1 = 32'd2550
; 
32'd135586: dataIn1 = 32'd2551
; 
32'd135587: dataIn1 = 32'd2552
; 
32'd135588: dataIn1 = 32'd3472
; 
32'd135589: dataIn1 = 32'd3476
; 
32'd135590: dataIn1 = 32'd4639
; 
32'd135591: dataIn1 = 32'd1071
; 
32'd135592: dataIn1 = 32'd2550
; 
32'd135593: dataIn1 = 32'd2551
; 
32'd135594: dataIn1 = 32'd4639
; 
32'd135595: dataIn1 = 32'd4641
; 
32'd135596: dataIn1 = 32'd4808
; 
32'd135597: dataIn1 = 32'd4810
; 
32'd135598: dataIn1 = 32'd1070
; 
32'd135599: dataIn1 = 32'd2550
; 
32'd135600: dataIn1 = 32'd2552
; 
32'd135601: dataIn1 = 32'd4639
; 
32'd135602: dataIn1 = 32'd4640
; 
32'd135603: dataIn1 = 32'd4795
; 
32'd135604: dataIn1 = 32'd4796
; 
32'd135605: dataIn1 = 32'd202
; 
32'd135606: dataIn1 = 32'd1039
; 
32'd135607: dataIn1 = 32'd1073
; 
32'd135608: dataIn1 = 32'd2553
; 
32'd135609: dataIn1 = 32'd2554
; 
32'd135610: dataIn1 = 32'd2556
; 
32'd135611: dataIn1 = 32'd3430
; 
32'd135612: dataIn1 = 32'd4642
; 
32'd135613: dataIn1 = 32'd5512
; 
32'd135614: dataIn1 = 32'd2553
; 
32'd135615: dataIn1 = 32'd2554
; 
32'd135616: dataIn1 = 32'd4642
; 
32'd135617: dataIn1 = 32'd4643
; 
32'd135618: dataIn1 = 32'd4838
; 
32'd135619: dataIn1 = 32'd5430
; 
32'd135620: dataIn1 = 32'd5512
; 
32'd135621: dataIn1 = 32'd5948
; 
32'd135622: dataIn1 = 32'd2555
; 
32'd135623: dataIn1 = 32'd2556
; 
32'd135624: dataIn1 = 32'd4645
; 
32'd135625: dataIn1 = 32'd4646
; 
32'd135626: dataIn1 = 32'd4832
; 
32'd135627: dataIn1 = 32'd4833
; 
32'd135628: dataIn1 = 32'd4835
; 
32'd135629: dataIn1 = 32'd1072
; 
32'd135630: dataIn1 = 32'd1073
; 
32'd135631: dataIn1 = 32'd2553
; 
32'd135632: dataIn1 = 32'd2555
; 
32'd135633: dataIn1 = 32'd2556
; 
32'd135634: dataIn1 = 32'd2557
; 
32'd135635: dataIn1 = 32'd3430
; 
32'd135636: dataIn1 = 32'd4645
; 
32'd135637: dataIn1 = 32'd4835
; 
32'd135638: dataIn1 = 32'd1072
; 
32'd135639: dataIn1 = 32'd2556
; 
32'd135640: dataIn1 = 32'd2557
; 
32'd135641: dataIn1 = 32'd4644
; 
32'd135642: dataIn1 = 32'd4645
; 
32'd135643: dataIn1 = 32'd4813
; 
32'd135644: dataIn1 = 32'd4815
; 
32'd135645: dataIn1 = 32'd2558
; 
32'd135646: dataIn1 = 32'd4648
; 
32'd135647: dataIn1 = 32'd4649
; 
32'd135648: dataIn1 = 32'd4653
; 
32'd135649: dataIn1 = 32'd4655
; 
32'd135650: dataIn1 = 32'd4657
; 
32'd135651: dataIn1 = 32'd4658
; 
32'd135652: dataIn1 = 32'd5892
; 
32'd135653: dataIn1 = 32'd5906
; 
32'd135654: dataIn1 = 32'd2559
; 
32'd135655: dataIn1 = 32'd4647
; 
32'd135656: dataIn1 = 32'd4649
; 
32'd135657: dataIn1 = 32'd4651
; 
32'd135658: dataIn1 = 32'd4654
; 
32'd135659: dataIn1 = 32'd4663
; 
32'd135660: dataIn1 = 32'd4665
; 
32'd135661: dataIn1 = 32'd5918
; 
32'd135662: dataIn1 = 32'd2560
; 
32'd135663: dataIn1 = 32'd4647
; 
32'd135664: dataIn1 = 32'd4648
; 
32'd135665: dataIn1 = 32'd4650
; 
32'd135666: dataIn1 = 32'd4652
; 
32'd135667: dataIn1 = 32'd4668
; 
32'd135668: dataIn1 = 32'd4669
; 
32'd135669: dataIn1 = 32'd5929
; 
32'd135670: dataIn1 = 32'd2561
; 
32'd135671: dataIn1 = 32'd5895
; 
32'd135672: dataIn1 = 32'd5896
; 
32'd135673: dataIn1 = 32'd5904
; 
32'd135674: dataIn1 = 32'd5913
; 
32'd135675: dataIn1 = 32'd5965
; 
32'd135676: dataIn1 = 32'd5966
; 
32'd135677: dataIn1 = 32'd2562
; 
32'd135678: dataIn1 = 32'd5897
; 
32'd135679: dataIn1 = 32'd5898
; 
32'd135680: dataIn1 = 32'd5905
; 
32'd135681: dataIn1 = 32'd5911
; 
32'd135682: dataIn1 = 32'd6028
; 
32'd135683: dataIn1 = 32'd6029
; 
32'd135684: dataIn1 = 32'd2563
; 
32'd135685: dataIn1 = 32'd4664
; 
32'd135686: dataIn1 = 32'd4665
; 
32'd135687: dataIn1 = 32'd4666
; 
32'd135688: dataIn1 = 32'd4667
; 
32'd135689: dataIn1 = 32'd4854
; 
32'd135690: dataIn1 = 32'd4855
; 
32'd135691: dataIn1 = 32'd5921
; 
32'd135692: dataIn1 = 32'd2564
; 
32'd135693: dataIn1 = 32'd4669
; 
32'd135694: dataIn1 = 32'd4670
; 
32'd135695: dataIn1 = 32'd4671
; 
32'd135696: dataIn1 = 32'd4672
; 
32'd135697: dataIn1 = 32'd4882
; 
32'd135698: dataIn1 = 32'd4883
; 
32'd135699: dataIn1 = 32'd5932
; 
32'd135700: dataIn1 = 32'd6061
; 
32'd135701: dataIn1 = 32'd212
; 
32'd135702: dataIn1 = 32'd1043
; 
32'd135703: dataIn1 = 32'd1077
; 
32'd135704: dataIn1 = 32'd2565
; 
32'd135705: dataIn1 = 32'd2566
; 
32'd135706: dataIn1 = 32'd2567
; 
32'd135707: dataIn1 = 32'd3431
; 
32'd135708: dataIn1 = 32'd4680
; 
32'd135709: dataIn1 = 32'd10274
; 
32'd135710: dataIn1 = 32'd10275
; 
32'd135711: dataIn1 = 32'd2565
; 
32'd135712: dataIn1 = 32'd2566
; 
32'd135713: dataIn1 = 32'd4673
; 
32'd135714: dataIn1 = 32'd4675
; 
32'd135715: dataIn1 = 32'd4677
; 
32'd135716: dataIn1 = 32'd4680
; 
32'd135717: dataIn1 = 32'd10274
; 
32'd135718: dataIn1 = 32'd2565
; 
32'd135719: dataIn1 = 32'd2567
; 
32'd135720: dataIn1 = 32'd10266
; 
32'd135721: dataIn1 = 32'd10267
; 
32'd135722: dataIn1 = 32'd10268
; 
32'd135723: dataIn1 = 32'd10274
; 
32'd135724: dataIn1 = 32'd10275
; 
32'd135725: dataIn1 = 32'd2568
; 
32'd135726: dataIn1 = 32'd4674
; 
32'd135727: dataIn1 = 32'd4675
; 
32'd135728: dataIn1 = 32'd4679
; 
32'd135729: dataIn1 = 32'd4681
; 
32'd135730: dataIn1 = 32'd4898
; 
32'd135731: dataIn1 = 32'd4899
; 
32'd135732: dataIn1 = 32'd2569
; 
32'd135733: dataIn1 = 32'd4673
; 
32'd135734: dataIn1 = 32'd4674
; 
32'd135735: dataIn1 = 32'd4676
; 
32'd135736: dataIn1 = 32'd4678
; 
32'd135737: dataIn1 = 32'd4857
; 
32'd135738: dataIn1 = 32'd4859
; 
32'd135739: dataIn1 = 32'd5992
; 
32'd135740: dataIn1 = 32'd2570
; 
32'd135741: dataIn1 = 32'd4682
; 
32'd135742: dataIn1 = 32'd4683
; 
32'd135743: dataIn1 = 32'd4853
; 
32'd135744: dataIn1 = 32'd4854
; 
32'd135745: dataIn1 = 32'd4856
; 
32'd135746: dataIn1 = 32'd10266
; 
32'd135747: dataIn1 = 32'd2571
; 
32'd135748: dataIn1 = 32'd3456
; 
32'd135749: dataIn1 = 32'd3466
; 
32'd135750: dataIn1 = 32'd4685
; 
32'd135751: dataIn1 = 32'd4686
; 
32'd135752: dataIn1 = 32'd4690
; 
32'd135753: dataIn1 = 32'd4692
; 
32'd135754: dataIn1 = 32'd2572
; 
32'd135755: dataIn1 = 32'd4684
; 
32'd135756: dataIn1 = 32'd4686
; 
32'd135757: dataIn1 = 32'd4688
; 
32'd135758: dataIn1 = 32'd4691
; 
32'd135759: dataIn1 = 32'd4912
; 
32'd135760: dataIn1 = 32'd4914
; 
32'd135761: dataIn1 = 32'd9630
; 
32'd135762: dataIn1 = 32'd2573
; 
32'd135763: dataIn1 = 32'd4684
; 
32'd135764: dataIn1 = 32'd4685
; 
32'd135765: dataIn1 = 32'd4687
; 
32'd135766: dataIn1 = 32'd4689
; 
32'd135767: dataIn1 = 32'd4893
; 
32'd135768: dataIn1 = 32'd4894
; 
32'd135769: dataIn1 = 32'd9619
; 
32'd135770: dataIn1 = 32'd2574
; 
32'd135771: dataIn1 = 32'd4694
; 
32'd135772: dataIn1 = 32'd4695
; 
32'd135773: dataIn1 = 32'd4699
; 
32'd135774: dataIn1 = 32'd4701
; 
32'd135775: dataIn1 = 32'd4936
; 
32'd135776: dataIn1 = 32'd4937
; 
32'd135777: dataIn1 = 32'd9661
; 
32'd135778: dataIn1 = 32'd2575
; 
32'd135779: dataIn1 = 32'd3481
; 
32'd135780: dataIn1 = 32'd3485
; 
32'd135781: dataIn1 = 32'd4693
; 
32'd135782: dataIn1 = 32'd4695
; 
32'd135783: dataIn1 = 32'd4697
; 
32'd135784: dataIn1 = 32'd4700
; 
32'd135785: dataIn1 = 32'd2576
; 
32'd135786: dataIn1 = 32'd4693
; 
32'd135787: dataIn1 = 32'd4694
; 
32'd135788: dataIn1 = 32'd4696
; 
32'd135789: dataIn1 = 32'd4698
; 
32'd135790: dataIn1 = 32'd4917
; 
32'd135791: dataIn1 = 32'd4919
; 
32'd135792: dataIn1 = 32'd9642
; 
32'd135793: dataIn1 = 32'd2577
; 
32'd135794: dataIn1 = 32'd3497
; 
32'd135795: dataIn1 = 32'd3500
; 
32'd135796: dataIn1 = 32'd4703
; 
32'd135797: dataIn1 = 32'd4704
; 
32'd135798: dataIn1 = 32'd4708
; 
32'd135799: dataIn1 = 32'd4710
; 
32'd135800: dataIn1 = 32'd2578
; 
32'd135801: dataIn1 = 32'd4702
; 
32'd135802: dataIn1 = 32'd4704
; 
32'd135803: dataIn1 = 32'd4706
; 
32'd135804: dataIn1 = 32'd4709
; 
32'd135805: dataIn1 = 32'd4950
; 
32'd135806: dataIn1 = 32'd4952
; 
32'd135807: dataIn1 = 32'd9666
; 
32'd135808: dataIn1 = 32'd2579
; 
32'd135809: dataIn1 = 32'd4702
; 
32'd135810: dataIn1 = 32'd4703
; 
32'd135811: dataIn1 = 32'd4705
; 
32'd135812: dataIn1 = 32'd4707
; 
32'd135813: dataIn1 = 32'd4931
; 
32'd135814: dataIn1 = 32'd4932
; 
32'd135815: dataIn1 = 32'd9652
; 
32'd135816: dataIn1 = 32'd2580
; 
32'd135817: dataIn1 = 32'd4712
; 
32'd135818: dataIn1 = 32'd4713
; 
32'd135819: dataIn1 = 32'd4717
; 
32'd135820: dataIn1 = 32'd4719
; 
32'd135821: dataIn1 = 32'd4974
; 
32'd135822: dataIn1 = 32'd4975
; 
32'd135823: dataIn1 = 32'd2581
; 
32'd135824: dataIn1 = 32'd3507
; 
32'd135825: dataIn1 = 32'd3509
; 
32'd135826: dataIn1 = 32'd4711
; 
32'd135827: dataIn1 = 32'd4713
; 
32'd135828: dataIn1 = 32'd4715
; 
32'd135829: dataIn1 = 32'd4718
; 
32'd135830: dataIn1 = 32'd2582
; 
32'd135831: dataIn1 = 32'd4711
; 
32'd135832: dataIn1 = 32'd4712
; 
32'd135833: dataIn1 = 32'd4714
; 
32'd135834: dataIn1 = 32'd4716
; 
32'd135835: dataIn1 = 32'd4955
; 
32'd135836: dataIn1 = 32'd4957
; 
32'd135837: dataIn1 = 32'd2583
; 
32'd135838: dataIn1 = 32'd3515
; 
32'd135839: dataIn1 = 32'd3517
; 
32'd135840: dataIn1 = 32'd4721
; 
32'd135841: dataIn1 = 32'd4722
; 
32'd135842: dataIn1 = 32'd4726
; 
32'd135843: dataIn1 = 32'd4728
; 
32'd135844: dataIn1 = 32'd2584
; 
32'd135845: dataIn1 = 32'd4720
; 
32'd135846: dataIn1 = 32'd4722
; 
32'd135847: dataIn1 = 32'd4724
; 
32'd135848: dataIn1 = 32'd4727
; 
32'd135849: dataIn1 = 32'd4988
; 
32'd135850: dataIn1 = 32'd4990
; 
32'd135851: dataIn1 = 32'd2585
; 
32'd135852: dataIn1 = 32'd4720
; 
32'd135853: dataIn1 = 32'd4721
; 
32'd135854: dataIn1 = 32'd4723
; 
32'd135855: dataIn1 = 32'd4725
; 
32'd135856: dataIn1 = 32'd4969
; 
32'd135857: dataIn1 = 32'd4970
; 
32'd135858: dataIn1 = 32'd2586
; 
32'd135859: dataIn1 = 32'd4730
; 
32'd135860: dataIn1 = 32'd4731
; 
32'd135861: dataIn1 = 32'd4735
; 
32'd135862: dataIn1 = 32'd4737
; 
32'd135863: dataIn1 = 32'd5012
; 
32'd135864: dataIn1 = 32'd5013
; 
32'd135865: dataIn1 = 32'd2587
; 
32'd135866: dataIn1 = 32'd3523
; 
32'd135867: dataIn1 = 32'd3525
; 
32'd135868: dataIn1 = 32'd4729
; 
32'd135869: dataIn1 = 32'd4731
; 
32'd135870: dataIn1 = 32'd4733
; 
32'd135871: dataIn1 = 32'd4736
; 
32'd135872: dataIn1 = 32'd2588
; 
32'd135873: dataIn1 = 32'd4729
; 
32'd135874: dataIn1 = 32'd4730
; 
32'd135875: dataIn1 = 32'd4732
; 
32'd135876: dataIn1 = 32'd4734
; 
32'd135877: dataIn1 = 32'd4993
; 
32'd135878: dataIn1 = 32'd4995
; 
32'd135879: dataIn1 = 32'd2589
; 
32'd135880: dataIn1 = 32'd3531
; 
32'd135881: dataIn1 = 32'd3533
; 
32'd135882: dataIn1 = 32'd4739
; 
32'd135883: dataIn1 = 32'd4740
; 
32'd135884: dataIn1 = 32'd4744
; 
32'd135885: dataIn1 = 32'd4746
; 
32'd135886: dataIn1 = 32'd2590
; 
32'd135887: dataIn1 = 32'd4738
; 
32'd135888: dataIn1 = 32'd4740
; 
32'd135889: dataIn1 = 32'd4742
; 
32'd135890: dataIn1 = 32'd4745
; 
32'd135891: dataIn1 = 32'd5026
; 
32'd135892: dataIn1 = 32'd5028
; 
32'd135893: dataIn1 = 32'd2591
; 
32'd135894: dataIn1 = 32'd4738
; 
32'd135895: dataIn1 = 32'd4739
; 
32'd135896: dataIn1 = 32'd4741
; 
32'd135897: dataIn1 = 32'd4743
; 
32'd135898: dataIn1 = 32'd5007
; 
32'd135899: dataIn1 = 32'd5008
; 
32'd135900: dataIn1 = 32'd2592
; 
32'd135901: dataIn1 = 32'd4748
; 
32'd135902: dataIn1 = 32'd4749
; 
32'd135903: dataIn1 = 32'd4753
; 
32'd135904: dataIn1 = 32'd4755
; 
32'd135905: dataIn1 = 32'd5050
; 
32'd135906: dataIn1 = 32'd5051
; 
32'd135907: dataIn1 = 32'd2593
; 
32'd135908: dataIn1 = 32'd3539
; 
32'd135909: dataIn1 = 32'd3541
; 
32'd135910: dataIn1 = 32'd4747
; 
32'd135911: dataIn1 = 32'd4749
; 
32'd135912: dataIn1 = 32'd4751
; 
32'd135913: dataIn1 = 32'd4754
; 
32'd135914: dataIn1 = 32'd2594
; 
32'd135915: dataIn1 = 32'd4747
; 
32'd135916: dataIn1 = 32'd4748
; 
32'd135917: dataIn1 = 32'd4750
; 
32'd135918: dataIn1 = 32'd4752
; 
32'd135919: dataIn1 = 32'd5031
; 
32'd135920: dataIn1 = 32'd5033
; 
32'd135921: dataIn1 = 32'd2595
; 
32'd135922: dataIn1 = 32'd3547
; 
32'd135923: dataIn1 = 32'd3549
; 
32'd135924: dataIn1 = 32'd4757
; 
32'd135925: dataIn1 = 32'd4758
; 
32'd135926: dataIn1 = 32'd4762
; 
32'd135927: dataIn1 = 32'd4764
; 
32'd135928: dataIn1 = 32'd2596
; 
32'd135929: dataIn1 = 32'd4756
; 
32'd135930: dataIn1 = 32'd4758
; 
32'd135931: dataIn1 = 32'd4760
; 
32'd135932: dataIn1 = 32'd4763
; 
32'd135933: dataIn1 = 32'd5064
; 
32'd135934: dataIn1 = 32'd5066
; 
32'd135935: dataIn1 = 32'd2597
; 
32'd135936: dataIn1 = 32'd4756
; 
32'd135937: dataIn1 = 32'd4757
; 
32'd135938: dataIn1 = 32'd4759
; 
32'd135939: dataIn1 = 32'd4761
; 
32'd135940: dataIn1 = 32'd5045
; 
32'd135941: dataIn1 = 32'd5046
; 
32'd135942: dataIn1 = 32'd2598
; 
32'd135943: dataIn1 = 32'd4766
; 
32'd135944: dataIn1 = 32'd4767
; 
32'd135945: dataIn1 = 32'd4771
; 
32'd135946: dataIn1 = 32'd4773
; 
32'd135947: dataIn1 = 32'd5088
; 
32'd135948: dataIn1 = 32'd5089
; 
32'd135949: dataIn1 = 32'd2599
; 
32'd135950: dataIn1 = 32'd3555
; 
32'd135951: dataIn1 = 32'd3557
; 
32'd135952: dataIn1 = 32'd4765
; 
32'd135953: dataIn1 = 32'd4767
; 
32'd135954: dataIn1 = 32'd4769
; 
32'd135955: dataIn1 = 32'd4772
; 
32'd135956: dataIn1 = 32'd2600
; 
32'd135957: dataIn1 = 32'd4765
; 
32'd135958: dataIn1 = 32'd4766
; 
32'd135959: dataIn1 = 32'd4768
; 
32'd135960: dataIn1 = 32'd4770
; 
32'd135961: dataIn1 = 32'd5069
; 
32'd135962: dataIn1 = 32'd5071
; 
32'd135963: dataIn1 = 32'd2601
; 
32'd135964: dataIn1 = 32'd3563
; 
32'd135965: dataIn1 = 32'd3565
; 
32'd135966: dataIn1 = 32'd4775
; 
32'd135967: dataIn1 = 32'd4776
; 
32'd135968: dataIn1 = 32'd4780
; 
32'd135969: dataIn1 = 32'd4782
; 
32'd135970: dataIn1 = 32'd2602
; 
32'd135971: dataIn1 = 32'd4774
; 
32'd135972: dataIn1 = 32'd4776
; 
32'd135973: dataIn1 = 32'd4778
; 
32'd135974: dataIn1 = 32'd4781
; 
32'd135975: dataIn1 = 32'd5102
; 
32'd135976: dataIn1 = 32'd5104
; 
32'd135977: dataIn1 = 32'd2603
; 
32'd135978: dataIn1 = 32'd4774
; 
32'd135979: dataIn1 = 32'd4775
; 
32'd135980: dataIn1 = 32'd4777
; 
32'd135981: dataIn1 = 32'd4779
; 
32'd135982: dataIn1 = 32'd5083
; 
32'd135983: dataIn1 = 32'd5084
; 
32'd135984: dataIn1 = 32'd2604
; 
32'd135985: dataIn1 = 32'd4784
; 
32'd135986: dataIn1 = 32'd4785
; 
32'd135987: dataIn1 = 32'd4789
; 
32'd135988: dataIn1 = 32'd4791
; 
32'd135989: dataIn1 = 32'd2605
; 
32'd135990: dataIn1 = 32'd3573
; 
32'd135991: dataIn1 = 32'd4783
; 
32'd135992: dataIn1 = 32'd4785
; 
32'd135993: dataIn1 = 32'd4787
; 
32'd135994: dataIn1 = 32'd4790
; 
32'd135995: dataIn1 = 32'd2606
; 
32'd135996: dataIn1 = 32'd4783
; 
32'd135997: dataIn1 = 32'd4784
; 
32'd135998: dataIn1 = 32'd4786
; 
32'd135999: dataIn1 = 32'd4788
; 
32'd136000: dataIn1 = 32'd5107
; 
32'd136001: dataIn1 = 32'd5109
; 
32'd136002: dataIn1 = 32'd1070
; 
32'd136003: dataIn1 = 32'd2607
; 
32'd136004: dataIn1 = 32'd2609
; 
32'd136005: dataIn1 = 32'd4793
; 
32'd136006: dataIn1 = 32'd4794
; 
32'd136007: dataIn1 = 32'd4796
; 
32'd136008: dataIn1 = 32'd4797
; 
32'd136009: dataIn1 = 32'd1069
; 
32'd136010: dataIn1 = 32'd2608
; 
32'd136011: dataIn1 = 32'd2609
; 
32'd136012: dataIn1 = 32'd4792
; 
32'd136013: dataIn1 = 32'd4794
; 
32'd136014: dataIn1 = 32'd4800
; 
32'd136015: dataIn1 = 32'd4802
; 
32'd136016: dataIn1 = 32'd1069
; 
32'd136017: dataIn1 = 32'd1070
; 
32'd136018: dataIn1 = 32'd2607
; 
32'd136019: dataIn1 = 32'd2608
; 
32'd136020: dataIn1 = 32'd2609
; 
32'd136021: dataIn1 = 32'd3480
; 
32'd136022: dataIn1 = 32'd3484
; 
32'd136023: dataIn1 = 32'd4794
; 
32'd136024: dataIn1 = 32'd2610
; 
32'd136025: dataIn1 = 32'd4795
; 
32'd136026: dataIn1 = 32'd4797
; 
32'd136027: dataIn1 = 32'd9698
; 
32'd136028: dataIn1 = 32'd9699
; 
32'd136029: dataIn1 = 32'd9703
; 
32'd136030: dataIn1 = 32'd9708
; 
32'd136031: dataIn1 = 32'd2611
; 
32'd136032: dataIn1 = 32'd4801
; 
32'd136033: dataIn1 = 32'd4802
; 
32'd136034: dataIn1 = 32'd9683
; 
32'd136035: dataIn1 = 32'd9685
; 
32'd136036: dataIn1 = 32'd9691
; 
32'd136037: dataIn1 = 32'd9695
; 
32'd136038: dataIn1 = 32'd1071
; 
32'd136039: dataIn1 = 32'd2612
; 
32'd136040: dataIn1 = 32'd2613
; 
32'd136041: dataIn1 = 32'd4806
; 
32'd136042: dataIn1 = 32'd4807
; 
32'd136043: dataIn1 = 32'd4809
; 
32'd136044: dataIn1 = 32'd4810
; 
32'd136045: dataIn1 = 32'd1071
; 
32'd136046: dataIn1 = 32'd1072
; 
32'd136047: dataIn1 = 32'd2612
; 
32'd136048: dataIn1 = 32'd2613
; 
32'd136049: dataIn1 = 32'd2614
; 
32'd136050: dataIn1 = 32'd3455
; 
32'd136051: dataIn1 = 32'd3465
; 
32'd136052: dataIn1 = 32'd4806
; 
32'd136053: dataIn1 = 32'd1072
; 
32'd136054: dataIn1 = 32'd2613
; 
32'd136055: dataIn1 = 32'd2614
; 
32'd136056: dataIn1 = 32'd4805
; 
32'd136057: dataIn1 = 32'd4806
; 
32'd136058: dataIn1 = 32'd4813
; 
32'd136059: dataIn1 = 32'd4814
; 
32'd136060: dataIn1 = 32'd2615
; 
32'd136061: dataIn1 = 32'd4808
; 
32'd136062: dataIn1 = 32'd4809
; 
32'd136063: dataIn1 = 32'd9713
; 
32'd136064: dataIn1 = 32'd9714
; 
32'd136065: dataIn1 = 32'd9720
; 
32'd136066: dataIn1 = 32'd9725
; 
32'd136067: dataIn1 = 32'd2616
; 
32'd136068: dataIn1 = 32'd4814
; 
32'd136069: dataIn1 = 32'd4815
; 
32'd136070: dataIn1 = 32'd4817
; 
32'd136071: dataIn1 = 32'd9730
; 
32'd136072: dataIn1 = 32'd9731
; 
32'd136073: dataIn1 = 32'd9758
; 
32'd136074: dataIn1 = 32'd2617
; 
32'd136075: dataIn1 = 32'd4819
; 
32'd136076: dataIn1 = 32'd4820
; 
32'd136077: dataIn1 = 32'd4824
; 
32'd136078: dataIn1 = 32'd4826
; 
32'd136079: dataIn1 = 32'd4828
; 
32'd136080: dataIn1 = 32'd4829
; 
32'd136081: dataIn1 = 32'd2618
; 
32'd136082: dataIn1 = 32'd4818
; 
32'd136083: dataIn1 = 32'd4820
; 
32'd136084: dataIn1 = 32'd4822
; 
32'd136085: dataIn1 = 32'd4825
; 
32'd136086: dataIn1 = 32'd4832
; 
32'd136087: dataIn1 = 32'd4834
; 
32'd136088: dataIn1 = 32'd2619
; 
32'd136089: dataIn1 = 32'd4818
; 
32'd136090: dataIn1 = 32'd4819
; 
32'd136091: dataIn1 = 32'd4821
; 
32'd136092: dataIn1 = 32'd4823
; 
32'd136093: dataIn1 = 32'd5318
; 
32'd136094: dataIn1 = 32'd5430
; 
32'd136095: dataIn1 = 32'd2620
; 
32'd136096: dataIn1 = 32'd4829
; 
32'd136097: dataIn1 = 32'd5945
; 
32'd136098: dataIn1 = 32'd5946
; 
32'd136099: dataIn1 = 32'd6955
; 
32'd136100: dataIn1 = 32'd6956
; 
32'd136101: dataIn1 = 32'd6970
; 
32'd136102: dataIn1 = 32'd2621
; 
32'd136103: dataIn1 = 32'd4833
; 
32'd136104: dataIn1 = 32'd4834
; 
32'd136105: dataIn1 = 32'd4836
; 
32'd136106: dataIn1 = 32'd4837
; 
32'd136107: dataIn1 = 32'd5858
; 
32'd136108: dataIn1 = 32'd5860
; 
32'd136109: dataIn1 = 32'd6938
; 
32'd136110: dataIn1 = 32'd2622
; 
32'd136111: dataIn1 = 32'd4841
; 
32'd136112: dataIn1 = 32'd4847
; 
32'd136113: dataIn1 = 32'd5956
; 
32'd136114: dataIn1 = 32'd5957
; 
32'd136115: dataIn1 = 32'd5963
; 
32'd136116: dataIn1 = 32'd5964
; 
32'd136117: dataIn1 = 32'd2623
; 
32'd136118: dataIn1 = 32'd4839
; 
32'd136119: dataIn1 = 32'd4841
; 
32'd136120: dataIn1 = 32'd4843
; 
32'd136121: dataIn1 = 32'd4846
; 
32'd136122: dataIn1 = 32'd4853
; 
32'd136123: dataIn1 = 32'd4855
; 
32'd136124: dataIn1 = 32'd2624
; 
32'd136125: dataIn1 = 32'd4839
; 
32'd136126: dataIn1 = 32'd4840
; 
32'd136127: dataIn1 = 32'd4842
; 
32'd136128: dataIn1 = 32'd4844
; 
32'd136129: dataIn1 = 32'd4857
; 
32'd136130: dataIn1 = 32'd4858
; 
32'd136131: dataIn1 = 32'd5955
; 
32'd136132: dataIn1 = 32'd5988
; 
32'd136133: dataIn1 = 32'd2625
; 
32'd136134: dataIn1 = 32'd5967
; 
32'd136135: dataIn1 = 32'd5968
; 
32'd136136: dataIn1 = 32'd5973
; 
32'd136137: dataIn1 = 32'd5978
; 
32'd136138: dataIn1 = 32'd7324
; 
32'd136139: dataIn1 = 32'd7325
; 
32'd136140: dataIn1 = 32'd2626
; 
32'd136141: dataIn1 = 32'd5984
; 
32'd136142: dataIn1 = 32'd5985
; 
32'd136143: dataIn1 = 32'd5989
; 
32'd136144: dataIn1 = 32'd5994
; 
32'd136145: dataIn1 = 32'd7340
; 
32'd136146: dataIn1 = 32'd7341
; 
32'd136147: dataIn1 = 32'd2627
; 
32'd136148: dataIn1 = 32'd5999
; 
32'd136149: dataIn1 = 32'd6000
; 
32'd136150: dataIn1 = 32'd6012
; 
32'd136151: dataIn1 = 32'd6017
; 
32'd136152: dataIn1 = 32'd6024
; 
32'd136153: dataIn1 = 32'd6025
; 
32'd136154: dataIn1 = 32'd2628
; 
32'd136155: dataIn1 = 32'd6001
; 
32'd136156: dataIn1 = 32'd6002
; 
32'd136157: dataIn1 = 32'd6005
; 
32'd136158: dataIn1 = 32'd6018
; 
32'd136159: dataIn1 = 32'd6046
; 
32'd136160: dataIn1 = 32'd6048
; 
32'd136161: dataIn1 = 32'd2629
; 
32'd136162: dataIn1 = 32'd4881
; 
32'd136163: dataIn1 = 32'd4882
; 
32'd136164: dataIn1 = 32'd6003
; 
32'd136165: dataIn1 = 32'd6004
; 
32'd136166: dataIn1 = 32'd6007
; 
32'd136167: dataIn1 = 32'd6013
; 
32'd136168: dataIn1 = 32'd2630
; 
32'd136169: dataIn1 = 32'd6026
; 
32'd136170: dataIn1 = 32'd6027
; 
32'd136171: dataIn1 = 32'd6034
; 
32'd136172: dataIn1 = 32'd6041
; 
32'd136173: dataIn1 = 32'd7266
; 
32'd136174: dataIn1 = 32'd7267
; 
32'd136175: dataIn1 = 32'd2631
; 
32'd136176: dataIn1 = 32'd6044
; 
32'd136177: dataIn1 = 32'd6045
; 
32'd136178: dataIn1 = 32'd6059
; 
32'd136179: dataIn1 = 32'd6703
; 
32'd136180: dataIn1 = 32'd9232
; 
32'd136181: dataIn1 = 32'd9274
; 
32'd136182: dataIn1 = 32'd2632
; 
32'd136183: dataIn1 = 32'd4885
; 
32'd136184: dataIn1 = 32'd4886
; 
32'd136185: dataIn1 = 32'd4890
; 
32'd136186: dataIn1 = 32'd4892
; 
32'd136187: dataIn1 = 32'd4894
; 
32'd136188: dataIn1 = 32'd4895
; 
32'd136189: dataIn1 = 32'd9620
; 
32'd136190: dataIn1 = 32'd2633
; 
32'd136191: dataIn1 = 32'd4884
; 
32'd136192: dataIn1 = 32'd4886
; 
32'd136193: dataIn1 = 32'd4888
; 
32'd136194: dataIn1 = 32'd4891
; 
32'd136195: dataIn1 = 32'd4898
; 
32'd136196: dataIn1 = 32'd4900
; 
32'd136197: dataIn1 = 32'd2634
; 
32'd136198: dataIn1 = 32'd3431
; 
32'd136199: dataIn1 = 32'd3432
; 
32'd136200: dataIn1 = 32'd4884
; 
32'd136201: dataIn1 = 32'd4885
; 
32'd136202: dataIn1 = 32'd4887
; 
32'd136203: dataIn1 = 32'd4889
; 
32'd136204: dataIn1 = 32'd2635
; 
32'd136205: dataIn1 = 32'd7476
; 
32'd136206: dataIn1 = 32'd7477
; 
32'd136207: dataIn1 = 32'd7488
; 
32'd136208: dataIn1 = 32'd7493
; 
32'd136209: dataIn1 = 32'd9614
; 
32'd136210: dataIn1 = 32'd9616
; 
32'd136211: dataIn1 = 32'd2636
; 
32'd136212: dataIn1 = 32'd4899
; 
32'd136213: dataIn1 = 32'd4900
; 
32'd136214: dataIn1 = 32'd7454
; 
32'd136215: dataIn1 = 32'd7455
; 
32'd136216: dataIn1 = 32'd7461
; 
32'd136217: dataIn1 = 32'd7471
; 
32'd136218: dataIn1 = 32'd2637
; 
32'd136219: dataIn1 = 32'd4904
; 
32'd136220: dataIn1 = 32'd4905
; 
32'd136221: dataIn1 = 32'd4909
; 
32'd136222: dataIn1 = 32'd4911
; 
32'd136223: dataIn1 = 32'd4913
; 
32'd136224: dataIn1 = 32'd4914
; 
32'd136225: dataIn1 = 32'd9632
; 
32'd136226: dataIn1 = 32'd2638
; 
32'd136227: dataIn1 = 32'd3473
; 
32'd136228: dataIn1 = 32'd3477
; 
32'd136229: dataIn1 = 32'd4903
; 
32'd136230: dataIn1 = 32'd4905
; 
32'd136231: dataIn1 = 32'd4907
; 
32'd136232: dataIn1 = 32'd4910
; 
32'd136233: dataIn1 = 32'd2639
; 
32'd136234: dataIn1 = 32'd4903
; 
32'd136235: dataIn1 = 32'd4904
; 
32'd136236: dataIn1 = 32'd4906
; 
32'd136237: dataIn1 = 32'd4908
; 
32'd136238: dataIn1 = 32'd4917
; 
32'd136239: dataIn1 = 32'd4918
; 
32'd136240: dataIn1 = 32'd9640
; 
32'd136241: dataIn1 = 32'd2640
; 
32'd136242: dataIn1 = 32'd7566
; 
32'd136243: dataIn1 = 32'd7567
; 
32'd136244: dataIn1 = 32'd7572
; 
32'd136245: dataIn1 = 32'd7577
; 
32'd136246: dataIn1 = 32'd9626
; 
32'd136247: dataIn1 = 32'd9627
; 
32'd136248: dataIn1 = 32'd2641
; 
32'd136249: dataIn1 = 32'd7586
; 
32'd136250: dataIn1 = 32'd7587
; 
32'd136251: dataIn1 = 32'd7594
; 
32'd136252: dataIn1 = 32'd7604
; 
32'd136253: dataIn1 = 32'd9636
; 
32'd136254: dataIn1 = 32'd9637
; 
32'd136255: dataIn1 = 32'd2642
; 
32'd136256: dataIn1 = 32'd4923
; 
32'd136257: dataIn1 = 32'd4924
; 
32'd136258: dataIn1 = 32'd4928
; 
32'd136259: dataIn1 = 32'd4930
; 
32'd136260: dataIn1 = 32'd4932
; 
32'd136261: dataIn1 = 32'd4933
; 
32'd136262: dataIn1 = 32'd9653
; 
32'd136263: dataIn1 = 32'd2643
; 
32'd136264: dataIn1 = 32'd4922
; 
32'd136265: dataIn1 = 32'd4924
; 
32'd136266: dataIn1 = 32'd4926
; 
32'd136267: dataIn1 = 32'd4929
; 
32'd136268: dataIn1 = 32'd4936
; 
32'd136269: dataIn1 = 32'd4938
; 
32'd136270: dataIn1 = 32'd9663
; 
32'd136271: dataIn1 = 32'd2644
; 
32'd136272: dataIn1 = 32'd3489
; 
32'd136273: dataIn1 = 32'd3493
; 
32'd136274: dataIn1 = 32'd4922
; 
32'd136275: dataIn1 = 32'd4923
; 
32'd136276: dataIn1 = 32'd4925
; 
32'd136277: dataIn1 = 32'd4927
; 
32'd136278: dataIn1 = 32'd2645
; 
32'd136279: dataIn1 = 32'd7729
; 
32'd136280: dataIn1 = 32'd7730
; 
32'd136281: dataIn1 = 32'd7741
; 
32'd136282: dataIn1 = 32'd7746
; 
32'd136283: dataIn1 = 32'd9647
; 
32'd136284: dataIn1 = 32'd9649
; 
32'd136285: dataIn1 = 32'd2646
; 
32'd136286: dataIn1 = 32'd7705
; 
32'd136287: dataIn1 = 32'd7706
; 
32'd136288: dataIn1 = 32'd7714
; 
32'd136289: dataIn1 = 32'd7724
; 
32'd136290: dataIn1 = 32'd9657
; 
32'd136291: dataIn1 = 32'd9658
; 
32'd136292: dataIn1 = 32'd2647
; 
32'd136293: dataIn1 = 32'd4942
; 
32'd136294: dataIn1 = 32'd4943
; 
32'd136295: dataIn1 = 32'd4947
; 
32'd136296: dataIn1 = 32'd4949
; 
32'd136297: dataIn1 = 32'd4951
; 
32'd136298: dataIn1 = 32'd4952
; 
32'd136299: dataIn1 = 32'd2648
; 
32'd136300: dataIn1 = 32'd3503
; 
32'd136301: dataIn1 = 32'd3505
; 
32'd136302: dataIn1 = 32'd4941
; 
32'd136303: dataIn1 = 32'd4943
; 
32'd136304: dataIn1 = 32'd4945
; 
32'd136305: dataIn1 = 32'd4948
; 
32'd136306: dataIn1 = 32'd2649
; 
32'd136307: dataIn1 = 32'd4941
; 
32'd136308: dataIn1 = 32'd4942
; 
32'd136309: dataIn1 = 32'd4944
; 
32'd136310: dataIn1 = 32'd4946
; 
32'd136311: dataIn1 = 32'd4955
; 
32'd136312: dataIn1 = 32'd4956
; 
32'd136313: dataIn1 = 32'd2650
; 
32'd136314: dataIn1 = 32'd4951
; 
32'd136315: dataIn1 = 32'd7819
; 
32'd136316: dataIn1 = 32'd7820
; 
32'd136317: dataIn1 = 32'd7825
; 
32'd136318: dataIn1 = 32'd7830
; 
32'd136319: dataIn1 = 32'd9764
; 
32'd136320: dataIn1 = 32'd2651
; 
32'd136321: dataIn1 = 32'd4956
; 
32'd136322: dataIn1 = 32'd4957
; 
32'd136323: dataIn1 = 32'd7839
; 
32'd136324: dataIn1 = 32'd7840
; 
32'd136325: dataIn1 = 32'd7847
; 
32'd136326: dataIn1 = 32'd7857
; 
32'd136327: dataIn1 = 32'd2652
; 
32'd136328: dataIn1 = 32'd4961
; 
32'd136329: dataIn1 = 32'd4962
; 
32'd136330: dataIn1 = 32'd4966
; 
32'd136331: dataIn1 = 32'd4968
; 
32'd136332: dataIn1 = 32'd4970
; 
32'd136333: dataIn1 = 32'd4971
; 
32'd136334: dataIn1 = 32'd2653
; 
32'd136335: dataIn1 = 32'd4960
; 
32'd136336: dataIn1 = 32'd4962
; 
32'd136337: dataIn1 = 32'd4964
; 
32'd136338: dataIn1 = 32'd4967
; 
32'd136339: dataIn1 = 32'd4974
; 
32'd136340: dataIn1 = 32'd4976
; 
32'd136341: dataIn1 = 32'd2654
; 
32'd136342: dataIn1 = 32'd3511
; 
32'd136343: dataIn1 = 32'd3513
; 
32'd136344: dataIn1 = 32'd4960
; 
32'd136345: dataIn1 = 32'd4961
; 
32'd136346: dataIn1 = 32'd4963
; 
32'd136347: dataIn1 = 32'd4965
; 
32'd136348: dataIn1 = 32'd2655
; 
32'd136349: dataIn1 = 32'd4969
; 
32'd136350: dataIn1 = 32'd4971
; 
32'd136351: dataIn1 = 32'd7982
; 
32'd136352: dataIn1 = 32'd7983
; 
32'd136353: dataIn1 = 32'd7994
; 
32'd136354: dataIn1 = 32'd7999
; 
32'd136355: dataIn1 = 32'd2656
; 
32'd136356: dataIn1 = 32'd4975
; 
32'd136357: dataIn1 = 32'd4976
; 
32'd136358: dataIn1 = 32'd7958
; 
32'd136359: dataIn1 = 32'd7959
; 
32'd136360: dataIn1 = 32'd7967
; 
32'd136361: dataIn1 = 32'd7977
; 
32'd136362: dataIn1 = 32'd2657
; 
32'd136363: dataIn1 = 32'd4980
; 
32'd136364: dataIn1 = 32'd4981
; 
32'd136365: dataIn1 = 32'd4985
; 
32'd136366: dataIn1 = 32'd4987
; 
32'd136367: dataIn1 = 32'd4989
; 
32'd136368: dataIn1 = 32'd4990
; 
32'd136369: dataIn1 = 32'd2658
; 
32'd136370: dataIn1 = 32'd3519
; 
32'd136371: dataIn1 = 32'd3521
; 
32'd136372: dataIn1 = 32'd4979
; 
32'd136373: dataIn1 = 32'd4981
; 
32'd136374: dataIn1 = 32'd4983
; 
32'd136375: dataIn1 = 32'd4986
; 
32'd136376: dataIn1 = 32'd2659
; 
32'd136377: dataIn1 = 32'd4979
; 
32'd136378: dataIn1 = 32'd4980
; 
32'd136379: dataIn1 = 32'd4982
; 
32'd136380: dataIn1 = 32'd4984
; 
32'd136381: dataIn1 = 32'd4993
; 
32'd136382: dataIn1 = 32'd4994
; 
32'd136383: dataIn1 = 32'd2660
; 
32'd136384: dataIn1 = 32'd4988
; 
32'd136385: dataIn1 = 32'd4989
; 
32'd136386: dataIn1 = 32'd8072
; 
32'd136387: dataIn1 = 32'd8073
; 
32'd136388: dataIn1 = 32'd8078
; 
32'd136389: dataIn1 = 32'd8083
; 
32'd136390: dataIn1 = 32'd2661
; 
32'd136391: dataIn1 = 32'd4994
; 
32'd136392: dataIn1 = 32'd4995
; 
32'd136393: dataIn1 = 32'd8092
; 
32'd136394: dataIn1 = 32'd8093
; 
32'd136395: dataIn1 = 32'd8100
; 
32'd136396: dataIn1 = 32'd8110
; 
32'd136397: dataIn1 = 32'd2662
; 
32'd136398: dataIn1 = 32'd4999
; 
32'd136399: dataIn1 = 32'd5000
; 
32'd136400: dataIn1 = 32'd5004
; 
32'd136401: dataIn1 = 32'd5006
; 
32'd136402: dataIn1 = 32'd5008
; 
32'd136403: dataIn1 = 32'd5009
; 
32'd136404: dataIn1 = 32'd2663
; 
32'd136405: dataIn1 = 32'd4998
; 
32'd136406: dataIn1 = 32'd5000
; 
32'd136407: dataIn1 = 32'd5002
; 
32'd136408: dataIn1 = 32'd5005
; 
32'd136409: dataIn1 = 32'd5012
; 
32'd136410: dataIn1 = 32'd5014
; 
32'd136411: dataIn1 = 32'd2664
; 
32'd136412: dataIn1 = 32'd3527
; 
32'd136413: dataIn1 = 32'd3529
; 
32'd136414: dataIn1 = 32'd4998
; 
32'd136415: dataIn1 = 32'd4999
; 
32'd136416: dataIn1 = 32'd5001
; 
32'd136417: dataIn1 = 32'd5003
; 
32'd136418: dataIn1 = 32'd2665
; 
32'd136419: dataIn1 = 32'd5007
; 
32'd136420: dataIn1 = 32'd5009
; 
32'd136421: dataIn1 = 32'd8235
; 
32'd136422: dataIn1 = 32'd8236
; 
32'd136423: dataIn1 = 32'd8247
; 
32'd136424: dataIn1 = 32'd8252
; 
32'd136425: dataIn1 = 32'd2666
; 
32'd136426: dataIn1 = 32'd5013
; 
32'd136427: dataIn1 = 32'd5014
; 
32'd136428: dataIn1 = 32'd8211
; 
32'd136429: dataIn1 = 32'd8212
; 
32'd136430: dataIn1 = 32'd8220
; 
32'd136431: dataIn1 = 32'd8230
; 
32'd136432: dataIn1 = 32'd2667
; 
32'd136433: dataIn1 = 32'd5018
; 
32'd136434: dataIn1 = 32'd5019
; 
32'd136435: dataIn1 = 32'd5023
; 
32'd136436: dataIn1 = 32'd5025
; 
32'd136437: dataIn1 = 32'd5027
; 
32'd136438: dataIn1 = 32'd5028
; 
32'd136439: dataIn1 = 32'd2668
; 
32'd136440: dataIn1 = 32'd3535
; 
32'd136441: dataIn1 = 32'd3537
; 
32'd136442: dataIn1 = 32'd5017
; 
32'd136443: dataIn1 = 32'd5019
; 
32'd136444: dataIn1 = 32'd5021
; 
32'd136445: dataIn1 = 32'd5024
; 
32'd136446: dataIn1 = 32'd2669
; 
32'd136447: dataIn1 = 32'd5017
; 
32'd136448: dataIn1 = 32'd5018
; 
32'd136449: dataIn1 = 32'd5020
; 
32'd136450: dataIn1 = 32'd5022
; 
32'd136451: dataIn1 = 32'd5031
; 
32'd136452: dataIn1 = 32'd5032
; 
32'd136453: dataIn1 = 32'd2670
; 
32'd136454: dataIn1 = 32'd5026
; 
32'd136455: dataIn1 = 32'd5027
; 
32'd136456: dataIn1 = 32'd8324
; 
32'd136457: dataIn1 = 32'd8325
; 
32'd136458: dataIn1 = 32'd8330
; 
32'd136459: dataIn1 = 32'd8335
; 
32'd136460: dataIn1 = 32'd2671
; 
32'd136461: dataIn1 = 32'd5032
; 
32'd136462: dataIn1 = 32'd5033
; 
32'd136463: dataIn1 = 32'd8344
; 
32'd136464: dataIn1 = 32'd8345
; 
32'd136465: dataIn1 = 32'd8352
; 
32'd136466: dataIn1 = 32'd8362
; 
32'd136467: dataIn1 = 32'd2672
; 
32'd136468: dataIn1 = 32'd5037
; 
32'd136469: dataIn1 = 32'd5038
; 
32'd136470: dataIn1 = 32'd5042
; 
32'd136471: dataIn1 = 32'd5044
; 
32'd136472: dataIn1 = 32'd5046
; 
32'd136473: dataIn1 = 32'd5047
; 
32'd136474: dataIn1 = 32'd2673
; 
32'd136475: dataIn1 = 32'd5036
; 
32'd136476: dataIn1 = 32'd5038
; 
32'd136477: dataIn1 = 32'd5040
; 
32'd136478: dataIn1 = 32'd5043
; 
32'd136479: dataIn1 = 32'd5050
; 
32'd136480: dataIn1 = 32'd5052
; 
32'd136481: dataIn1 = 32'd2674
; 
32'd136482: dataIn1 = 32'd3543
; 
32'd136483: dataIn1 = 32'd3545
; 
32'd136484: dataIn1 = 32'd5036
; 
32'd136485: dataIn1 = 32'd5037
; 
32'd136486: dataIn1 = 32'd5039
; 
32'd136487: dataIn1 = 32'd5041
; 
32'd136488: dataIn1 = 32'd2675
; 
32'd136489: dataIn1 = 32'd5045
; 
32'd136490: dataIn1 = 32'd5047
; 
32'd136491: dataIn1 = 32'd8487
; 
32'd136492: dataIn1 = 32'd8488
; 
32'd136493: dataIn1 = 32'd8499
; 
32'd136494: dataIn1 = 32'd8504
; 
32'd136495: dataIn1 = 32'd2676
; 
32'd136496: dataIn1 = 32'd5051
; 
32'd136497: dataIn1 = 32'd5052
; 
32'd136498: dataIn1 = 32'd8463
; 
32'd136499: dataIn1 = 32'd8464
; 
32'd136500: dataIn1 = 32'd8472
; 
32'd136501: dataIn1 = 32'd8482
; 
32'd136502: dataIn1 = 32'd2677
; 
32'd136503: dataIn1 = 32'd5056
; 
32'd136504: dataIn1 = 32'd5057
; 
32'd136505: dataIn1 = 32'd5061
; 
32'd136506: dataIn1 = 32'd5063
; 
32'd136507: dataIn1 = 32'd5065
; 
32'd136508: dataIn1 = 32'd5066
; 
32'd136509: dataIn1 = 32'd2678
; 
32'd136510: dataIn1 = 32'd3551
; 
32'd136511: dataIn1 = 32'd3553
; 
32'd136512: dataIn1 = 32'd5055
; 
32'd136513: dataIn1 = 32'd5057
; 
32'd136514: dataIn1 = 32'd5059
; 
32'd136515: dataIn1 = 32'd5062
; 
32'd136516: dataIn1 = 32'd2679
; 
32'd136517: dataIn1 = 32'd5055
; 
32'd136518: dataIn1 = 32'd5056
; 
32'd136519: dataIn1 = 32'd5058
; 
32'd136520: dataIn1 = 32'd5060
; 
32'd136521: dataIn1 = 32'd5069
; 
32'd136522: dataIn1 = 32'd5070
; 
32'd136523: dataIn1 = 32'd2680
; 
32'd136524: dataIn1 = 32'd5064
; 
32'd136525: dataIn1 = 32'd5065
; 
32'd136526: dataIn1 = 32'd8577
; 
32'd136527: dataIn1 = 32'd8578
; 
32'd136528: dataIn1 = 32'd8583
; 
32'd136529: dataIn1 = 32'd8588
; 
32'd136530: dataIn1 = 32'd2681
; 
32'd136531: dataIn1 = 32'd5070
; 
32'd136532: dataIn1 = 32'd5071
; 
32'd136533: dataIn1 = 32'd8597
; 
32'd136534: dataIn1 = 32'd8598
; 
32'd136535: dataIn1 = 32'd8605
; 
32'd136536: dataIn1 = 32'd8615
; 
32'd136537: dataIn1 = 32'd2682
; 
32'd136538: dataIn1 = 32'd5075
; 
32'd136539: dataIn1 = 32'd5076
; 
32'd136540: dataIn1 = 32'd5080
; 
32'd136541: dataIn1 = 32'd5082
; 
32'd136542: dataIn1 = 32'd5084
; 
32'd136543: dataIn1 = 32'd5085
; 
32'd136544: dataIn1 = 32'd2683
; 
32'd136545: dataIn1 = 32'd5074
; 
32'd136546: dataIn1 = 32'd5076
; 
32'd136547: dataIn1 = 32'd5078
; 
32'd136548: dataIn1 = 32'd5081
; 
32'd136549: dataIn1 = 32'd5088
; 
32'd136550: dataIn1 = 32'd5090
; 
32'd136551: dataIn1 = 32'd2684
; 
32'd136552: dataIn1 = 32'd3559
; 
32'd136553: dataIn1 = 32'd3561
; 
32'd136554: dataIn1 = 32'd5074
; 
32'd136555: dataIn1 = 32'd5075
; 
32'd136556: dataIn1 = 32'd5077
; 
32'd136557: dataIn1 = 32'd5079
; 
32'd136558: dataIn1 = 32'd2685
; 
32'd136559: dataIn1 = 32'd5083
; 
32'd136560: dataIn1 = 32'd5085
; 
32'd136561: dataIn1 = 32'd8740
; 
32'd136562: dataIn1 = 32'd8741
; 
32'd136563: dataIn1 = 32'd8752
; 
32'd136564: dataIn1 = 32'd8757
; 
32'd136565: dataIn1 = 32'd2686
; 
32'd136566: dataIn1 = 32'd5089
; 
32'd136567: dataIn1 = 32'd5090
; 
32'd136568: dataIn1 = 32'd8716
; 
32'd136569: dataIn1 = 32'd8717
; 
32'd136570: dataIn1 = 32'd8725
; 
32'd136571: dataIn1 = 32'd8735
; 
32'd136572: dataIn1 = 32'd2687
; 
32'd136573: dataIn1 = 32'd5094
; 
32'd136574: dataIn1 = 32'd5095
; 
32'd136575: dataIn1 = 32'd5099
; 
32'd136576: dataIn1 = 32'd5101
; 
32'd136577: dataIn1 = 32'd5103
; 
32'd136578: dataIn1 = 32'd5104
; 
32'd136579: dataIn1 = 32'd2688
; 
32'd136580: dataIn1 = 32'd3567
; 
32'd136581: dataIn1 = 32'd3569
; 
32'd136582: dataIn1 = 32'd5093
; 
32'd136583: dataIn1 = 32'd5095
; 
32'd136584: dataIn1 = 32'd5097
; 
32'd136585: dataIn1 = 32'd5100
; 
32'd136586: dataIn1 = 32'd2689
; 
32'd136587: dataIn1 = 32'd5093
; 
32'd136588: dataIn1 = 32'd5094
; 
32'd136589: dataIn1 = 32'd5096
; 
32'd136590: dataIn1 = 32'd5098
; 
32'd136591: dataIn1 = 32'd5107
; 
32'd136592: dataIn1 = 32'd5108
; 
32'd136593: dataIn1 = 32'd2690
; 
32'd136594: dataIn1 = 32'd5102
; 
32'd136595: dataIn1 = 32'd5103
; 
32'd136596: dataIn1 = 32'd8829
; 
32'd136597: dataIn1 = 32'd8830
; 
32'd136598: dataIn1 = 32'd8835
; 
32'd136599: dataIn1 = 32'd8840
; 
32'd136600: dataIn1 = 32'd2691
; 
32'd136601: dataIn1 = 32'd5108
; 
32'd136602: dataIn1 = 32'd5109
; 
32'd136603: dataIn1 = 32'd8849
; 
32'd136604: dataIn1 = 32'd8850
; 
32'd136605: dataIn1 = 32'd8857
; 
32'd136606: dataIn1 = 32'd8867
; 
32'd136607: dataIn1 = 32'd2692
; 
32'd136608: dataIn1 = 32'd7067
; 
32'd136609: dataIn1 = 32'd7068
; 
32'd136610: dataIn1 = 32'd7097
; 
32'd136611: dataIn1 = 32'd7107
; 
32'd136612: dataIn1 = 32'd7123
; 
32'd136613: dataIn1 = 32'd7124
; 
32'd136614: dataIn1 = 32'd2693
; 
32'd136615: dataIn1 = 32'd6072
; 
32'd136616: dataIn1 = 32'd6073
; 
32'd136617: dataIn1 = 32'd6081
; 
32'd136618: dataIn1 = 32'd6094
; 
32'd136619: dataIn1 = 32'd6704
; 
32'd136620: dataIn1 = 32'd6707
; 
32'd136621: dataIn1 = 32'd2694
; 
32'd136622: dataIn1 = 32'd7076
; 
32'd136623: dataIn1 = 32'd7077
; 
32'd136624: dataIn1 = 32'd7084
; 
32'd136625: dataIn1 = 32'd7103
; 
32'd136626: dataIn1 = 32'd7184
; 
32'd136627: dataIn1 = 32'd7185
; 
32'd136628: dataIn1 = 32'd2695
; 
32'd136629: dataIn1 = 32'd7131
; 
32'd136630: dataIn1 = 32'd7132
; 
32'd136631: dataIn1 = 32'd7138
; 
32'd136632: dataIn1 = 32'd7162
; 
32'd136633: dataIn1 = 32'd9361
; 
32'd136634: dataIn1 = 32'd9362
; 
32'd136635: dataIn1 = 32'd2696
; 
32'd136636: dataIn1 = 32'd7176
; 
32'd136637: dataIn1 = 32'd7177
; 
32'd136638: dataIn1 = 32'd7198
; 
32'd136639: dataIn1 = 32'd7219
; 
32'd136640: dataIn1 = 32'd8883
; 
32'd136641: dataIn1 = 32'd8884
; 
32'd136642: dataIn1 = 32'd2697
; 
32'd136643: dataIn1 = 32'd5133
; 
32'd136644: dataIn1 = 32'd5139
; 
32'd136645: dataIn1 = 32'd6149
; 
32'd136646: dataIn1 = 32'd6150
; 
32'd136647: dataIn1 = 32'd6157
; 
32'd136648: dataIn1 = 32'd6158
; 
32'd136649: dataIn1 = 32'd7272
; 
32'd136650: dataIn1 = 32'd2698
; 
32'd136651: dataIn1 = 32'd2701
; 
32'd136652: dataIn1 = 32'd2702
; 
32'd136653: dataIn1 = 32'd5131
; 
32'd136654: dataIn1 = 32'd5133
; 
32'd136655: dataIn1 = 32'd5135
; 
32'd136656: dataIn1 = 32'd5138
; 
32'd136657: dataIn1 = 32'd2699
; 
32'd136658: dataIn1 = 32'd6142
; 
32'd136659: dataIn1 = 32'd6144
; 
32'd136660: dataIn1 = 32'd7245
; 
32'd136661: dataIn1 = 32'd7246
; 
32'd136662: dataIn1 = 32'd7310
; 
32'd136663: dataIn1 = 32'd7311
; 
32'd136664: dataIn1 = 32'd2700
; 
32'd136665: dataIn1 = 32'd5144
; 
32'd136666: dataIn1 = 32'd5270
; 
32'd136667: dataIn1 = 32'd9668
; 
32'd136668: dataIn1 = 32'd9669
; 
32'd136669: dataIn1 = 32'd9670
; 
32'd136670: dataIn1 = 32'd9671
; 
32'd136671: dataIn1 = 32'd10120
; 
32'd136672: dataIn1 = 32'd16
; 
32'd136673: dataIn1 = 32'd1122
; 
32'd136674: dataIn1 = 32'd2698
; 
32'd136675: dataIn1 = 32'd2701
; 
32'd136676: dataIn1 = 32'd2702
; 
32'd136677: dataIn1 = 32'd2740
; 
32'd136678: dataIn1 = 32'd2742
; 
32'd136679: dataIn1 = 32'd5138
; 
32'd136680: dataIn1 = 32'd16
; 
32'd136681: dataIn1 = 32'd1121
; 
32'd136682: dataIn1 = 32'd2698
; 
32'd136683: dataIn1 = 32'd2701
; 
32'd136684: dataIn1 = 32'd2702
; 
32'd136685: dataIn1 = 32'd2744
; 
32'd136686: dataIn1 = 32'd2746
; 
32'd136687: dataIn1 = 32'd5135
; 
32'd136688: dataIn1 = 32'd2703
; 
32'd136689: dataIn1 = 32'd7302
; 
32'd136690: dataIn1 = 32'd7303
; 
32'd136691: dataIn1 = 32'd7316
; 
32'd136692: dataIn1 = 32'd7351
; 
32'd136693: dataIn1 = 32'd8940
; 
32'd136694: dataIn1 = 32'd8941
; 
32'd136695: dataIn1 = 32'd2704
; 
32'd136696: dataIn1 = 32'd7368
; 
32'd136697: dataIn1 = 32'd7369
; 
32'd136698: dataIn1 = 32'd7398
; 
32'd136699: dataIn1 = 32'd7415
; 
32'd136700: dataIn1 = 32'd7431
; 
32'd136701: dataIn1 = 32'd7432
; 
32'd136702: dataIn1 = 32'd2705
; 
32'd136703: dataIn1 = 32'd6744
; 
32'd136704: dataIn1 = 32'd6745
; 
32'd136705: dataIn1 = 32'd9235
; 
32'd136706: dataIn1 = 32'd9236
; 
32'd136707: dataIn1 = 32'd9287
; 
32'd136708: dataIn1 = 32'd9290
; 
32'd136709: dataIn1 = 32'd2706
; 
32'd136710: dataIn1 = 32'd7377
; 
32'd136711: dataIn1 = 32'd7378
; 
32'd136712: dataIn1 = 32'd7385
; 
32'd136713: dataIn1 = 32'd7411
; 
32'd136714: dataIn1 = 32'd7540
; 
32'd136715: dataIn1 = 32'd7541
; 
32'd136716: dataIn1 = 32'd2707
; 
32'd136717: dataIn1 = 32'd7439
; 
32'd136718: dataIn1 = 32'd7440
; 
32'd136719: dataIn1 = 32'd7466
; 
32'd136720: dataIn1 = 32'd7511
; 
32'd136721: dataIn1 = 32'd8948
; 
32'd136722: dataIn1 = 32'd8949
; 
32'd136723: dataIn1 = 32'd2708
; 
32'd136724: dataIn1 = 32'd7532
; 
32'd136725: dataIn1 = 32'd7533
; 
32'd136726: dataIn1 = 32'd7554
; 
32'd136727: dataIn1 = 32'd7599
; 
32'd136728: dataIn1 = 32'd8989
; 
32'd136729: dataIn1 = 32'd8990
; 
32'd136730: dataIn1 = 32'd2709
; 
32'd136731: dataIn1 = 32'd7619
; 
32'd136732: dataIn1 = 32'd7620
; 
32'd136733: dataIn1 = 32'd7649
; 
32'd136734: dataIn1 = 32'd7666
; 
32'd136735: dataIn1 = 32'd7682
; 
32'd136736: dataIn1 = 32'd7683
; 
32'd136737: dataIn1 = 32'd2710
; 
32'd136738: dataIn1 = 32'd6754
; 
32'd136739: dataIn1 = 32'd6755
; 
32'd136740: dataIn1 = 32'd9240
; 
32'd136741: dataIn1 = 32'd9241
; 
32'd136742: dataIn1 = 32'd9293
; 
32'd136743: dataIn1 = 32'd9296
; 
32'd136744: dataIn1 = 32'd2711
; 
32'd136745: dataIn1 = 32'd7628
; 
32'd136746: dataIn1 = 32'd7629
; 
32'd136747: dataIn1 = 32'd7636
; 
32'd136748: dataIn1 = 32'd7662
; 
32'd136749: dataIn1 = 32'd7793
; 
32'd136750: dataIn1 = 32'd7794
; 
32'd136751: dataIn1 = 32'd2712
; 
32'd136752: dataIn1 = 32'd7690
; 
32'd136753: dataIn1 = 32'd7691
; 
32'd136754: dataIn1 = 32'd7719
; 
32'd136755: dataIn1 = 32'd7764
; 
32'd136756: dataIn1 = 32'd8997
; 
32'd136757: dataIn1 = 32'd8998
; 
32'd136758: dataIn1 = 32'd2713
; 
32'd136759: dataIn1 = 32'd7785
; 
32'd136760: dataIn1 = 32'd7786
; 
32'd136761: dataIn1 = 32'd7807
; 
32'd136762: dataIn1 = 32'd7852
; 
32'd136763: dataIn1 = 32'd9041
; 
32'd136764: dataIn1 = 32'd9042
; 
32'd136765: dataIn1 = 32'd2714
; 
32'd136766: dataIn1 = 32'd7872
; 
32'd136767: dataIn1 = 32'd7873
; 
32'd136768: dataIn1 = 32'd7902
; 
32'd136769: dataIn1 = 32'd7919
; 
32'd136770: dataIn1 = 32'd7935
; 
32'd136771: dataIn1 = 32'd7936
; 
32'd136772: dataIn1 = 32'd2715
; 
32'd136773: dataIn1 = 32'd6314
; 
32'd136774: dataIn1 = 32'd6315
; 
32'd136775: dataIn1 = 32'd6321
; 
32'd136776: dataIn1 = 32'd6335
; 
32'd136777: dataIn1 = 32'd6708
; 
32'd136778: dataIn1 = 32'd6711
; 
32'd136779: dataIn1 = 32'd2716
; 
32'd136780: dataIn1 = 32'd7881
; 
32'd136781: dataIn1 = 32'd7882
; 
32'd136782: dataIn1 = 32'd7889
; 
32'd136783: dataIn1 = 32'd7915
; 
32'd136784: dataIn1 = 32'd8046
; 
32'd136785: dataIn1 = 32'd8047
; 
32'd136786: dataIn1 = 32'd2717
; 
32'd136787: dataIn1 = 32'd7943
; 
32'd136788: dataIn1 = 32'd7944
; 
32'd136789: dataIn1 = 32'd7972
; 
32'd136790: dataIn1 = 32'd8017
; 
32'd136791: dataIn1 = 32'd9049
; 
32'd136792: dataIn1 = 32'd9050
; 
32'd136793: dataIn1 = 32'd2718
; 
32'd136794: dataIn1 = 32'd8038
; 
32'd136795: dataIn1 = 32'd8039
; 
32'd136796: dataIn1 = 32'd8060
; 
32'd136797: dataIn1 = 32'd8105
; 
32'd136798: dataIn1 = 32'd9092
; 
32'd136799: dataIn1 = 32'd9093
; 
32'd136800: dataIn1 = 32'd2719
; 
32'd136801: dataIn1 = 32'd8125
; 
32'd136802: dataIn1 = 32'd8126
; 
32'd136803: dataIn1 = 32'd8155
; 
32'd136804: dataIn1 = 32'd8172
; 
32'd136805: dataIn1 = 32'd8188
; 
32'd136806: dataIn1 = 32'd8189
; 
32'd136807: dataIn1 = 32'd2720
; 
32'd136808: dataIn1 = 32'd6388
; 
32'd136809: dataIn1 = 32'd6389
; 
32'd136810: dataIn1 = 32'd6397
; 
32'd136811: dataIn1 = 32'd6409
; 
32'd136812: dataIn1 = 32'd6716
; 
32'd136813: dataIn1 = 32'd9776
; 
32'd136814: dataIn1 = 32'd2721
; 
32'd136815: dataIn1 = 32'd8134
; 
32'd136816: dataIn1 = 32'd8135
; 
32'd136817: dataIn1 = 32'd8142
; 
32'd136818: dataIn1 = 32'd8168
; 
32'd136819: dataIn1 = 32'd8299
; 
32'd136820: dataIn1 = 32'd8300
; 
32'd136821: dataIn1 = 32'd2722
; 
32'd136822: dataIn1 = 32'd8196
; 
32'd136823: dataIn1 = 32'd8197
; 
32'd136824: dataIn1 = 32'd8225
; 
32'd136825: dataIn1 = 32'd8270
; 
32'd136826: dataIn1 = 32'd9100
; 
32'd136827: dataIn1 = 32'd9101
; 
32'd136828: dataIn1 = 32'd2723
; 
32'd136829: dataIn1 = 32'd8291
; 
32'd136830: dataIn1 = 32'd8292
; 
32'd136831: dataIn1 = 32'd8313
; 
32'd136832: dataIn1 = 32'd8357
; 
32'd136833: dataIn1 = 32'd9144
; 
32'd136834: dataIn1 = 32'd9145
; 
32'd136835: dataIn1 = 32'd2724
; 
32'd136836: dataIn1 = 32'd8377
; 
32'd136837: dataIn1 = 32'd8378
; 
32'd136838: dataIn1 = 32'd8407
; 
32'd136839: dataIn1 = 32'd8424
; 
32'd136840: dataIn1 = 32'd8440
; 
32'd136841: dataIn1 = 32'd8441
; 
32'd136842: dataIn1 = 32'd2725
; 
32'd136843: dataIn1 = 32'd6766
; 
32'd136844: dataIn1 = 32'd6767
; 
32'd136845: dataIn1 = 32'd9246
; 
32'd136846: dataIn1 = 32'd9247
; 
32'd136847: dataIn1 = 32'd9299
; 
32'd136848: dataIn1 = 32'd9302
; 
32'd136849: dataIn1 = 32'd2726
; 
32'd136850: dataIn1 = 32'd8386
; 
32'd136851: dataIn1 = 32'd8387
; 
32'd136852: dataIn1 = 32'd8394
; 
32'd136853: dataIn1 = 32'd8420
; 
32'd136854: dataIn1 = 32'd8551
; 
32'd136855: dataIn1 = 32'd8552
; 
32'd136856: dataIn1 = 32'd2727
; 
32'd136857: dataIn1 = 32'd8448
; 
32'd136858: dataIn1 = 32'd8449
; 
32'd136859: dataIn1 = 32'd8477
; 
32'd136860: dataIn1 = 32'd8522
; 
32'd136861: dataIn1 = 32'd9152
; 
32'd136862: dataIn1 = 32'd9153
; 
32'd136863: dataIn1 = 32'd2728
; 
32'd136864: dataIn1 = 32'd8543
; 
32'd136865: dataIn1 = 32'd8544
; 
32'd136866: dataIn1 = 32'd8565
; 
32'd136867: dataIn1 = 32'd8610
; 
32'd136868: dataIn1 = 32'd9194
; 
32'd136869: dataIn1 = 32'd9195
; 
32'd136870: dataIn1 = 32'd2729
; 
32'd136871: dataIn1 = 32'd8630
; 
32'd136872: dataIn1 = 32'd8631
; 
32'd136873: dataIn1 = 32'd8660
; 
32'd136874: dataIn1 = 32'd8677
; 
32'd136875: dataIn1 = 32'd8693
; 
32'd136876: dataIn1 = 32'd8694
; 
32'd136877: dataIn1 = 32'd2730
; 
32'd136878: dataIn1 = 32'd6776
; 
32'd136879: dataIn1 = 32'd6777
; 
32'd136880: dataIn1 = 32'd9252
; 
32'd136881: dataIn1 = 32'd9253
; 
32'd136882: dataIn1 = 32'd9305
; 
32'd136883: dataIn1 = 32'd9308
; 
32'd136884: dataIn1 = 32'd2731
; 
32'd136885: dataIn1 = 32'd8639
; 
32'd136886: dataIn1 = 32'd8640
; 
32'd136887: dataIn1 = 32'd8647
; 
32'd136888: dataIn1 = 32'd8673
; 
32'd136889: dataIn1 = 32'd8804
; 
32'd136890: dataIn1 = 32'd8805
; 
32'd136891: dataIn1 = 32'd2732
; 
32'd136892: dataIn1 = 32'd8701
; 
32'd136893: dataIn1 = 32'd8702
; 
32'd136894: dataIn1 = 32'd8730
; 
32'd136895: dataIn1 = 32'd8775
; 
32'd136896: dataIn1 = 32'd9202
; 
32'd136897: dataIn1 = 32'd9203
; 
32'd136898: dataIn1 = 32'd2733
; 
32'd136899: dataIn1 = 32'd8796
; 
32'd136900: dataIn1 = 32'd8797
; 
32'd136901: dataIn1 = 32'd8862
; 
32'd136902: dataIn1 = 32'd9276
; 
32'd136903: dataIn1 = 32'd9404
; 
32'd136904: dataIn1 = 32'd9405
; 
32'd136905: dataIn1 = 32'd2734
; 
32'd136906: dataIn1 = 32'd6576
; 
32'd136907: dataIn1 = 32'd6577
; 
32'd136908: dataIn1 = 32'd6588
; 
32'd136909: dataIn1 = 32'd6593
; 
32'd136910: dataIn1 = 32'd6718
; 
32'd136911: dataIn1 = 32'd6720
; 
32'd136912: dataIn1 = 32'd1135
; 
32'd136913: dataIn1 = 32'd2735
; 
32'd136914: dataIn1 = 32'd5513
; 
32'd136915: dataIn1 = 32'd6719
; 
32'd136916: dataIn1 = 32'd6720
; 
32'd136917: dataIn1 = 32'd6733
; 
32'd136918: dataIn1 = 32'd6741
; 
32'd136919: dataIn1 = 32'd1135
; 
32'd136920: dataIn1 = 32'd2736
; 
32'd136921: dataIn1 = 32'd2737
; 
32'd136922: dataIn1 = 32'd6717
; 
32'd136923: dataIn1 = 32'd6718
; 
32'd136924: dataIn1 = 32'd6741
; 
32'd136925: dataIn1 = 32'd6742
; 
32'd136926: dataIn1 = 32'd15
; 
32'd136927: dataIn1 = 32'd1135
; 
32'd136928: dataIn1 = 32'd2323
; 
32'd136929: dataIn1 = 32'd2736
; 
32'd136930: dataIn1 = 32'd2737
; 
32'd136931: dataIn1 = 32'd3433
; 
32'd136932: dataIn1 = 32'd6742
; 
32'd136933: dataIn1 = 32'd2738
; 
32'd136934: dataIn1 = 32'd2740
; 
32'd136935: dataIn1 = 32'd5270
; 
32'd136936: dataIn1 = 32'd5271
; 
32'd136937: dataIn1 = 32'd5272
; 
32'd136938: dataIn1 = 32'd5273
; 
32'd136939: dataIn1 = 32'd5634
; 
32'd136940: dataIn1 = 32'd1136
; 
32'd136941: dataIn1 = 32'd2739
; 
32'd136942: dataIn1 = 32'd2740
; 
32'd136943: dataIn1 = 32'd2741
; 
32'd136944: dataIn1 = 32'd5633
; 
32'd136945: dataIn1 = 32'd5634
; 
32'd136946: dataIn1 = 32'd6691
; 
32'd136947: dataIn1 = 32'd1122
; 
32'd136948: dataIn1 = 32'd1136
; 
32'd136949: dataIn1 = 32'd2701
; 
32'd136950: dataIn1 = 32'd2738
; 
32'd136951: dataIn1 = 32'd2739
; 
32'd136952: dataIn1 = 32'd2740
; 
32'd136953: dataIn1 = 32'd2742
; 
32'd136954: dataIn1 = 32'd5272
; 
32'd136955: dataIn1 = 32'd5634
; 
32'd136956: dataIn1 = 32'd15
; 
32'd136957: dataIn1 = 32'd1136
; 
32'd136958: dataIn1 = 32'd2324
; 
32'd136959: dataIn1 = 32'd2739
; 
32'd136960: dataIn1 = 32'd2741
; 
32'd136961: dataIn1 = 32'd3436
; 
32'd136962: dataIn1 = 32'd6691
; 
32'd136963: dataIn1 = 32'd16
; 
32'd136964: dataIn1 = 32'd1136
; 
32'd136965: dataIn1 = 32'd2701
; 
32'd136966: dataIn1 = 32'd2740
; 
32'd136967: dataIn1 = 32'd2742
; 
32'd136968: dataIn1 = 32'd3435
; 
32'd136969: dataIn1 = 32'd2743
; 
32'd136970: dataIn1 = 32'd2744
; 
32'd136971: dataIn1 = 32'd5278
; 
32'd136972: dataIn1 = 32'd9277
; 
32'd136973: dataIn1 = 32'd9278
; 
32'd136974: dataIn1 = 32'd9321
; 
32'd136975: dataIn1 = 32'd9338
; 
32'd136976: dataIn1 = 32'd1121
; 
32'd136977: dataIn1 = 32'd1137
; 
32'd136978: dataIn1 = 32'd2702
; 
32'd136979: dataIn1 = 32'd2743
; 
32'd136980: dataIn1 = 32'd2744
; 
32'd136981: dataIn1 = 32'd2745
; 
32'd136982: dataIn1 = 32'd2746
; 
32'd136983: dataIn1 = 32'd5278
; 
32'd136984: dataIn1 = 32'd9338
; 
32'd136985: dataIn1 = 32'd1137
; 
32'd136986: dataIn1 = 32'd2744
; 
32'd136987: dataIn1 = 32'd2745
; 
32'd136988: dataIn1 = 32'd5515
; 
32'd136989: dataIn1 = 32'd9337
; 
32'd136990: dataIn1 = 32'd9338
; 
32'd136991: dataIn1 = 32'd9339
; 
32'd136992: dataIn1 = 32'd16
; 
32'd136993: dataIn1 = 32'd1137
; 
32'd136994: dataIn1 = 32'd2702
; 
32'd136995: dataIn1 = 32'd2744
; 
32'd136996: dataIn1 = 32'd2746
; 
32'd136997: dataIn1 = 32'd3437
; 
32'd136998: dataIn1 = 32'd2747
; 
32'd136999: dataIn1 = 32'd6786
; 
32'd137000: dataIn1 = 32'd6787
; 
32'd137001: dataIn1 = 32'd9258
; 
32'd137002: dataIn1 = 32'd9259
; 
32'd137003: dataIn1 = 32'd9292
; 
32'd137004: dataIn1 = 32'd9298
; 
32'd137005: dataIn1 = 32'd17
; 
32'd137006: dataIn1 = 32'd28
; 
32'd137007: dataIn1 = 32'd1138
; 
32'd137008: dataIn1 = 32'd2108
; 
32'd137009: dataIn1 = 32'd2138
; 
32'd137010: dataIn1 = 32'd2748
; 
32'd137011: dataIn1 = 32'd3419
; 
32'd137012: dataIn1 = 32'd5514
; 
32'd137013: dataIn1 = 32'd2749
; 
32'd137014: dataIn1 = 32'd6626
; 
32'd137015: dataIn1 = 32'd6627
; 
32'd137016: dataIn1 = 32'd6636
; 
32'd137017: dataIn1 = 32'd6722
; 
32'd137018: dataIn1 = 32'd9036
; 
32'd137019: dataIn1 = 32'd9282
; 
32'd137020: dataIn1 = 32'd2750
; 
32'd137021: dataIn1 = 32'd6644
; 
32'd137022: dataIn1 = 32'd6645
; 
32'd137023: dataIn1 = 32'd6654
; 
32'd137024: dataIn1 = 32'd6657
; 
32'd137025: dataIn1 = 32'd6724
; 
32'd137026: dataIn1 = 32'd6727
; 
32'd137027: dataIn1 = 32'd2751
; 
32'd137028: dataIn1 = 32'd6664
; 
32'd137029: dataIn1 = 32'd6665
; 
32'd137030: dataIn1 = 32'd6677
; 
32'd137031: dataIn1 = 32'd6729
; 
32'd137032: dataIn1 = 32'd9139
; 
32'd137033: dataIn1 = 32'd9284
; 
32'd137034: dataIn1 = 32'd2752
; 
32'd137035: dataIn1 = 32'd6796
; 
32'd137036: dataIn1 = 32'd6797
; 
32'd137037: dataIn1 = 32'd9260
; 
32'd137038: dataIn1 = 32'd9261
; 
32'd137039: dataIn1 = 32'd9304
; 
32'd137040: dataIn1 = 32'd9310
; 
32'd137041: dataIn1 = 32'd541
; 
32'd137042: dataIn1 = 32'd542
; 
32'd137043: dataIn1 = 32'd1244
; 
32'd137044: dataIn1 = 32'd1248
; 
32'd137045: dataIn1 = 32'd2481
; 
32'd137046: dataIn1 = 32'd2753
; 
32'd137047: dataIn1 = 32'd2754
; 
32'd137048: dataIn1 = 32'd541
; 
32'd137049: dataIn1 = 32'd543
; 
32'd137050: dataIn1 = 32'd1243
; 
32'd137051: dataIn1 = 32'd1248
; 
32'd137052: dataIn1 = 32'd2753
; 
32'd137053: dataIn1 = 32'd2754
; 
32'd137054: dataIn1 = 32'd3438
; 
32'd137055: dataIn1 = 32'd547
; 
32'd137056: dataIn1 = 32'd548
; 
32'd137057: dataIn1 = 32'd1260
; 
32'd137058: dataIn1 = 32'd2480
; 
32'd137059: dataIn1 = 32'd2755
; 
32'd137060: dataIn1 = 32'd10250
; 
32'd137061: dataIn1 = 32'd10269
; 
32'd137062: dataIn1 = 32'd266
; 
32'd137063: dataIn1 = 32'd548
; 
32'd137064: dataIn1 = 32'd549
; 
32'd137065: dataIn1 = 32'd1262
; 
32'd137066: dataIn1 = 32'd2482
; 
32'd137067: dataIn1 = 32'd2756
; 
32'd137068: dataIn1 = 32'd285
; 
32'd137069: dataIn1 = 32'd583
; 
32'd137070: dataIn1 = 32'd2484
; 
32'd137071: dataIn1 = 32'd2757
; 
32'd137072: dataIn1 = 32'd2766
; 
32'd137073: dataIn1 = 32'd2769
; 
32'd137074: dataIn1 = 32'd10985
; 
32'd137075: dataIn1 = 32'd768
; 
32'd137076: dataIn1 = 32'd783
; 
32'd137077: dataIn1 = 32'd1462
; 
32'd137078: dataIn1 = 32'd1490
; 
32'd137079: dataIn1 = 32'd2498
; 
32'd137080: dataIn1 = 32'd2758
; 
32'd137081: dataIn1 = 32'd3439
; 
32'd137082: dataIn1 = 32'd798
; 
32'd137083: dataIn1 = 32'd800
; 
32'd137084: dataIn1 = 32'd1506
; 
32'd137085: dataIn1 = 32'd1872
; 
32'd137086: dataIn1 = 32'd2512
; 
32'd137087: dataIn1 = 32'd2759
; 
32'd137088: dataIn1 = 32'd3040
; 
32'd137089: dataIn1 = 32'd806
; 
32'd137090: dataIn1 = 32'd1514
; 
32'd137091: dataIn1 = 32'd1518
; 
32'd137092: dataIn1 = 32'd2522
; 
32'd137093: dataIn1 = 32'd2760
; 
32'd137094: dataIn1 = 32'd3440
; 
32'd137095: dataIn1 = 32'd10976
; 
32'd137096: dataIn1 = 32'd1723
; 
32'd137097: dataIn1 = 32'd1724
; 
32'd137098: dataIn1 = 32'd2761
; 
32'd137099: dataIn1 = 32'd2762
; 
32'd137100: dataIn1 = 32'd2763
; 
32'd137101: dataIn1 = 32'd2764
; 
32'd137102: dataIn1 = 32'd2765
; 
32'd137103: dataIn1 = 32'd1724
; 
32'd137104: dataIn1 = 32'd2761
; 
32'd137105: dataIn1 = 32'd2762
; 
32'd137106: dataIn1 = 32'd2763
; 
32'd137107: dataIn1 = 32'd3045
; 
32'd137108: dataIn1 = 32'd10991
; 
32'd137109: dataIn1 = 32'd10992
; 
32'd137110: dataIn1 = 32'd1723
; 
32'd137111: dataIn1 = 32'd2761
; 
32'd137112: dataIn1 = 32'd2762
; 
32'd137113: dataIn1 = 32'd2763
; 
32'd137114: dataIn1 = 32'd3053
; 
32'd137115: dataIn1 = 32'd10990
; 
32'd137116: dataIn1 = 32'd10991
; 
32'd137117: dataIn1 = 32'd279
; 
32'd137118: dataIn1 = 32'd1724
; 
32'd137119: dataIn1 = 32'd2761
; 
32'd137120: dataIn1 = 32'd2764
; 
32'd137121: dataIn1 = 32'd2765
; 
32'd137122: dataIn1 = 32'd3041
; 
32'd137123: dataIn1 = 32'd3044
; 
32'd137124: dataIn1 = 32'd279
; 
32'd137125: dataIn1 = 32'd1723
; 
32'd137126: dataIn1 = 32'd2761
; 
32'd137127: dataIn1 = 32'd2764
; 
32'd137128: dataIn1 = 32'd2765
; 
32'd137129: dataIn1 = 32'd3048
; 
32'd137130: dataIn1 = 32'd3051
; 
32'd137131: dataIn1 = 32'd583
; 
32'd137132: dataIn1 = 32'd1726
; 
32'd137133: dataIn1 = 32'd2757
; 
32'd137134: dataIn1 = 32'd2766
; 
32'd137135: dataIn1 = 32'd2767
; 
32'd137136: dataIn1 = 32'd2768
; 
32'd137137: dataIn1 = 32'd2769
; 
32'd137138: dataIn1 = 32'd1725
; 
32'd137139: dataIn1 = 32'd1726
; 
32'd137140: dataIn1 = 32'd2766
; 
32'd137141: dataIn1 = 32'd2767
; 
32'd137142: dataIn1 = 32'd2768
; 
32'd137143: dataIn1 = 32'd2770
; 
32'd137144: dataIn1 = 32'd2771
; 
32'd137145: dataIn1 = 32'd583
; 
32'd137146: dataIn1 = 32'd1299
; 
32'd137147: dataIn1 = 32'd1725
; 
32'd137148: dataIn1 = 32'd2766
; 
32'd137149: dataIn1 = 32'd2767
; 
32'd137150: dataIn1 = 32'd2768
; 
32'd137151: dataIn1 = 32'd3054
; 
32'd137152: dataIn1 = 32'd285
; 
32'd137153: dataIn1 = 32'd1726
; 
32'd137154: dataIn1 = 32'd2757
; 
32'd137155: dataIn1 = 32'd2766
; 
32'd137156: dataIn1 = 32'd2769
; 
32'd137157: dataIn1 = 32'd3868
; 
32'd137158: dataIn1 = 32'd5304
; 
32'd137159: dataIn1 = 32'd154
; 
32'd137160: dataIn1 = 32'd1726
; 
32'd137161: dataIn1 = 32'd2767
; 
32'd137162: dataIn1 = 32'd2770
; 
32'd137163: dataIn1 = 32'd2771
; 
32'd137164: dataIn1 = 32'd3869
; 
32'd137165: dataIn1 = 32'd3933
; 
32'd137166: dataIn1 = 32'd154
; 
32'd137167: dataIn1 = 32'd1725
; 
32'd137168: dataIn1 = 32'd2767
; 
32'd137169: dataIn1 = 32'd2770
; 
32'd137170: dataIn1 = 32'd2771
; 
32'd137171: dataIn1 = 32'd3049
; 
32'd137172: dataIn1 = 32'd3052
; 
32'd137173: dataIn1 = 32'd1728
; 
32'd137174: dataIn1 = 32'd2772
; 
32'd137175: dataIn1 = 32'd2773
; 
32'd137176: dataIn1 = 32'd2774
; 
32'd137177: dataIn1 = 32'd3058
; 
32'd137178: dataIn1 = 32'd10998
; 
32'd137179: dataIn1 = 32'd10999
; 
32'd137180: dataIn1 = 32'd1727
; 
32'd137181: dataIn1 = 32'd1728
; 
32'd137182: dataIn1 = 32'd2772
; 
32'd137183: dataIn1 = 32'd2773
; 
32'd137184: dataIn1 = 32'd2774
; 
32'd137185: dataIn1 = 32'd2775
; 
32'd137186: dataIn1 = 32'd2776
; 
32'd137187: dataIn1 = 32'd1727
; 
32'd137188: dataIn1 = 32'd2772
; 
32'd137189: dataIn1 = 32'd2773
; 
32'd137190: dataIn1 = 32'd2774
; 
32'd137191: dataIn1 = 32'd3068
; 
32'd137192: dataIn1 = 32'd10999
; 
32'd137193: dataIn1 = 32'd11000
; 
32'd137194: dataIn1 = 32'd286
; 
32'd137195: dataIn1 = 32'd1728
; 
32'd137196: dataIn1 = 32'd2773
; 
32'd137197: dataIn1 = 32'd2775
; 
32'd137198: dataIn1 = 32'd2776
; 
32'd137199: dataIn1 = 32'd3056
; 
32'd137200: dataIn1 = 32'd3060
; 
32'd137201: dataIn1 = 32'd286
; 
32'd137202: dataIn1 = 32'd1727
; 
32'd137203: dataIn1 = 32'd2773
; 
32'd137204: dataIn1 = 32'd2775
; 
32'd137205: dataIn1 = 32'd2776
; 
32'd137206: dataIn1 = 32'd3063
; 
32'd137207: dataIn1 = 32'd3066
; 
32'd137208: dataIn1 = 32'd1730
; 
32'd137209: dataIn1 = 32'd2777
; 
32'd137210: dataIn1 = 32'd2778
; 
32'd137211: dataIn1 = 32'd2779
; 
32'd137212: dataIn1 = 32'd3059
; 
32'd137213: dataIn1 = 32'd10995
; 
32'd137214: dataIn1 = 32'd10996
; 
32'd137215: dataIn1 = 32'd1729
; 
32'd137216: dataIn1 = 32'd2777
; 
32'd137217: dataIn1 = 32'd2778
; 
32'd137218: dataIn1 = 32'd2779
; 
32'd137219: dataIn1 = 32'd3046
; 
32'd137220: dataIn1 = 32'd10994
; 
32'd137221: dataIn1 = 32'd10995
; 
32'd137222: dataIn1 = 32'd1729
; 
32'd137223: dataIn1 = 32'd1730
; 
32'd137224: dataIn1 = 32'd2777
; 
32'd137225: dataIn1 = 32'd2778
; 
32'd137226: dataIn1 = 32'd2779
; 
32'd137227: dataIn1 = 32'd2780
; 
32'd137228: dataIn1 = 32'd2781
; 
32'd137229: dataIn1 = 32'd155
; 
32'd137230: dataIn1 = 32'd1730
; 
32'd137231: dataIn1 = 32'd2779
; 
32'd137232: dataIn1 = 32'd2780
; 
32'd137233: dataIn1 = 32'd2781
; 
32'd137234: dataIn1 = 32'd3057
; 
32'd137235: dataIn1 = 32'd3061
; 
32'd137236: dataIn1 = 32'd155
; 
32'd137237: dataIn1 = 32'd1729
; 
32'd137238: dataIn1 = 32'd2779
; 
32'd137239: dataIn1 = 32'd2780
; 
32'd137240: dataIn1 = 32'd2781
; 
32'd137241: dataIn1 = 32'd3043
; 
32'd137242: dataIn1 = 32'd3047
; 
32'd137243: dataIn1 = 32'd1731
; 
32'd137244: dataIn1 = 32'd1732
; 
32'd137245: dataIn1 = 32'd2782
; 
32'd137246: dataIn1 = 32'd2783
; 
32'd137247: dataIn1 = 32'd2784
; 
32'd137248: dataIn1 = 32'd2785
; 
32'd137249: dataIn1 = 32'd2786
; 
32'd137250: dataIn1 = 32'd1732
; 
32'd137251: dataIn1 = 32'd2782
; 
32'd137252: dataIn1 = 32'd2783
; 
32'd137253: dataIn1 = 32'd2784
; 
32'd137254: dataIn1 = 32'd3074
; 
32'd137255: dataIn1 = 32'd11003
; 
32'd137256: dataIn1 = 32'd11004
; 
32'd137257: dataIn1 = 32'd1731
; 
32'd137258: dataIn1 = 32'd2782
; 
32'd137259: dataIn1 = 32'd2783
; 
32'd137260: dataIn1 = 32'd2784
; 
32'd137261: dataIn1 = 32'd3067
; 
32'd137262: dataIn1 = 32'd11002
; 
32'd137263: dataIn1 = 32'd11003
; 
32'd137264: dataIn1 = 32'd157
; 
32'd137265: dataIn1 = 32'd1732
; 
32'd137266: dataIn1 = 32'd2782
; 
32'd137267: dataIn1 = 32'd2785
; 
32'd137268: dataIn1 = 32'd2786
; 
32'd137269: dataIn1 = 32'd3069
; 
32'd137270: dataIn1 = 32'd3072
; 
32'd137271: dataIn1 = 32'd157
; 
32'd137272: dataIn1 = 32'd1731
; 
32'd137273: dataIn1 = 32'd2782
; 
32'd137274: dataIn1 = 32'd2785
; 
32'd137275: dataIn1 = 32'd2786
; 
32'd137276: dataIn1 = 32'd3062
; 
32'd137277: dataIn1 = 32'd3065
; 
32'd137278: dataIn1 = 32'd1734
; 
32'd137279: dataIn1 = 32'd2787
; 
32'd137280: dataIn1 = 32'd2788
; 
32'd137281: dataIn1 = 32'd2789
; 
32'd137282: dataIn1 = 32'd3079
; 
32'd137283: dataIn1 = 32'd11007
; 
32'd137284: dataIn1 = 32'd11008
; 
32'd137285: dataIn1 = 32'd1733
; 
32'd137286: dataIn1 = 32'd1734
; 
32'd137287: dataIn1 = 32'd2787
; 
32'd137288: dataIn1 = 32'd2788
; 
32'd137289: dataIn1 = 32'd2789
; 
32'd137290: dataIn1 = 32'd2790
; 
32'd137291: dataIn1 = 32'd2791
; 
32'd137292: dataIn1 = 32'd1733
; 
32'd137293: dataIn1 = 32'd2787
; 
32'd137294: dataIn1 = 32'd2788
; 
32'd137295: dataIn1 = 32'd2789
; 
32'd137296: dataIn1 = 32'd3075
; 
32'd137297: dataIn1 = 32'd11006
; 
32'd137298: dataIn1 = 32'd11007
; 
32'd137299: dataIn1 = 32'd293
; 
32'd137300: dataIn1 = 32'd1734
; 
32'd137301: dataIn1 = 32'd2788
; 
32'd137302: dataIn1 = 32'd2790
; 
32'd137303: dataIn1 = 32'd2791
; 
32'd137304: dataIn1 = 32'd3077
; 
32'd137305: dataIn1 = 32'd3081
; 
32'd137306: dataIn1 = 32'd293
; 
32'd137307: dataIn1 = 32'd1733
; 
32'd137308: dataIn1 = 32'd2788
; 
32'd137309: dataIn1 = 32'd2790
; 
32'd137310: dataIn1 = 32'd2791
; 
32'd137311: dataIn1 = 32'd3070
; 
32'd137312: dataIn1 = 32'd3073
; 
32'd137313: dataIn1 = 32'd1735
; 
32'd137314: dataIn1 = 32'd1736
; 
32'd137315: dataIn1 = 32'd2792
; 
32'd137316: dataIn1 = 32'd2793
; 
32'd137317: dataIn1 = 32'd2794
; 
32'd137318: dataIn1 = 32'd2795
; 
32'd137319: dataIn1 = 32'd2796
; 
32'd137320: dataIn1 = 32'd1736
; 
32'd137321: dataIn1 = 32'd2792
; 
32'd137322: dataIn1 = 32'd2793
; 
32'd137323: dataIn1 = 32'd2794
; 
32'd137324: dataIn1 = 32'd3087
; 
32'd137325: dataIn1 = 32'd11023
; 
32'd137326: dataIn1 = 32'd11024
; 
32'd137327: dataIn1 = 32'd1735
; 
32'd137328: dataIn1 = 32'd2792
; 
32'd137329: dataIn1 = 32'd2793
; 
32'd137330: dataIn1 = 32'd2794
; 
32'd137331: dataIn1 = 32'd3095
; 
32'd137332: dataIn1 = 32'd11022
; 
32'd137333: dataIn1 = 32'd11023
; 
32'd137334: dataIn1 = 32'd295
; 
32'd137335: dataIn1 = 32'd1736
; 
32'd137336: dataIn1 = 32'd2792
; 
32'd137337: dataIn1 = 32'd2795
; 
32'd137338: dataIn1 = 32'd2796
; 
32'd137339: dataIn1 = 32'd3083
; 
32'd137340: dataIn1 = 32'd3086
; 
32'd137341: dataIn1 = 32'd295
; 
32'd137342: dataIn1 = 32'd1735
; 
32'd137343: dataIn1 = 32'd2792
; 
32'd137344: dataIn1 = 32'd2795
; 
32'd137345: dataIn1 = 32'd2796
; 
32'd137346: dataIn1 = 32'd3090
; 
32'd137347: dataIn1 = 32'd3093
; 
32'd137348: dataIn1 = 32'd1738
; 
32'd137349: dataIn1 = 32'd2797
; 
32'd137350: dataIn1 = 32'd2798
; 
32'd137351: dataIn1 = 32'd2799
; 
32'd137352: dataIn1 = 32'd3101
; 
32'd137353: dataIn1 = 32'd11015
; 
32'd137354: dataIn1 = 32'd11016
; 
32'd137355: dataIn1 = 32'd1737
; 
32'd137356: dataIn1 = 32'd2797
; 
32'd137357: dataIn1 = 32'd2798
; 
32'd137358: dataIn1 = 32'd2799
; 
32'd137359: dataIn1 = 32'd3109
; 
32'd137360: dataIn1 = 32'd11014
; 
32'd137361: dataIn1 = 32'd11015
; 
32'd137362: dataIn1 = 32'd1737
; 
32'd137363: dataIn1 = 32'd1738
; 
32'd137364: dataIn1 = 32'd2797
; 
32'd137365: dataIn1 = 32'd2798
; 
32'd137366: dataIn1 = 32'd2799
; 
32'd137367: dataIn1 = 32'd2800
; 
32'd137368: dataIn1 = 32'd2801
; 
32'd137369: dataIn1 = 32'd301
; 
32'd137370: dataIn1 = 32'd1738
; 
32'd137371: dataIn1 = 32'd2799
; 
32'd137372: dataIn1 = 32'd2800
; 
32'd137373: dataIn1 = 32'd2801
; 
32'd137374: dataIn1 = 32'd3099
; 
32'd137375: dataIn1 = 32'd3103
; 
32'd137376: dataIn1 = 32'd301
; 
32'd137377: dataIn1 = 32'd1737
; 
32'd137378: dataIn1 = 32'd2799
; 
32'd137379: dataIn1 = 32'd2800
; 
32'd137380: dataIn1 = 32'd2801
; 
32'd137381: dataIn1 = 32'd3106
; 
32'd137382: dataIn1 = 32'd3110
; 
32'd137383: dataIn1 = 32'd1740
; 
32'd137384: dataIn1 = 32'd2802
; 
32'd137385: dataIn1 = 32'd2803
; 
32'd137386: dataIn1 = 32'd2804
; 
32'd137387: dataIn1 = 32'd3100
; 
32'd137388: dataIn1 = 32'd11018
; 
32'd137389: dataIn1 = 32'd11019
; 
32'd137390: dataIn1 = 32'd1739
; 
32'd137391: dataIn1 = 32'd1740
; 
32'd137392: dataIn1 = 32'd2802
; 
32'd137393: dataIn1 = 32'd2803
; 
32'd137394: dataIn1 = 32'd2804
; 
32'd137395: dataIn1 = 32'd2805
; 
32'd137396: dataIn1 = 32'd2806
; 
32'd137397: dataIn1 = 32'd1739
; 
32'd137398: dataIn1 = 32'd2802
; 
32'd137399: dataIn1 = 32'd2803
; 
32'd137400: dataIn1 = 32'd2804
; 
32'd137401: dataIn1 = 32'd3096
; 
32'd137402: dataIn1 = 32'd11019
; 
32'd137403: dataIn1 = 32'd11020
; 
32'd137404: dataIn1 = 32'd161
; 
32'd137405: dataIn1 = 32'd1740
; 
32'd137406: dataIn1 = 32'd2803
; 
32'd137407: dataIn1 = 32'd2805
; 
32'd137408: dataIn1 = 32'd2806
; 
32'd137409: dataIn1 = 32'd3098
; 
32'd137410: dataIn1 = 32'd3102
; 
32'd137411: dataIn1 = 32'd161
; 
32'd137412: dataIn1 = 32'd1739
; 
32'd137413: dataIn1 = 32'd2803
; 
32'd137414: dataIn1 = 32'd2805
; 
32'd137415: dataIn1 = 32'd2806
; 
32'd137416: dataIn1 = 32'd3091
; 
32'd137417: dataIn1 = 32'd3094
; 
32'd137418: dataIn1 = 32'd1741
; 
32'd137419: dataIn1 = 32'd1742
; 
32'd137420: dataIn1 = 32'd2807
; 
32'd137421: dataIn1 = 32'd2808
; 
32'd137422: dataIn1 = 32'd2809
; 
32'd137423: dataIn1 = 32'd2810
; 
32'd137424: dataIn1 = 32'd2811
; 
32'd137425: dataIn1 = 32'd1742
; 
32'd137426: dataIn1 = 32'd2807
; 
32'd137427: dataIn1 = 32'd2808
; 
32'd137428: dataIn1 = 32'd2809
; 
32'd137429: dataIn1 = 32'd3108
; 
32'd137430: dataIn1 = 32'd11011
; 
32'd137431: dataIn1 = 32'd11012
; 
32'd137432: dataIn1 = 32'd1741
; 
32'd137433: dataIn1 = 32'd2807
; 
32'd137434: dataIn1 = 32'd2808
; 
32'd137435: dataIn1 = 32'd2809
; 
32'd137436: dataIn1 = 32'd3080
; 
32'd137437: dataIn1 = 32'd11010
; 
32'd137438: dataIn1 = 32'd11011
; 
32'd137439: dataIn1 = 32'd159
; 
32'd137440: dataIn1 = 32'd1742
; 
32'd137441: dataIn1 = 32'd2807
; 
32'd137442: dataIn1 = 32'd2810
; 
32'd137443: dataIn1 = 32'd2811
; 
32'd137444: dataIn1 = 32'd3104
; 
32'd137445: dataIn1 = 32'd3107
; 
32'd137446: dataIn1 = 32'd159
; 
32'd137447: dataIn1 = 32'd1741
; 
32'd137448: dataIn1 = 32'd2807
; 
32'd137449: dataIn1 = 32'd2810
; 
32'd137450: dataIn1 = 32'd2811
; 
32'd137451: dataIn1 = 32'd3078
; 
32'd137452: dataIn1 = 32'd3082
; 
32'd137453: dataIn1 = 32'd1744
; 
32'd137454: dataIn1 = 32'd2812
; 
32'd137455: dataIn1 = 32'd2813
; 
32'd137456: dataIn1 = 32'd2814
; 
32'd137457: dataIn1 = 32'd3114
; 
32'd137458: dataIn1 = 32'd11030
; 
32'd137459: dataIn1 = 32'd11031
; 
32'd137460: dataIn1 = 32'd1743
; 
32'd137461: dataIn1 = 32'd1744
; 
32'd137462: dataIn1 = 32'd2812
; 
32'd137463: dataIn1 = 32'd2813
; 
32'd137464: dataIn1 = 32'd2814
; 
32'd137465: dataIn1 = 32'd2815
; 
32'd137466: dataIn1 = 32'd2816
; 
32'd137467: dataIn1 = 32'd1743
; 
32'd137468: dataIn1 = 32'd2812
; 
32'd137469: dataIn1 = 32'd2813
; 
32'd137470: dataIn1 = 32'd2814
; 
32'd137471: dataIn1 = 32'd3124
; 
32'd137472: dataIn1 = 32'd11031
; 
32'd137473: dataIn1 = 32'd11032
; 
32'd137474: dataIn1 = 32'd302
; 
32'd137475: dataIn1 = 32'd1744
; 
32'd137476: dataIn1 = 32'd2813
; 
32'd137477: dataIn1 = 32'd2815
; 
32'd137478: dataIn1 = 32'd2816
; 
32'd137479: dataIn1 = 32'd3112
; 
32'd137480: dataIn1 = 32'd3116
; 
32'd137481: dataIn1 = 32'd302
; 
32'd137482: dataIn1 = 32'd1743
; 
32'd137483: dataIn1 = 32'd2813
; 
32'd137484: dataIn1 = 32'd2815
; 
32'd137485: dataIn1 = 32'd2816
; 
32'd137486: dataIn1 = 32'd3119
; 
32'd137487: dataIn1 = 32'd3122
; 
32'd137488: dataIn1 = 32'd1746
; 
32'd137489: dataIn1 = 32'd2817
; 
32'd137490: dataIn1 = 32'd2818
; 
32'd137491: dataIn1 = 32'd2819
; 
32'd137492: dataIn1 = 32'd3115
; 
32'd137493: dataIn1 = 32'd11027
; 
32'd137494: dataIn1 = 32'd11028
; 
32'd137495: dataIn1 = 32'd1745
; 
32'd137496: dataIn1 = 32'd2817
; 
32'd137497: dataIn1 = 32'd2818
; 
32'd137498: dataIn1 = 32'd2819
; 
32'd137499: dataIn1 = 32'd3088
; 
32'd137500: dataIn1 = 32'd11026
; 
32'd137501: dataIn1 = 32'd11027
; 
32'd137502: dataIn1 = 32'd1745
; 
32'd137503: dataIn1 = 32'd1746
; 
32'd137504: dataIn1 = 32'd2817
; 
32'd137505: dataIn1 = 32'd2818
; 
32'd137506: dataIn1 = 32'd2819
; 
32'd137507: dataIn1 = 32'd2820
; 
32'd137508: dataIn1 = 32'd2821
; 
32'd137509: dataIn1 = 32'd162
; 
32'd137510: dataIn1 = 32'd1746
; 
32'd137511: dataIn1 = 32'd2819
; 
32'd137512: dataIn1 = 32'd2820
; 
32'd137513: dataIn1 = 32'd2821
; 
32'd137514: dataIn1 = 32'd3113
; 
32'd137515: dataIn1 = 32'd3117
; 
32'd137516: dataIn1 = 32'd162
; 
32'd137517: dataIn1 = 32'd1745
; 
32'd137518: dataIn1 = 32'd2819
; 
32'd137519: dataIn1 = 32'd2820
; 
32'd137520: dataIn1 = 32'd2821
; 
32'd137521: dataIn1 = 32'd3085
; 
32'd137522: dataIn1 = 32'd3089
; 
32'd137523: dataIn1 = 32'd1747
; 
32'd137524: dataIn1 = 32'd1748
; 
32'd137525: dataIn1 = 32'd2822
; 
32'd137526: dataIn1 = 32'd2823
; 
32'd137527: dataIn1 = 32'd2824
; 
32'd137528: dataIn1 = 32'd2825
; 
32'd137529: dataIn1 = 32'd2826
; 
32'd137530: dataIn1 = 32'd1748
; 
32'd137531: dataIn1 = 32'd2822
; 
32'd137532: dataIn1 = 32'd2823
; 
32'd137533: dataIn1 = 32'd2824
; 
32'd137534: dataIn1 = 32'd3130
; 
32'd137535: dataIn1 = 32'd11035
; 
32'd137536: dataIn1 = 32'd11036
; 
32'd137537: dataIn1 = 32'd1747
; 
32'd137538: dataIn1 = 32'd2822
; 
32'd137539: dataIn1 = 32'd2823
; 
32'd137540: dataIn1 = 32'd2824
; 
32'd137541: dataIn1 = 32'd3123
; 
32'd137542: dataIn1 = 32'd11034
; 
32'd137543: dataIn1 = 32'd11035
; 
32'd137544: dataIn1 = 32'd163
; 
32'd137545: dataIn1 = 32'd1748
; 
32'd137546: dataIn1 = 32'd2822
; 
32'd137547: dataIn1 = 32'd2825
; 
32'd137548: dataIn1 = 32'd2826
; 
32'd137549: dataIn1 = 32'd3125
; 
32'd137550: dataIn1 = 32'd3128
; 
32'd137551: dataIn1 = 32'd163
; 
32'd137552: dataIn1 = 32'd1747
; 
32'd137553: dataIn1 = 32'd2822
; 
32'd137554: dataIn1 = 32'd2825
; 
32'd137555: dataIn1 = 32'd2826
; 
32'd137556: dataIn1 = 32'd3118
; 
32'd137557: dataIn1 = 32'd3121
; 
32'd137558: dataIn1 = 32'd1750
; 
32'd137559: dataIn1 = 32'd2827
; 
32'd137560: dataIn1 = 32'd2828
; 
32'd137561: dataIn1 = 32'd2829
; 
32'd137562: dataIn1 = 32'd3135
; 
32'd137563: dataIn1 = 32'd11039
; 
32'd137564: dataIn1 = 32'd11040
; 
32'd137565: dataIn1 = 32'd1749
; 
32'd137566: dataIn1 = 32'd1750
; 
32'd137567: dataIn1 = 32'd2827
; 
32'd137568: dataIn1 = 32'd2828
; 
32'd137569: dataIn1 = 32'd2829
; 
32'd137570: dataIn1 = 32'd2830
; 
32'd137571: dataIn1 = 32'd2831
; 
32'd137572: dataIn1 = 32'd1749
; 
32'd137573: dataIn1 = 32'd2827
; 
32'd137574: dataIn1 = 32'd2828
; 
32'd137575: dataIn1 = 32'd2829
; 
32'd137576: dataIn1 = 32'd3131
; 
32'd137577: dataIn1 = 32'd11038
; 
32'd137578: dataIn1 = 32'd11039
; 
32'd137579: dataIn1 = 32'd309
; 
32'd137580: dataIn1 = 32'd1750
; 
32'd137581: dataIn1 = 32'd2828
; 
32'd137582: dataIn1 = 32'd2830
; 
32'd137583: dataIn1 = 32'd2831
; 
32'd137584: dataIn1 = 32'd3133
; 
32'd137585: dataIn1 = 32'd3137
; 
32'd137586: dataIn1 = 32'd309
; 
32'd137587: dataIn1 = 32'd1749
; 
32'd137588: dataIn1 = 32'd2828
; 
32'd137589: dataIn1 = 32'd2830
; 
32'd137590: dataIn1 = 32'd2831
; 
32'd137591: dataIn1 = 32'd3126
; 
32'd137592: dataIn1 = 32'd3129
; 
32'd137593: dataIn1 = 32'd1751
; 
32'd137594: dataIn1 = 32'd1752
; 
32'd137595: dataIn1 = 32'd2832
; 
32'd137596: dataIn1 = 32'd2833
; 
32'd137597: dataIn1 = 32'd2834
; 
32'd137598: dataIn1 = 32'd2835
; 
32'd137599: dataIn1 = 32'd2836
; 
32'd137600: dataIn1 = 32'd1752
; 
32'd137601: dataIn1 = 32'd2832
; 
32'd137602: dataIn1 = 32'd2833
; 
32'd137603: dataIn1 = 32'd2834
; 
32'd137604: dataIn1 = 32'd3143
; 
32'd137605: dataIn1 = 32'd11055
; 
32'd137606: dataIn1 = 32'd11056
; 
32'd137607: dataIn1 = 32'd1751
; 
32'd137608: dataIn1 = 32'd2832
; 
32'd137609: dataIn1 = 32'd2833
; 
32'd137610: dataIn1 = 32'd2834
; 
32'd137611: dataIn1 = 32'd3151
; 
32'd137612: dataIn1 = 32'd11054
; 
32'd137613: dataIn1 = 32'd11055
; 
32'd137614: dataIn1 = 32'd311
; 
32'd137615: dataIn1 = 32'd1752
; 
32'd137616: dataIn1 = 32'd2832
; 
32'd137617: dataIn1 = 32'd2835
; 
32'd137618: dataIn1 = 32'd2836
; 
32'd137619: dataIn1 = 32'd3139
; 
32'd137620: dataIn1 = 32'd3142
; 
32'd137621: dataIn1 = 32'd311
; 
32'd137622: dataIn1 = 32'd1751
; 
32'd137623: dataIn1 = 32'd2832
; 
32'd137624: dataIn1 = 32'd2835
; 
32'd137625: dataIn1 = 32'd2836
; 
32'd137626: dataIn1 = 32'd3146
; 
32'd137627: dataIn1 = 32'd3149
; 
32'd137628: dataIn1 = 32'd1754
; 
32'd137629: dataIn1 = 32'd2837
; 
32'd137630: dataIn1 = 32'd2838
; 
32'd137631: dataIn1 = 32'd2839
; 
32'd137632: dataIn1 = 32'd3157
; 
32'd137633: dataIn1 = 32'd11047
; 
32'd137634: dataIn1 = 32'd11048
; 
32'd137635: dataIn1 = 32'd1753
; 
32'd137636: dataIn1 = 32'd2837
; 
32'd137637: dataIn1 = 32'd2838
; 
32'd137638: dataIn1 = 32'd2839
; 
32'd137639: dataIn1 = 32'd3165
; 
32'd137640: dataIn1 = 32'd11046
; 
32'd137641: dataIn1 = 32'd11047
; 
32'd137642: dataIn1 = 32'd1753
; 
32'd137643: dataIn1 = 32'd1754
; 
32'd137644: dataIn1 = 32'd2837
; 
32'd137645: dataIn1 = 32'd2838
; 
32'd137646: dataIn1 = 32'd2839
; 
32'd137647: dataIn1 = 32'd2840
; 
32'd137648: dataIn1 = 32'd2841
; 
32'd137649: dataIn1 = 32'd317
; 
32'd137650: dataIn1 = 32'd1754
; 
32'd137651: dataIn1 = 32'd2839
; 
32'd137652: dataIn1 = 32'd2840
; 
32'd137653: dataIn1 = 32'd2841
; 
32'd137654: dataIn1 = 32'd3155
; 
32'd137655: dataIn1 = 32'd3159
; 
32'd137656: dataIn1 = 32'd317
; 
32'd137657: dataIn1 = 32'd1753
; 
32'd137658: dataIn1 = 32'd2839
; 
32'd137659: dataIn1 = 32'd2840
; 
32'd137660: dataIn1 = 32'd2841
; 
32'd137661: dataIn1 = 32'd3162
; 
32'd137662: dataIn1 = 32'd3166
; 
32'd137663: dataIn1 = 32'd1756
; 
32'd137664: dataIn1 = 32'd2842
; 
32'd137665: dataIn1 = 32'd2843
; 
32'd137666: dataIn1 = 32'd2844
; 
32'd137667: dataIn1 = 32'd3156
; 
32'd137668: dataIn1 = 32'd11050
; 
32'd137669: dataIn1 = 32'd11051
; 
32'd137670: dataIn1 = 32'd1755
; 
32'd137671: dataIn1 = 32'd1756
; 
32'd137672: dataIn1 = 32'd2842
; 
32'd137673: dataIn1 = 32'd2843
; 
32'd137674: dataIn1 = 32'd2844
; 
32'd137675: dataIn1 = 32'd2845
; 
32'd137676: dataIn1 = 32'd2846
; 
32'd137677: dataIn1 = 32'd1755
; 
32'd137678: dataIn1 = 32'd2842
; 
32'd137679: dataIn1 = 32'd2843
; 
32'd137680: dataIn1 = 32'd2844
; 
32'd137681: dataIn1 = 32'd3152
; 
32'd137682: dataIn1 = 32'd11051
; 
32'd137683: dataIn1 = 32'd11052
; 
32'd137684: dataIn1 = 32'd167
; 
32'd137685: dataIn1 = 32'd1756
; 
32'd137686: dataIn1 = 32'd2843
; 
32'd137687: dataIn1 = 32'd2845
; 
32'd137688: dataIn1 = 32'd2846
; 
32'd137689: dataIn1 = 32'd3154
; 
32'd137690: dataIn1 = 32'd3158
; 
32'd137691: dataIn1 = 32'd167
; 
32'd137692: dataIn1 = 32'd1755
; 
32'd137693: dataIn1 = 32'd2843
; 
32'd137694: dataIn1 = 32'd2845
; 
32'd137695: dataIn1 = 32'd2846
; 
32'd137696: dataIn1 = 32'd3147
; 
32'd137697: dataIn1 = 32'd3150
; 
32'd137698: dataIn1 = 32'd1757
; 
32'd137699: dataIn1 = 32'd1758
; 
32'd137700: dataIn1 = 32'd2847
; 
32'd137701: dataIn1 = 32'd2848
; 
32'd137702: dataIn1 = 32'd2849
; 
32'd137703: dataIn1 = 32'd2850
; 
32'd137704: dataIn1 = 32'd2851
; 
32'd137705: dataIn1 = 32'd1758
; 
32'd137706: dataIn1 = 32'd2847
; 
32'd137707: dataIn1 = 32'd2848
; 
32'd137708: dataIn1 = 32'd2849
; 
32'd137709: dataIn1 = 32'd3164
; 
32'd137710: dataIn1 = 32'd11043
; 
32'd137711: dataIn1 = 32'd11044
; 
32'd137712: dataIn1 = 32'd1757
; 
32'd137713: dataIn1 = 32'd2847
; 
32'd137714: dataIn1 = 32'd2848
; 
32'd137715: dataIn1 = 32'd2849
; 
32'd137716: dataIn1 = 32'd3136
; 
32'd137717: dataIn1 = 32'd11042
; 
32'd137718: dataIn1 = 32'd11043
; 
32'd137719: dataIn1 = 32'd165
; 
32'd137720: dataIn1 = 32'd1758
; 
32'd137721: dataIn1 = 32'd2847
; 
32'd137722: dataIn1 = 32'd2850
; 
32'd137723: dataIn1 = 32'd2851
; 
32'd137724: dataIn1 = 32'd3160
; 
32'd137725: dataIn1 = 32'd3163
; 
32'd137726: dataIn1 = 32'd165
; 
32'd137727: dataIn1 = 32'd1757
; 
32'd137728: dataIn1 = 32'd2847
; 
32'd137729: dataIn1 = 32'd2850
; 
32'd137730: dataIn1 = 32'd2851
; 
32'd137731: dataIn1 = 32'd3134
; 
32'd137732: dataIn1 = 32'd3138
; 
32'd137733: dataIn1 = 32'd1760
; 
32'd137734: dataIn1 = 32'd2852
; 
32'd137735: dataIn1 = 32'd2853
; 
32'd137736: dataIn1 = 32'd2854
; 
32'd137737: dataIn1 = 32'd3170
; 
32'd137738: dataIn1 = 32'd11062
; 
32'd137739: dataIn1 = 32'd11063
; 
32'd137740: dataIn1 = 32'd1759
; 
32'd137741: dataIn1 = 32'd1760
; 
32'd137742: dataIn1 = 32'd2852
; 
32'd137743: dataIn1 = 32'd2853
; 
32'd137744: dataIn1 = 32'd2854
; 
32'd137745: dataIn1 = 32'd2855
; 
32'd137746: dataIn1 = 32'd2856
; 
32'd137747: dataIn1 = 32'd1759
; 
32'd137748: dataIn1 = 32'd2852
; 
32'd137749: dataIn1 = 32'd2853
; 
32'd137750: dataIn1 = 32'd2854
; 
32'd137751: dataIn1 = 32'd3180
; 
32'd137752: dataIn1 = 32'd11063
; 
32'd137753: dataIn1 = 32'd11064
; 
32'd137754: dataIn1 = 32'd318
; 
32'd137755: dataIn1 = 32'd1760
; 
32'd137756: dataIn1 = 32'd2853
; 
32'd137757: dataIn1 = 32'd2855
; 
32'd137758: dataIn1 = 32'd2856
; 
32'd137759: dataIn1 = 32'd3168
; 
32'd137760: dataIn1 = 32'd3172
; 
32'd137761: dataIn1 = 32'd318
; 
32'd137762: dataIn1 = 32'd1759
; 
32'd137763: dataIn1 = 32'd2853
; 
32'd137764: dataIn1 = 32'd2855
; 
32'd137765: dataIn1 = 32'd2856
; 
32'd137766: dataIn1 = 32'd3175
; 
32'd137767: dataIn1 = 32'd3178
; 
32'd137768: dataIn1 = 32'd1762
; 
32'd137769: dataIn1 = 32'd2857
; 
32'd137770: dataIn1 = 32'd2858
; 
32'd137771: dataIn1 = 32'd2859
; 
32'd137772: dataIn1 = 32'd3171
; 
32'd137773: dataIn1 = 32'd11059
; 
32'd137774: dataIn1 = 32'd11060
; 
32'd137775: dataIn1 = 32'd1761
; 
32'd137776: dataIn1 = 32'd2857
; 
32'd137777: dataIn1 = 32'd2858
; 
32'd137778: dataIn1 = 32'd2859
; 
32'd137779: dataIn1 = 32'd3144
; 
32'd137780: dataIn1 = 32'd11058
; 
32'd137781: dataIn1 = 32'd11059
; 
32'd137782: dataIn1 = 32'd1761
; 
32'd137783: dataIn1 = 32'd1762
; 
32'd137784: dataIn1 = 32'd2857
; 
32'd137785: dataIn1 = 32'd2858
; 
32'd137786: dataIn1 = 32'd2859
; 
32'd137787: dataIn1 = 32'd2860
; 
32'd137788: dataIn1 = 32'd2861
; 
32'd137789: dataIn1 = 32'd168
; 
32'd137790: dataIn1 = 32'd1762
; 
32'd137791: dataIn1 = 32'd2859
; 
32'd137792: dataIn1 = 32'd2860
; 
32'd137793: dataIn1 = 32'd2861
; 
32'd137794: dataIn1 = 32'd3169
; 
32'd137795: dataIn1 = 32'd3173
; 
32'd137796: dataIn1 = 32'd168
; 
32'd137797: dataIn1 = 32'd1761
; 
32'd137798: dataIn1 = 32'd2859
; 
32'd137799: dataIn1 = 32'd2860
; 
32'd137800: dataIn1 = 32'd2861
; 
32'd137801: dataIn1 = 32'd3141
; 
32'd137802: dataIn1 = 32'd3145
; 
32'd137803: dataIn1 = 32'd1763
; 
32'd137804: dataIn1 = 32'd1764
; 
32'd137805: dataIn1 = 32'd2862
; 
32'd137806: dataIn1 = 32'd2863
; 
32'd137807: dataIn1 = 32'd2864
; 
32'd137808: dataIn1 = 32'd2865
; 
32'd137809: dataIn1 = 32'd2866
; 
32'd137810: dataIn1 = 32'd1764
; 
32'd137811: dataIn1 = 32'd2862
; 
32'd137812: dataIn1 = 32'd2863
; 
32'd137813: dataIn1 = 32'd2864
; 
32'd137814: dataIn1 = 32'd3186
; 
32'd137815: dataIn1 = 32'd11067
; 
32'd137816: dataIn1 = 32'd11068
; 
32'd137817: dataIn1 = 32'd1763
; 
32'd137818: dataIn1 = 32'd2862
; 
32'd137819: dataIn1 = 32'd2863
; 
32'd137820: dataIn1 = 32'd2864
; 
32'd137821: dataIn1 = 32'd3179
; 
32'd137822: dataIn1 = 32'd11066
; 
32'd137823: dataIn1 = 32'd11067
; 
32'd137824: dataIn1 = 32'd169
; 
32'd137825: dataIn1 = 32'd1764
; 
32'd137826: dataIn1 = 32'd2862
; 
32'd137827: dataIn1 = 32'd2865
; 
32'd137828: dataIn1 = 32'd2866
; 
32'd137829: dataIn1 = 32'd3181
; 
32'd137830: dataIn1 = 32'd3184
; 
32'd137831: dataIn1 = 32'd169
; 
32'd137832: dataIn1 = 32'd1763
; 
32'd137833: dataIn1 = 32'd2862
; 
32'd137834: dataIn1 = 32'd2865
; 
32'd137835: dataIn1 = 32'd2866
; 
32'd137836: dataIn1 = 32'd3174
; 
32'd137837: dataIn1 = 32'd3177
; 
32'd137838: dataIn1 = 32'd1766
; 
32'd137839: dataIn1 = 32'd2867
; 
32'd137840: dataIn1 = 32'd2868
; 
32'd137841: dataIn1 = 32'd2869
; 
32'd137842: dataIn1 = 32'd3191
; 
32'd137843: dataIn1 = 32'd11071
; 
32'd137844: dataIn1 = 32'd11072
; 
32'd137845: dataIn1 = 32'd1765
; 
32'd137846: dataIn1 = 32'd1766
; 
32'd137847: dataIn1 = 32'd2867
; 
32'd137848: dataIn1 = 32'd2868
; 
32'd137849: dataIn1 = 32'd2869
; 
32'd137850: dataIn1 = 32'd2870
; 
32'd137851: dataIn1 = 32'd2871
; 
32'd137852: dataIn1 = 32'd1765
; 
32'd137853: dataIn1 = 32'd2867
; 
32'd137854: dataIn1 = 32'd2868
; 
32'd137855: dataIn1 = 32'd2869
; 
32'd137856: dataIn1 = 32'd3187
; 
32'd137857: dataIn1 = 32'd11070
; 
32'd137858: dataIn1 = 32'd11071
; 
32'd137859: dataIn1 = 32'd325
; 
32'd137860: dataIn1 = 32'd1766
; 
32'd137861: dataIn1 = 32'd2868
; 
32'd137862: dataIn1 = 32'd2870
; 
32'd137863: dataIn1 = 32'd2871
; 
32'd137864: dataIn1 = 32'd3189
; 
32'd137865: dataIn1 = 32'd3193
; 
32'd137866: dataIn1 = 32'd325
; 
32'd137867: dataIn1 = 32'd1765
; 
32'd137868: dataIn1 = 32'd2868
; 
32'd137869: dataIn1 = 32'd2870
; 
32'd137870: dataIn1 = 32'd2871
; 
32'd137871: dataIn1 = 32'd3182
; 
32'd137872: dataIn1 = 32'd3185
; 
32'd137873: dataIn1 = 32'd1767
; 
32'd137874: dataIn1 = 32'd1768
; 
32'd137875: dataIn1 = 32'd2872
; 
32'd137876: dataIn1 = 32'd2873
; 
32'd137877: dataIn1 = 32'd2874
; 
32'd137878: dataIn1 = 32'd2875
; 
32'd137879: dataIn1 = 32'd2876
; 
32'd137880: dataIn1 = 32'd1768
; 
32'd137881: dataIn1 = 32'd2872
; 
32'd137882: dataIn1 = 32'd2873
; 
32'd137883: dataIn1 = 32'd2874
; 
32'd137884: dataIn1 = 32'd3199
; 
32'd137885: dataIn1 = 32'd11087
; 
32'd137886: dataIn1 = 32'd11088
; 
32'd137887: dataIn1 = 32'd1767
; 
32'd137888: dataIn1 = 32'd2872
; 
32'd137889: dataIn1 = 32'd2873
; 
32'd137890: dataIn1 = 32'd2874
; 
32'd137891: dataIn1 = 32'd3207
; 
32'd137892: dataIn1 = 32'd11086
; 
32'd137893: dataIn1 = 32'd11087
; 
32'd137894: dataIn1 = 32'd327
; 
32'd137895: dataIn1 = 32'd1768
; 
32'd137896: dataIn1 = 32'd2872
; 
32'd137897: dataIn1 = 32'd2875
; 
32'd137898: dataIn1 = 32'd2876
; 
32'd137899: dataIn1 = 32'd3195
; 
32'd137900: dataIn1 = 32'd3198
; 
32'd137901: dataIn1 = 32'd327
; 
32'd137902: dataIn1 = 32'd1767
; 
32'd137903: dataIn1 = 32'd2872
; 
32'd137904: dataIn1 = 32'd2875
; 
32'd137905: dataIn1 = 32'd2876
; 
32'd137906: dataIn1 = 32'd3202
; 
32'd137907: dataIn1 = 32'd3205
; 
32'd137908: dataIn1 = 32'd1770
; 
32'd137909: dataIn1 = 32'd2877
; 
32'd137910: dataIn1 = 32'd2878
; 
32'd137911: dataIn1 = 32'd2879
; 
32'd137912: dataIn1 = 32'd3213
; 
32'd137913: dataIn1 = 32'd11079
; 
32'd137914: dataIn1 = 32'd11080
; 
32'd137915: dataIn1 = 32'd1769
; 
32'd137916: dataIn1 = 32'd2877
; 
32'd137917: dataIn1 = 32'd2878
; 
32'd137918: dataIn1 = 32'd2879
; 
32'd137919: dataIn1 = 32'd3221
; 
32'd137920: dataIn1 = 32'd11078
; 
32'd137921: dataIn1 = 32'd11079
; 
32'd137922: dataIn1 = 32'd1769
; 
32'd137923: dataIn1 = 32'd1770
; 
32'd137924: dataIn1 = 32'd2877
; 
32'd137925: dataIn1 = 32'd2878
; 
32'd137926: dataIn1 = 32'd2879
; 
32'd137927: dataIn1 = 32'd2880
; 
32'd137928: dataIn1 = 32'd2881
; 
32'd137929: dataIn1 = 32'd333
; 
32'd137930: dataIn1 = 32'd1770
; 
32'd137931: dataIn1 = 32'd2879
; 
32'd137932: dataIn1 = 32'd2880
; 
32'd137933: dataIn1 = 32'd2881
; 
32'd137934: dataIn1 = 32'd3211
; 
32'd137935: dataIn1 = 32'd3215
; 
32'd137936: dataIn1 = 32'd333
; 
32'd137937: dataIn1 = 32'd1769
; 
32'd137938: dataIn1 = 32'd2879
; 
32'd137939: dataIn1 = 32'd2880
; 
32'd137940: dataIn1 = 32'd2881
; 
32'd137941: dataIn1 = 32'd3218
; 
32'd137942: dataIn1 = 32'd3222
; 
32'd137943: dataIn1 = 32'd1772
; 
32'd137944: dataIn1 = 32'd2882
; 
32'd137945: dataIn1 = 32'd2883
; 
32'd137946: dataIn1 = 32'd2884
; 
32'd137947: dataIn1 = 32'd3212
; 
32'd137948: dataIn1 = 32'd11082
; 
32'd137949: dataIn1 = 32'd11083
; 
32'd137950: dataIn1 = 32'd1771
; 
32'd137951: dataIn1 = 32'd1772
; 
32'd137952: dataIn1 = 32'd2882
; 
32'd137953: dataIn1 = 32'd2883
; 
32'd137954: dataIn1 = 32'd2884
; 
32'd137955: dataIn1 = 32'd2885
; 
32'd137956: dataIn1 = 32'd2886
; 
32'd137957: dataIn1 = 32'd1771
; 
32'd137958: dataIn1 = 32'd2882
; 
32'd137959: dataIn1 = 32'd2883
; 
32'd137960: dataIn1 = 32'd2884
; 
32'd137961: dataIn1 = 32'd3208
; 
32'd137962: dataIn1 = 32'd11083
; 
32'd137963: dataIn1 = 32'd11084
; 
32'd137964: dataIn1 = 32'd173
; 
32'd137965: dataIn1 = 32'd1772
; 
32'd137966: dataIn1 = 32'd2883
; 
32'd137967: dataIn1 = 32'd2885
; 
32'd137968: dataIn1 = 32'd2886
; 
32'd137969: dataIn1 = 32'd3210
; 
32'd137970: dataIn1 = 32'd3214
; 
32'd137971: dataIn1 = 32'd173
; 
32'd137972: dataIn1 = 32'd1771
; 
32'd137973: dataIn1 = 32'd2883
; 
32'd137974: dataIn1 = 32'd2885
; 
32'd137975: dataIn1 = 32'd2886
; 
32'd137976: dataIn1 = 32'd3203
; 
32'd137977: dataIn1 = 32'd3206
; 
32'd137978: dataIn1 = 32'd1773
; 
32'd137979: dataIn1 = 32'd1774
; 
32'd137980: dataIn1 = 32'd2887
; 
32'd137981: dataIn1 = 32'd2888
; 
32'd137982: dataIn1 = 32'd2889
; 
32'd137983: dataIn1 = 32'd2890
; 
32'd137984: dataIn1 = 32'd2891
; 
32'd137985: dataIn1 = 32'd1774
; 
32'd137986: dataIn1 = 32'd2887
; 
32'd137987: dataIn1 = 32'd2888
; 
32'd137988: dataIn1 = 32'd2889
; 
32'd137989: dataIn1 = 32'd3220
; 
32'd137990: dataIn1 = 32'd11075
; 
32'd137991: dataIn1 = 32'd11076
; 
32'd137992: dataIn1 = 32'd1773
; 
32'd137993: dataIn1 = 32'd2887
; 
32'd137994: dataIn1 = 32'd2888
; 
32'd137995: dataIn1 = 32'd2889
; 
32'd137996: dataIn1 = 32'd3192
; 
32'd137997: dataIn1 = 32'd11074
; 
32'd137998: dataIn1 = 32'd11075
; 
32'd137999: dataIn1 = 32'd171
; 
32'd138000: dataIn1 = 32'd1774
; 
32'd138001: dataIn1 = 32'd2887
; 
32'd138002: dataIn1 = 32'd2890
; 
32'd138003: dataIn1 = 32'd2891
; 
32'd138004: dataIn1 = 32'd3216
; 
32'd138005: dataIn1 = 32'd3219
; 
32'd138006: dataIn1 = 32'd171
; 
32'd138007: dataIn1 = 32'd1773
; 
32'd138008: dataIn1 = 32'd2887
; 
32'd138009: dataIn1 = 32'd2890
; 
32'd138010: dataIn1 = 32'd2891
; 
32'd138011: dataIn1 = 32'd3190
; 
32'd138012: dataIn1 = 32'd3194
; 
32'd138013: dataIn1 = 32'd1776
; 
32'd138014: dataIn1 = 32'd2892
; 
32'd138015: dataIn1 = 32'd2893
; 
32'd138016: dataIn1 = 32'd2894
; 
32'd138017: dataIn1 = 32'd3226
; 
32'd138018: dataIn1 = 32'd11094
; 
32'd138019: dataIn1 = 32'd11095
; 
32'd138020: dataIn1 = 32'd1775
; 
32'd138021: dataIn1 = 32'd1776
; 
32'd138022: dataIn1 = 32'd2892
; 
32'd138023: dataIn1 = 32'd2893
; 
32'd138024: dataIn1 = 32'd2894
; 
32'd138025: dataIn1 = 32'd2895
; 
32'd138026: dataIn1 = 32'd2896
; 
32'd138027: dataIn1 = 32'd1775
; 
32'd138028: dataIn1 = 32'd2892
; 
32'd138029: dataIn1 = 32'd2893
; 
32'd138030: dataIn1 = 32'd2894
; 
32'd138031: dataIn1 = 32'd3236
; 
32'd138032: dataIn1 = 32'd11095
; 
32'd138033: dataIn1 = 32'd11096
; 
32'd138034: dataIn1 = 32'd334
; 
32'd138035: dataIn1 = 32'd1776
; 
32'd138036: dataIn1 = 32'd2893
; 
32'd138037: dataIn1 = 32'd2895
; 
32'd138038: dataIn1 = 32'd2896
; 
32'd138039: dataIn1 = 32'd3224
; 
32'd138040: dataIn1 = 32'd3228
; 
32'd138041: dataIn1 = 32'd334
; 
32'd138042: dataIn1 = 32'd1775
; 
32'd138043: dataIn1 = 32'd2893
; 
32'd138044: dataIn1 = 32'd2895
; 
32'd138045: dataIn1 = 32'd2896
; 
32'd138046: dataIn1 = 32'd3231
; 
32'd138047: dataIn1 = 32'd3234
; 
32'd138048: dataIn1 = 32'd1778
; 
32'd138049: dataIn1 = 32'd2897
; 
32'd138050: dataIn1 = 32'd2898
; 
32'd138051: dataIn1 = 32'd2899
; 
32'd138052: dataIn1 = 32'd3227
; 
32'd138053: dataIn1 = 32'd11091
; 
32'd138054: dataIn1 = 32'd11092
; 
32'd138055: dataIn1 = 32'd1777
; 
32'd138056: dataIn1 = 32'd2897
; 
32'd138057: dataIn1 = 32'd2898
; 
32'd138058: dataIn1 = 32'd2899
; 
32'd138059: dataIn1 = 32'd3200
; 
32'd138060: dataIn1 = 32'd11090
; 
32'd138061: dataIn1 = 32'd11091
; 
32'd138062: dataIn1 = 32'd1777
; 
32'd138063: dataIn1 = 32'd1778
; 
32'd138064: dataIn1 = 32'd2897
; 
32'd138065: dataIn1 = 32'd2898
; 
32'd138066: dataIn1 = 32'd2899
; 
32'd138067: dataIn1 = 32'd2900
; 
32'd138068: dataIn1 = 32'd2901
; 
32'd138069: dataIn1 = 32'd174
; 
32'd138070: dataIn1 = 32'd1778
; 
32'd138071: dataIn1 = 32'd2899
; 
32'd138072: dataIn1 = 32'd2900
; 
32'd138073: dataIn1 = 32'd2901
; 
32'd138074: dataIn1 = 32'd3225
; 
32'd138075: dataIn1 = 32'd3229
; 
32'd138076: dataIn1 = 32'd174
; 
32'd138077: dataIn1 = 32'd1777
; 
32'd138078: dataIn1 = 32'd2899
; 
32'd138079: dataIn1 = 32'd2900
; 
32'd138080: dataIn1 = 32'd2901
; 
32'd138081: dataIn1 = 32'd3197
; 
32'd138082: dataIn1 = 32'd3201
; 
32'd138083: dataIn1 = 32'd1779
; 
32'd138084: dataIn1 = 32'd1780
; 
32'd138085: dataIn1 = 32'd2902
; 
32'd138086: dataIn1 = 32'd2903
; 
32'd138087: dataIn1 = 32'd2904
; 
32'd138088: dataIn1 = 32'd2905
; 
32'd138089: dataIn1 = 32'd2906
; 
32'd138090: dataIn1 = 32'd1780
; 
32'd138091: dataIn1 = 32'd2902
; 
32'd138092: dataIn1 = 32'd2903
; 
32'd138093: dataIn1 = 32'd2904
; 
32'd138094: dataIn1 = 32'd3242
; 
32'd138095: dataIn1 = 32'd11099
; 
32'd138096: dataIn1 = 32'd11100
; 
32'd138097: dataIn1 = 32'd1779
; 
32'd138098: dataIn1 = 32'd2902
; 
32'd138099: dataIn1 = 32'd2903
; 
32'd138100: dataIn1 = 32'd2904
; 
32'd138101: dataIn1 = 32'd3235
; 
32'd138102: dataIn1 = 32'd11098
; 
32'd138103: dataIn1 = 32'd11099
; 
32'd138104: dataIn1 = 32'd175
; 
32'd138105: dataIn1 = 32'd1780
; 
32'd138106: dataIn1 = 32'd2902
; 
32'd138107: dataIn1 = 32'd2905
; 
32'd138108: dataIn1 = 32'd2906
; 
32'd138109: dataIn1 = 32'd3237
; 
32'd138110: dataIn1 = 32'd3240
; 
32'd138111: dataIn1 = 32'd175
; 
32'd138112: dataIn1 = 32'd1779
; 
32'd138113: dataIn1 = 32'd2902
; 
32'd138114: dataIn1 = 32'd2905
; 
32'd138115: dataIn1 = 32'd2906
; 
32'd138116: dataIn1 = 32'd3230
; 
32'd138117: dataIn1 = 32'd3233
; 
32'd138118: dataIn1 = 32'd1782
; 
32'd138119: dataIn1 = 32'd2907
; 
32'd138120: dataIn1 = 32'd2908
; 
32'd138121: dataIn1 = 32'd2909
; 
32'd138122: dataIn1 = 32'd3247
; 
32'd138123: dataIn1 = 32'd11103
; 
32'd138124: dataIn1 = 32'd11104
; 
32'd138125: dataIn1 = 32'd1781
; 
32'd138126: dataIn1 = 32'd1782
; 
32'd138127: dataIn1 = 32'd2907
; 
32'd138128: dataIn1 = 32'd2908
; 
32'd138129: dataIn1 = 32'd2909
; 
32'd138130: dataIn1 = 32'd2910
; 
32'd138131: dataIn1 = 32'd2911
; 
32'd138132: dataIn1 = 32'd1781
; 
32'd138133: dataIn1 = 32'd2907
; 
32'd138134: dataIn1 = 32'd2908
; 
32'd138135: dataIn1 = 32'd2909
; 
32'd138136: dataIn1 = 32'd3243
; 
32'd138137: dataIn1 = 32'd11102
; 
32'd138138: dataIn1 = 32'd11103
; 
32'd138139: dataIn1 = 32'd341
; 
32'd138140: dataIn1 = 32'd1782
; 
32'd138141: dataIn1 = 32'd2908
; 
32'd138142: dataIn1 = 32'd2910
; 
32'd138143: dataIn1 = 32'd2911
; 
32'd138144: dataIn1 = 32'd3245
; 
32'd138145: dataIn1 = 32'd3249
; 
32'd138146: dataIn1 = 32'd341
; 
32'd138147: dataIn1 = 32'd1781
; 
32'd138148: dataIn1 = 32'd2908
; 
32'd138149: dataIn1 = 32'd2910
; 
32'd138150: dataIn1 = 32'd2911
; 
32'd138151: dataIn1 = 32'd3238
; 
32'd138152: dataIn1 = 32'd3241
; 
32'd138153: dataIn1 = 32'd1783
; 
32'd138154: dataIn1 = 32'd1784
; 
32'd138155: dataIn1 = 32'd2912
; 
32'd138156: dataIn1 = 32'd2913
; 
32'd138157: dataIn1 = 32'd2914
; 
32'd138158: dataIn1 = 32'd2915
; 
32'd138159: dataIn1 = 32'd2916
; 
32'd138160: dataIn1 = 32'd1784
; 
32'd138161: dataIn1 = 32'd2912
; 
32'd138162: dataIn1 = 32'd2913
; 
32'd138163: dataIn1 = 32'd2914
; 
32'd138164: dataIn1 = 32'd3255
; 
32'd138165: dataIn1 = 32'd11119
; 
32'd138166: dataIn1 = 32'd11120
; 
32'd138167: dataIn1 = 32'd1783
; 
32'd138168: dataIn1 = 32'd2912
; 
32'd138169: dataIn1 = 32'd2913
; 
32'd138170: dataIn1 = 32'd2914
; 
32'd138171: dataIn1 = 32'd3263
; 
32'd138172: dataIn1 = 32'd11118
; 
32'd138173: dataIn1 = 32'd11119
; 
32'd138174: dataIn1 = 32'd343
; 
32'd138175: dataIn1 = 32'd1784
; 
32'd138176: dataIn1 = 32'd2912
; 
32'd138177: dataIn1 = 32'd2915
; 
32'd138178: dataIn1 = 32'd2916
; 
32'd138179: dataIn1 = 32'd3251
; 
32'd138180: dataIn1 = 32'd3254
; 
32'd138181: dataIn1 = 32'd343
; 
32'd138182: dataIn1 = 32'd1783
; 
32'd138183: dataIn1 = 32'd2912
; 
32'd138184: dataIn1 = 32'd2915
; 
32'd138185: dataIn1 = 32'd2916
; 
32'd138186: dataIn1 = 32'd3258
; 
32'd138187: dataIn1 = 32'd3261
; 
32'd138188: dataIn1 = 32'd1786
; 
32'd138189: dataIn1 = 32'd2917
; 
32'd138190: dataIn1 = 32'd2918
; 
32'd138191: dataIn1 = 32'd2919
; 
32'd138192: dataIn1 = 32'd3269
; 
32'd138193: dataIn1 = 32'd11111
; 
32'd138194: dataIn1 = 32'd11112
; 
32'd138195: dataIn1 = 32'd1785
; 
32'd138196: dataIn1 = 32'd2917
; 
32'd138197: dataIn1 = 32'd2918
; 
32'd138198: dataIn1 = 32'd2919
; 
32'd138199: dataIn1 = 32'd3277
; 
32'd138200: dataIn1 = 32'd11110
; 
32'd138201: dataIn1 = 32'd11111
; 
32'd138202: dataIn1 = 32'd1785
; 
32'd138203: dataIn1 = 32'd1786
; 
32'd138204: dataIn1 = 32'd2917
; 
32'd138205: dataIn1 = 32'd2918
; 
32'd138206: dataIn1 = 32'd2919
; 
32'd138207: dataIn1 = 32'd2920
; 
32'd138208: dataIn1 = 32'd2921
; 
32'd138209: dataIn1 = 32'd349
; 
32'd138210: dataIn1 = 32'd1786
; 
32'd138211: dataIn1 = 32'd2919
; 
32'd138212: dataIn1 = 32'd2920
; 
32'd138213: dataIn1 = 32'd2921
; 
32'd138214: dataIn1 = 32'd3267
; 
32'd138215: dataIn1 = 32'd3271
; 
32'd138216: dataIn1 = 32'd349
; 
32'd138217: dataIn1 = 32'd1785
; 
32'd138218: dataIn1 = 32'd2919
; 
32'd138219: dataIn1 = 32'd2920
; 
32'd138220: dataIn1 = 32'd2921
; 
32'd138221: dataIn1 = 32'd3274
; 
32'd138222: dataIn1 = 32'd3278
; 
32'd138223: dataIn1 = 32'd1788
; 
32'd138224: dataIn1 = 32'd2922
; 
32'd138225: dataIn1 = 32'd2923
; 
32'd138226: dataIn1 = 32'd2924
; 
32'd138227: dataIn1 = 32'd3268
; 
32'd138228: dataIn1 = 32'd11114
; 
32'd138229: dataIn1 = 32'd11115
; 
32'd138230: dataIn1 = 32'd1787
; 
32'd138231: dataIn1 = 32'd1788
; 
32'd138232: dataIn1 = 32'd2922
; 
32'd138233: dataIn1 = 32'd2923
; 
32'd138234: dataIn1 = 32'd2924
; 
32'd138235: dataIn1 = 32'd2925
; 
32'd138236: dataIn1 = 32'd2926
; 
32'd138237: dataIn1 = 32'd1787
; 
32'd138238: dataIn1 = 32'd2922
; 
32'd138239: dataIn1 = 32'd2923
; 
32'd138240: dataIn1 = 32'd2924
; 
32'd138241: dataIn1 = 32'd3264
; 
32'd138242: dataIn1 = 32'd11115
; 
32'd138243: dataIn1 = 32'd11116
; 
32'd138244: dataIn1 = 32'd179
; 
32'd138245: dataIn1 = 32'd1788
; 
32'd138246: dataIn1 = 32'd2923
; 
32'd138247: dataIn1 = 32'd2925
; 
32'd138248: dataIn1 = 32'd2926
; 
32'd138249: dataIn1 = 32'd3266
; 
32'd138250: dataIn1 = 32'd3270
; 
32'd138251: dataIn1 = 32'd179
; 
32'd138252: dataIn1 = 32'd1787
; 
32'd138253: dataIn1 = 32'd2923
; 
32'd138254: dataIn1 = 32'd2925
; 
32'd138255: dataIn1 = 32'd2926
; 
32'd138256: dataIn1 = 32'd3259
; 
32'd138257: dataIn1 = 32'd3262
; 
32'd138258: dataIn1 = 32'd1789
; 
32'd138259: dataIn1 = 32'd1790
; 
32'd138260: dataIn1 = 32'd2927
; 
32'd138261: dataIn1 = 32'd2928
; 
32'd138262: dataIn1 = 32'd2929
; 
32'd138263: dataIn1 = 32'd2930
; 
32'd138264: dataIn1 = 32'd2931
; 
32'd138265: dataIn1 = 32'd1790
; 
32'd138266: dataIn1 = 32'd2927
; 
32'd138267: dataIn1 = 32'd2928
; 
32'd138268: dataIn1 = 32'd2929
; 
32'd138269: dataIn1 = 32'd3276
; 
32'd138270: dataIn1 = 32'd11107
; 
32'd138271: dataIn1 = 32'd11108
; 
32'd138272: dataIn1 = 32'd1789
; 
32'd138273: dataIn1 = 32'd2927
; 
32'd138274: dataIn1 = 32'd2928
; 
32'd138275: dataIn1 = 32'd2929
; 
32'd138276: dataIn1 = 32'd3248
; 
32'd138277: dataIn1 = 32'd11106
; 
32'd138278: dataIn1 = 32'd11107
; 
32'd138279: dataIn1 = 32'd177
; 
32'd138280: dataIn1 = 32'd1790
; 
32'd138281: dataIn1 = 32'd2927
; 
32'd138282: dataIn1 = 32'd2930
; 
32'd138283: dataIn1 = 32'd2931
; 
32'd138284: dataIn1 = 32'd3272
; 
32'd138285: dataIn1 = 32'd3275
; 
32'd138286: dataIn1 = 32'd177
; 
32'd138287: dataIn1 = 32'd1789
; 
32'd138288: dataIn1 = 32'd2927
; 
32'd138289: dataIn1 = 32'd2930
; 
32'd138290: dataIn1 = 32'd2931
; 
32'd138291: dataIn1 = 32'd3246
; 
32'd138292: dataIn1 = 32'd3250
; 
32'd138293: dataIn1 = 32'd1792
; 
32'd138294: dataIn1 = 32'd2932
; 
32'd138295: dataIn1 = 32'd2933
; 
32'd138296: dataIn1 = 32'd2934
; 
32'd138297: dataIn1 = 32'd3282
; 
32'd138298: dataIn1 = 32'd11126
; 
32'd138299: dataIn1 = 32'd11127
; 
32'd138300: dataIn1 = 32'd1791
; 
32'd138301: dataIn1 = 32'd1792
; 
32'd138302: dataIn1 = 32'd2932
; 
32'd138303: dataIn1 = 32'd2933
; 
32'd138304: dataIn1 = 32'd2934
; 
32'd138305: dataIn1 = 32'd2935
; 
32'd138306: dataIn1 = 32'd2936
; 
32'd138307: dataIn1 = 32'd1791
; 
32'd138308: dataIn1 = 32'd2932
; 
32'd138309: dataIn1 = 32'd2933
; 
32'd138310: dataIn1 = 32'd2934
; 
32'd138311: dataIn1 = 32'd3292
; 
32'd138312: dataIn1 = 32'd11127
; 
32'd138313: dataIn1 = 32'd11128
; 
32'd138314: dataIn1 = 32'd350
; 
32'd138315: dataIn1 = 32'd1792
; 
32'd138316: dataIn1 = 32'd2933
; 
32'd138317: dataIn1 = 32'd2935
; 
32'd138318: dataIn1 = 32'd2936
; 
32'd138319: dataIn1 = 32'd3280
; 
32'd138320: dataIn1 = 32'd3284
; 
32'd138321: dataIn1 = 32'd350
; 
32'd138322: dataIn1 = 32'd1791
; 
32'd138323: dataIn1 = 32'd2933
; 
32'd138324: dataIn1 = 32'd2935
; 
32'd138325: dataIn1 = 32'd2936
; 
32'd138326: dataIn1 = 32'd3287
; 
32'd138327: dataIn1 = 32'd3290
; 
32'd138328: dataIn1 = 32'd1794
; 
32'd138329: dataIn1 = 32'd2937
; 
32'd138330: dataIn1 = 32'd2938
; 
32'd138331: dataIn1 = 32'd2939
; 
32'd138332: dataIn1 = 32'd3283
; 
32'd138333: dataIn1 = 32'd11123
; 
32'd138334: dataIn1 = 32'd11124
; 
32'd138335: dataIn1 = 32'd1793
; 
32'd138336: dataIn1 = 32'd2937
; 
32'd138337: dataIn1 = 32'd2938
; 
32'd138338: dataIn1 = 32'd2939
; 
32'd138339: dataIn1 = 32'd3256
; 
32'd138340: dataIn1 = 32'd11122
; 
32'd138341: dataIn1 = 32'd11123
; 
32'd138342: dataIn1 = 32'd1793
; 
32'd138343: dataIn1 = 32'd1794
; 
32'd138344: dataIn1 = 32'd2937
; 
32'd138345: dataIn1 = 32'd2938
; 
32'd138346: dataIn1 = 32'd2939
; 
32'd138347: dataIn1 = 32'd2940
; 
32'd138348: dataIn1 = 32'd2941
; 
32'd138349: dataIn1 = 32'd180
; 
32'd138350: dataIn1 = 32'd1794
; 
32'd138351: dataIn1 = 32'd2939
; 
32'd138352: dataIn1 = 32'd2940
; 
32'd138353: dataIn1 = 32'd2941
; 
32'd138354: dataIn1 = 32'd3281
; 
32'd138355: dataIn1 = 32'd3285
; 
32'd138356: dataIn1 = 32'd180
; 
32'd138357: dataIn1 = 32'd1793
; 
32'd138358: dataIn1 = 32'd2939
; 
32'd138359: dataIn1 = 32'd2940
; 
32'd138360: dataIn1 = 32'd2941
; 
32'd138361: dataIn1 = 32'd3253
; 
32'd138362: dataIn1 = 32'd3257
; 
32'd138363: dataIn1 = 32'd1795
; 
32'd138364: dataIn1 = 32'd1796
; 
32'd138365: dataIn1 = 32'd2942
; 
32'd138366: dataIn1 = 32'd2943
; 
32'd138367: dataIn1 = 32'd2944
; 
32'd138368: dataIn1 = 32'd2945
; 
32'd138369: dataIn1 = 32'd2946
; 
32'd138370: dataIn1 = 32'd1796
; 
32'd138371: dataIn1 = 32'd2942
; 
32'd138372: dataIn1 = 32'd2943
; 
32'd138373: dataIn1 = 32'd2944
; 
32'd138374: dataIn1 = 32'd3298
; 
32'd138375: dataIn1 = 32'd11131
; 
32'd138376: dataIn1 = 32'd11132
; 
32'd138377: dataIn1 = 32'd1795
; 
32'd138378: dataIn1 = 32'd2942
; 
32'd138379: dataIn1 = 32'd2943
; 
32'd138380: dataIn1 = 32'd2944
; 
32'd138381: dataIn1 = 32'd3291
; 
32'd138382: dataIn1 = 32'd11130
; 
32'd138383: dataIn1 = 32'd11131
; 
32'd138384: dataIn1 = 32'd181
; 
32'd138385: dataIn1 = 32'd1796
; 
32'd138386: dataIn1 = 32'd2942
; 
32'd138387: dataIn1 = 32'd2945
; 
32'd138388: dataIn1 = 32'd2946
; 
32'd138389: dataIn1 = 32'd3293
; 
32'd138390: dataIn1 = 32'd3296
; 
32'd138391: dataIn1 = 32'd181
; 
32'd138392: dataIn1 = 32'd1795
; 
32'd138393: dataIn1 = 32'd2942
; 
32'd138394: dataIn1 = 32'd2945
; 
32'd138395: dataIn1 = 32'd2946
; 
32'd138396: dataIn1 = 32'd3286
; 
32'd138397: dataIn1 = 32'd3289
; 
32'd138398: dataIn1 = 32'd1798
; 
32'd138399: dataIn1 = 32'd2947
; 
32'd138400: dataIn1 = 32'd2948
; 
32'd138401: dataIn1 = 32'd2949
; 
32'd138402: dataIn1 = 32'd3303
; 
32'd138403: dataIn1 = 32'd11135
; 
32'd138404: dataIn1 = 32'd11136
; 
32'd138405: dataIn1 = 32'd1797
; 
32'd138406: dataIn1 = 32'd1798
; 
32'd138407: dataIn1 = 32'd2947
; 
32'd138408: dataIn1 = 32'd2948
; 
32'd138409: dataIn1 = 32'd2949
; 
32'd138410: dataIn1 = 32'd2950
; 
32'd138411: dataIn1 = 32'd2951
; 
32'd138412: dataIn1 = 32'd1797
; 
32'd138413: dataIn1 = 32'd2947
; 
32'd138414: dataIn1 = 32'd2948
; 
32'd138415: dataIn1 = 32'd2949
; 
32'd138416: dataIn1 = 32'd3299
; 
32'd138417: dataIn1 = 32'd11134
; 
32'd138418: dataIn1 = 32'd11135
; 
32'd138419: dataIn1 = 32'd357
; 
32'd138420: dataIn1 = 32'd1798
; 
32'd138421: dataIn1 = 32'd2948
; 
32'd138422: dataIn1 = 32'd2950
; 
32'd138423: dataIn1 = 32'd2951
; 
32'd138424: dataIn1 = 32'd3301
; 
32'd138425: dataIn1 = 32'd3305
; 
32'd138426: dataIn1 = 32'd357
; 
32'd138427: dataIn1 = 32'd1797
; 
32'd138428: dataIn1 = 32'd2948
; 
32'd138429: dataIn1 = 32'd2950
; 
32'd138430: dataIn1 = 32'd2951
; 
32'd138431: dataIn1 = 32'd3294
; 
32'd138432: dataIn1 = 32'd3297
; 
32'd138433: dataIn1 = 32'd1799
; 
32'd138434: dataIn1 = 32'd1800
; 
32'd138435: dataIn1 = 32'd2952
; 
32'd138436: dataIn1 = 32'd2953
; 
32'd138437: dataIn1 = 32'd2954
; 
32'd138438: dataIn1 = 32'd2955
; 
32'd138439: dataIn1 = 32'd2956
; 
32'd138440: dataIn1 = 32'd1800
; 
32'd138441: dataIn1 = 32'd2952
; 
32'd138442: dataIn1 = 32'd2953
; 
32'd138443: dataIn1 = 32'd2954
; 
32'd138444: dataIn1 = 32'd3311
; 
32'd138445: dataIn1 = 32'd11151
; 
32'd138446: dataIn1 = 32'd11152
; 
32'd138447: dataIn1 = 32'd1799
; 
32'd138448: dataIn1 = 32'd2952
; 
32'd138449: dataIn1 = 32'd2953
; 
32'd138450: dataIn1 = 32'd2954
; 
32'd138451: dataIn1 = 32'd3319
; 
32'd138452: dataIn1 = 32'd11150
; 
32'd138453: dataIn1 = 32'd11151
; 
32'd138454: dataIn1 = 32'd359
; 
32'd138455: dataIn1 = 32'd1800
; 
32'd138456: dataIn1 = 32'd2952
; 
32'd138457: dataIn1 = 32'd2955
; 
32'd138458: dataIn1 = 32'd2956
; 
32'd138459: dataIn1 = 32'd3307
; 
32'd138460: dataIn1 = 32'd3310
; 
32'd138461: dataIn1 = 32'd359
; 
32'd138462: dataIn1 = 32'd1799
; 
32'd138463: dataIn1 = 32'd2952
; 
32'd138464: dataIn1 = 32'd2955
; 
32'd138465: dataIn1 = 32'd2956
; 
32'd138466: dataIn1 = 32'd3314
; 
32'd138467: dataIn1 = 32'd3317
; 
32'd138468: dataIn1 = 32'd1802
; 
32'd138469: dataIn1 = 32'd2957
; 
32'd138470: dataIn1 = 32'd2958
; 
32'd138471: dataIn1 = 32'd2959
; 
32'd138472: dataIn1 = 32'd3325
; 
32'd138473: dataIn1 = 32'd11143
; 
32'd138474: dataIn1 = 32'd11144
; 
32'd138475: dataIn1 = 32'd1801
; 
32'd138476: dataIn1 = 32'd2957
; 
32'd138477: dataIn1 = 32'd2958
; 
32'd138478: dataIn1 = 32'd2959
; 
32'd138479: dataIn1 = 32'd3333
; 
32'd138480: dataIn1 = 32'd11142
; 
32'd138481: dataIn1 = 32'd11143
; 
32'd138482: dataIn1 = 32'd1801
; 
32'd138483: dataIn1 = 32'd1802
; 
32'd138484: dataIn1 = 32'd2957
; 
32'd138485: dataIn1 = 32'd2958
; 
32'd138486: dataIn1 = 32'd2959
; 
32'd138487: dataIn1 = 32'd2960
; 
32'd138488: dataIn1 = 32'd2961
; 
32'd138489: dataIn1 = 32'd365
; 
32'd138490: dataIn1 = 32'd1802
; 
32'd138491: dataIn1 = 32'd2959
; 
32'd138492: dataIn1 = 32'd2960
; 
32'd138493: dataIn1 = 32'd2961
; 
32'd138494: dataIn1 = 32'd3323
; 
32'd138495: dataIn1 = 32'd3327
; 
32'd138496: dataIn1 = 32'd365
; 
32'd138497: dataIn1 = 32'd1801
; 
32'd138498: dataIn1 = 32'd2959
; 
32'd138499: dataIn1 = 32'd2960
; 
32'd138500: dataIn1 = 32'd2961
; 
32'd138501: dataIn1 = 32'd3330
; 
32'd138502: dataIn1 = 32'd3334
; 
32'd138503: dataIn1 = 32'd1804
; 
32'd138504: dataIn1 = 32'd2962
; 
32'd138505: dataIn1 = 32'd2963
; 
32'd138506: dataIn1 = 32'd2964
; 
32'd138507: dataIn1 = 32'd3324
; 
32'd138508: dataIn1 = 32'd11146
; 
32'd138509: dataIn1 = 32'd11147
; 
32'd138510: dataIn1 = 32'd1803
; 
32'd138511: dataIn1 = 32'd1804
; 
32'd138512: dataIn1 = 32'd2962
; 
32'd138513: dataIn1 = 32'd2963
; 
32'd138514: dataIn1 = 32'd2964
; 
32'd138515: dataIn1 = 32'd2965
; 
32'd138516: dataIn1 = 32'd2966
; 
32'd138517: dataIn1 = 32'd1803
; 
32'd138518: dataIn1 = 32'd2962
; 
32'd138519: dataIn1 = 32'd2963
; 
32'd138520: dataIn1 = 32'd2964
; 
32'd138521: dataIn1 = 32'd3320
; 
32'd138522: dataIn1 = 32'd11147
; 
32'd138523: dataIn1 = 32'd11148
; 
32'd138524: dataIn1 = 32'd185
; 
32'd138525: dataIn1 = 32'd1804
; 
32'd138526: dataIn1 = 32'd2963
; 
32'd138527: dataIn1 = 32'd2965
; 
32'd138528: dataIn1 = 32'd2966
; 
32'd138529: dataIn1 = 32'd3322
; 
32'd138530: dataIn1 = 32'd3326
; 
32'd138531: dataIn1 = 32'd185
; 
32'd138532: dataIn1 = 32'd1803
; 
32'd138533: dataIn1 = 32'd2963
; 
32'd138534: dataIn1 = 32'd2965
; 
32'd138535: dataIn1 = 32'd2966
; 
32'd138536: dataIn1 = 32'd3315
; 
32'd138537: dataIn1 = 32'd3318
; 
32'd138538: dataIn1 = 32'd1805
; 
32'd138539: dataIn1 = 32'd1806
; 
32'd138540: dataIn1 = 32'd2967
; 
32'd138541: dataIn1 = 32'd2968
; 
32'd138542: dataIn1 = 32'd2969
; 
32'd138543: dataIn1 = 32'd2970
; 
32'd138544: dataIn1 = 32'd2971
; 
32'd138545: dataIn1 = 32'd1806
; 
32'd138546: dataIn1 = 32'd2967
; 
32'd138547: dataIn1 = 32'd2968
; 
32'd138548: dataIn1 = 32'd2969
; 
32'd138549: dataIn1 = 32'd3332
; 
32'd138550: dataIn1 = 32'd11139
; 
32'd138551: dataIn1 = 32'd11140
; 
32'd138552: dataIn1 = 32'd1805
; 
32'd138553: dataIn1 = 32'd2967
; 
32'd138554: dataIn1 = 32'd2968
; 
32'd138555: dataIn1 = 32'd2969
; 
32'd138556: dataIn1 = 32'd3304
; 
32'd138557: dataIn1 = 32'd11138
; 
32'd138558: dataIn1 = 32'd11139
; 
32'd138559: dataIn1 = 32'd183
; 
32'd138560: dataIn1 = 32'd1806
; 
32'd138561: dataIn1 = 32'd2967
; 
32'd138562: dataIn1 = 32'd2970
; 
32'd138563: dataIn1 = 32'd2971
; 
32'd138564: dataIn1 = 32'd3328
; 
32'd138565: dataIn1 = 32'd3331
; 
32'd138566: dataIn1 = 32'd183
; 
32'd138567: dataIn1 = 32'd1805
; 
32'd138568: dataIn1 = 32'd2967
; 
32'd138569: dataIn1 = 32'd2970
; 
32'd138570: dataIn1 = 32'd2971
; 
32'd138571: dataIn1 = 32'd3302
; 
32'd138572: dataIn1 = 32'd3306
; 
32'd138573: dataIn1 = 32'd1808
; 
32'd138574: dataIn1 = 32'd2972
; 
32'd138575: dataIn1 = 32'd2973
; 
32'd138576: dataIn1 = 32'd2974
; 
32'd138577: dataIn1 = 32'd3338
; 
32'd138578: dataIn1 = 32'd11158
; 
32'd138579: dataIn1 = 32'd11159
; 
32'd138580: dataIn1 = 32'd1807
; 
32'd138581: dataIn1 = 32'd1808
; 
32'd138582: dataIn1 = 32'd2972
; 
32'd138583: dataIn1 = 32'd2973
; 
32'd138584: dataIn1 = 32'd2974
; 
32'd138585: dataIn1 = 32'd2975
; 
32'd138586: dataIn1 = 32'd2976
; 
32'd138587: dataIn1 = 32'd1807
; 
32'd138588: dataIn1 = 32'd2972
; 
32'd138589: dataIn1 = 32'd2973
; 
32'd138590: dataIn1 = 32'd2974
; 
32'd138591: dataIn1 = 32'd3348
; 
32'd138592: dataIn1 = 32'd11159
; 
32'd138593: dataIn1 = 32'd11160
; 
32'd138594: dataIn1 = 32'd366
; 
32'd138595: dataIn1 = 32'd1808
; 
32'd138596: dataIn1 = 32'd2973
; 
32'd138597: dataIn1 = 32'd2975
; 
32'd138598: dataIn1 = 32'd2976
; 
32'd138599: dataIn1 = 32'd3336
; 
32'd138600: dataIn1 = 32'd3340
; 
32'd138601: dataIn1 = 32'd366
; 
32'd138602: dataIn1 = 32'd1807
; 
32'd138603: dataIn1 = 32'd2973
; 
32'd138604: dataIn1 = 32'd2975
; 
32'd138605: dataIn1 = 32'd2976
; 
32'd138606: dataIn1 = 32'd3343
; 
32'd138607: dataIn1 = 32'd3346
; 
32'd138608: dataIn1 = 32'd1810
; 
32'd138609: dataIn1 = 32'd2977
; 
32'd138610: dataIn1 = 32'd2978
; 
32'd138611: dataIn1 = 32'd2979
; 
32'd138612: dataIn1 = 32'd3339
; 
32'd138613: dataIn1 = 32'd11155
; 
32'd138614: dataIn1 = 32'd11156
; 
32'd138615: dataIn1 = 32'd1809
; 
32'd138616: dataIn1 = 32'd2977
; 
32'd138617: dataIn1 = 32'd2978
; 
32'd138618: dataIn1 = 32'd2979
; 
32'd138619: dataIn1 = 32'd3312
; 
32'd138620: dataIn1 = 32'd11154
; 
32'd138621: dataIn1 = 32'd11155
; 
32'd138622: dataIn1 = 32'd1809
; 
32'd138623: dataIn1 = 32'd1810
; 
32'd138624: dataIn1 = 32'd2977
; 
32'd138625: dataIn1 = 32'd2978
; 
32'd138626: dataIn1 = 32'd2979
; 
32'd138627: dataIn1 = 32'd2980
; 
32'd138628: dataIn1 = 32'd2981
; 
32'd138629: dataIn1 = 32'd186
; 
32'd138630: dataIn1 = 32'd1810
; 
32'd138631: dataIn1 = 32'd2979
; 
32'd138632: dataIn1 = 32'd2980
; 
32'd138633: dataIn1 = 32'd2981
; 
32'd138634: dataIn1 = 32'd3337
; 
32'd138635: dataIn1 = 32'd3341
; 
32'd138636: dataIn1 = 32'd186
; 
32'd138637: dataIn1 = 32'd1809
; 
32'd138638: dataIn1 = 32'd2979
; 
32'd138639: dataIn1 = 32'd2980
; 
32'd138640: dataIn1 = 32'd2981
; 
32'd138641: dataIn1 = 32'd3309
; 
32'd138642: dataIn1 = 32'd3313
; 
32'd138643: dataIn1 = 32'd1811
; 
32'd138644: dataIn1 = 32'd1812
; 
32'd138645: dataIn1 = 32'd2982
; 
32'd138646: dataIn1 = 32'd2983
; 
32'd138647: dataIn1 = 32'd2984
; 
32'd138648: dataIn1 = 32'd2985
; 
32'd138649: dataIn1 = 32'd2986
; 
32'd138650: dataIn1 = 32'd1812
; 
32'd138651: dataIn1 = 32'd2982
; 
32'd138652: dataIn1 = 32'd2983
; 
32'd138653: dataIn1 = 32'd2984
; 
32'd138654: dataIn1 = 32'd3354
; 
32'd138655: dataIn1 = 32'd11163
; 
32'd138656: dataIn1 = 32'd11164
; 
32'd138657: dataIn1 = 32'd1811
; 
32'd138658: dataIn1 = 32'd2982
; 
32'd138659: dataIn1 = 32'd2983
; 
32'd138660: dataIn1 = 32'd2984
; 
32'd138661: dataIn1 = 32'd3347
; 
32'd138662: dataIn1 = 32'd11162
; 
32'd138663: dataIn1 = 32'd11163
; 
32'd138664: dataIn1 = 32'd187
; 
32'd138665: dataIn1 = 32'd1812
; 
32'd138666: dataIn1 = 32'd2982
; 
32'd138667: dataIn1 = 32'd2985
; 
32'd138668: dataIn1 = 32'd2986
; 
32'd138669: dataIn1 = 32'd3349
; 
32'd138670: dataIn1 = 32'd3352
; 
32'd138671: dataIn1 = 32'd187
; 
32'd138672: dataIn1 = 32'd1811
; 
32'd138673: dataIn1 = 32'd2982
; 
32'd138674: dataIn1 = 32'd2985
; 
32'd138675: dataIn1 = 32'd2986
; 
32'd138676: dataIn1 = 32'd3342
; 
32'd138677: dataIn1 = 32'd3345
; 
32'd138678: dataIn1 = 32'd1814
; 
32'd138679: dataIn1 = 32'd2987
; 
32'd138680: dataIn1 = 32'd2988
; 
32'd138681: dataIn1 = 32'd2989
; 
32'd138682: dataIn1 = 32'd3359
; 
32'd138683: dataIn1 = 32'd11167
; 
32'd138684: dataIn1 = 32'd11168
; 
32'd138685: dataIn1 = 32'd1813
; 
32'd138686: dataIn1 = 32'd1814
; 
32'd138687: dataIn1 = 32'd2987
; 
32'd138688: dataIn1 = 32'd2988
; 
32'd138689: dataIn1 = 32'd2989
; 
32'd138690: dataIn1 = 32'd2990
; 
32'd138691: dataIn1 = 32'd2991
; 
32'd138692: dataIn1 = 32'd1813
; 
32'd138693: dataIn1 = 32'd2987
; 
32'd138694: dataIn1 = 32'd2988
; 
32'd138695: dataIn1 = 32'd2989
; 
32'd138696: dataIn1 = 32'd3355
; 
32'd138697: dataIn1 = 32'd11166
; 
32'd138698: dataIn1 = 32'd11167
; 
32'd138699: dataIn1 = 32'd373
; 
32'd138700: dataIn1 = 32'd1814
; 
32'd138701: dataIn1 = 32'd2988
; 
32'd138702: dataIn1 = 32'd2990
; 
32'd138703: dataIn1 = 32'd2991
; 
32'd138704: dataIn1 = 32'd3357
; 
32'd138705: dataIn1 = 32'd3361
; 
32'd138706: dataIn1 = 32'd373
; 
32'd138707: dataIn1 = 32'd1813
; 
32'd138708: dataIn1 = 32'd2988
; 
32'd138709: dataIn1 = 32'd2990
; 
32'd138710: dataIn1 = 32'd2991
; 
32'd138711: dataIn1 = 32'd3350
; 
32'd138712: dataIn1 = 32'd3353
; 
32'd138713: dataIn1 = 32'd1815
; 
32'd138714: dataIn1 = 32'd1816
; 
32'd138715: dataIn1 = 32'd2992
; 
32'd138716: dataIn1 = 32'd2993
; 
32'd138717: dataIn1 = 32'd2994
; 
32'd138718: dataIn1 = 32'd2995
; 
32'd138719: dataIn1 = 32'd2996
; 
32'd138720: dataIn1 = 32'd1816
; 
32'd138721: dataIn1 = 32'd2992
; 
32'd138722: dataIn1 = 32'd2993
; 
32'd138723: dataIn1 = 32'd2994
; 
32'd138724: dataIn1 = 32'd3367
; 
32'd138725: dataIn1 = 32'd11184
; 
32'd138726: dataIn1 = 32'd11185
; 
32'd138727: dataIn1 = 32'd1815
; 
32'd138728: dataIn1 = 32'd2992
; 
32'd138729: dataIn1 = 32'd2993
; 
32'd138730: dataIn1 = 32'd2994
; 
32'd138731: dataIn1 = 32'd3375
; 
32'd138732: dataIn1 = 32'd11183
; 
32'd138733: dataIn1 = 32'd11184
; 
32'd138734: dataIn1 = 32'd375
; 
32'd138735: dataIn1 = 32'd1816
; 
32'd138736: dataIn1 = 32'd2992
; 
32'd138737: dataIn1 = 32'd2995
; 
32'd138738: dataIn1 = 32'd2996
; 
32'd138739: dataIn1 = 32'd3363
; 
32'd138740: dataIn1 = 32'd3366
; 
32'd138741: dataIn1 = 32'd375
; 
32'd138742: dataIn1 = 32'd1815
; 
32'd138743: dataIn1 = 32'd2992
; 
32'd138744: dataIn1 = 32'd2995
; 
32'd138745: dataIn1 = 32'd2996
; 
32'd138746: dataIn1 = 32'd3370
; 
32'd138747: dataIn1 = 32'd3373
; 
32'd138748: dataIn1 = 32'd1818
; 
32'd138749: dataIn1 = 32'd2997
; 
32'd138750: dataIn1 = 32'd2998
; 
32'd138751: dataIn1 = 32'd2999
; 
32'd138752: dataIn1 = 32'd3381
; 
32'd138753: dataIn1 = 32'd11175
; 
32'd138754: dataIn1 = 32'd11176
; 
32'd138755: dataIn1 = 32'd1817
; 
32'd138756: dataIn1 = 32'd2997
; 
32'd138757: dataIn1 = 32'd2998
; 
32'd138758: dataIn1 = 32'd2999
; 
32'd138759: dataIn1 = 32'd3389
; 
32'd138760: dataIn1 = 32'd11174
; 
32'd138761: dataIn1 = 32'd11175
; 
32'd138762: dataIn1 = 32'd1817
; 
32'd138763: dataIn1 = 32'd1818
; 
32'd138764: dataIn1 = 32'd2997
; 
32'd138765: dataIn1 = 32'd2998
; 
32'd138766: dataIn1 = 32'd2999
; 
32'd138767: dataIn1 = 32'd3000
; 
32'd138768: dataIn1 = 32'd3001
; 
32'd138769: dataIn1 = 32'd381
; 
32'd138770: dataIn1 = 32'd1818
; 
32'd138771: dataIn1 = 32'd2999
; 
32'd138772: dataIn1 = 32'd3000
; 
32'd138773: dataIn1 = 32'd3001
; 
32'd138774: dataIn1 = 32'd3379
; 
32'd138775: dataIn1 = 32'd3383
; 
32'd138776: dataIn1 = 32'd381
; 
32'd138777: dataIn1 = 32'd1817
; 
32'd138778: dataIn1 = 32'd2999
; 
32'd138779: dataIn1 = 32'd3000
; 
32'd138780: dataIn1 = 32'd3001
; 
32'd138781: dataIn1 = 32'd3386
; 
32'd138782: dataIn1 = 32'd3390
; 
32'd138783: dataIn1 = 32'd1820
; 
32'd138784: dataIn1 = 32'd3002
; 
32'd138785: dataIn1 = 32'd3003
; 
32'd138786: dataIn1 = 32'd3004
; 
32'd138787: dataIn1 = 32'd3380
; 
32'd138788: dataIn1 = 32'd11178
; 
32'd138789: dataIn1 = 32'd11179
; 
32'd138790: dataIn1 = 32'd11180
; 
32'd138791: dataIn1 = 32'd1819
; 
32'd138792: dataIn1 = 32'd1820
; 
32'd138793: dataIn1 = 32'd3002
; 
32'd138794: dataIn1 = 32'd3003
; 
32'd138795: dataIn1 = 32'd3004
; 
32'd138796: dataIn1 = 32'd3005
; 
32'd138797: dataIn1 = 32'd3006
; 
32'd138798: dataIn1 = 32'd1819
; 
32'd138799: dataIn1 = 32'd3002
; 
32'd138800: dataIn1 = 32'd3003
; 
32'd138801: dataIn1 = 32'd3004
; 
32'd138802: dataIn1 = 32'd3376
; 
32'd138803: dataIn1 = 32'd11180
; 
32'd138804: dataIn1 = 32'd11181
; 
32'd138805: dataIn1 = 32'd191
; 
32'd138806: dataIn1 = 32'd1820
; 
32'd138807: dataIn1 = 32'd3003
; 
32'd138808: dataIn1 = 32'd3005
; 
32'd138809: dataIn1 = 32'd3006
; 
32'd138810: dataIn1 = 32'd3378
; 
32'd138811: dataIn1 = 32'd3382
; 
32'd138812: dataIn1 = 32'd191
; 
32'd138813: dataIn1 = 32'd1819
; 
32'd138814: dataIn1 = 32'd3003
; 
32'd138815: dataIn1 = 32'd3005
; 
32'd138816: dataIn1 = 32'd3006
; 
32'd138817: dataIn1 = 32'd3371
; 
32'd138818: dataIn1 = 32'd3374
; 
32'd138819: dataIn1 = 32'd1821
; 
32'd138820: dataIn1 = 32'd1822
; 
32'd138821: dataIn1 = 32'd3007
; 
32'd138822: dataIn1 = 32'd3008
; 
32'd138823: dataIn1 = 32'd3009
; 
32'd138824: dataIn1 = 32'd3010
; 
32'd138825: dataIn1 = 32'd3011
; 
32'd138826: dataIn1 = 32'd1822
; 
32'd138827: dataIn1 = 32'd3007
; 
32'd138828: dataIn1 = 32'd3008
; 
32'd138829: dataIn1 = 32'd3009
; 
32'd138830: dataIn1 = 32'd3388
; 
32'd138831: dataIn1 = 32'd11172
; 
32'd138832: dataIn1 = 32'd1821
; 
32'd138833: dataIn1 = 32'd3007
; 
32'd138834: dataIn1 = 32'd3008
; 
32'd138835: dataIn1 = 32'd3009
; 
32'd138836: dataIn1 = 32'd3360
; 
32'd138837: dataIn1 = 32'd11171
; 
32'd138838: dataIn1 = 32'd11172
; 
32'd138839: dataIn1 = 32'd189
; 
32'd138840: dataIn1 = 32'd1822
; 
32'd138841: dataIn1 = 32'd3007
; 
32'd138842: dataIn1 = 32'd3010
; 
32'd138843: dataIn1 = 32'd3011
; 
32'd138844: dataIn1 = 32'd3384
; 
32'd138845: dataIn1 = 32'd3387
; 
32'd138846: dataIn1 = 32'd189
; 
32'd138847: dataIn1 = 32'd1821
; 
32'd138848: dataIn1 = 32'd3007
; 
32'd138849: dataIn1 = 32'd3010
; 
32'd138850: dataIn1 = 32'd3011
; 
32'd138851: dataIn1 = 32'd3358
; 
32'd138852: dataIn1 = 32'd3362
; 
32'd138853: dataIn1 = 32'd1824
; 
32'd138854: dataIn1 = 32'd3012
; 
32'd138855: dataIn1 = 32'd3013
; 
32'd138856: dataIn1 = 32'd3014
; 
32'd138857: dataIn1 = 32'd3394
; 
32'd138858: dataIn1 = 32'd11191
; 
32'd138859: dataIn1 = 32'd11192
; 
32'd138860: dataIn1 = 32'd1823
; 
32'd138861: dataIn1 = 32'd1824
; 
32'd138862: dataIn1 = 32'd3012
; 
32'd138863: dataIn1 = 32'd3013
; 
32'd138864: dataIn1 = 32'd3014
; 
32'd138865: dataIn1 = 32'd3015
; 
32'd138866: dataIn1 = 32'd3016
; 
32'd138867: dataIn1 = 32'd1823
; 
32'd138868: dataIn1 = 32'd3012
; 
32'd138869: dataIn1 = 32'd3013
; 
32'd138870: dataIn1 = 32'd3014
; 
32'd138871: dataIn1 = 32'd3404
; 
32'd138872: dataIn1 = 32'd11192
; 
32'd138873: dataIn1 = 32'd11193
; 
32'd138874: dataIn1 = 32'd382
; 
32'd138875: dataIn1 = 32'd1824
; 
32'd138876: dataIn1 = 32'd3013
; 
32'd138877: dataIn1 = 32'd3015
; 
32'd138878: dataIn1 = 32'd3016
; 
32'd138879: dataIn1 = 32'd3392
; 
32'd138880: dataIn1 = 32'd3396
; 
32'd138881: dataIn1 = 32'd382
; 
32'd138882: dataIn1 = 32'd1823
; 
32'd138883: dataIn1 = 32'd3013
; 
32'd138884: dataIn1 = 32'd3015
; 
32'd138885: dataIn1 = 32'd3016
; 
32'd138886: dataIn1 = 32'd3399
; 
32'd138887: dataIn1 = 32'd3402
; 
32'd138888: dataIn1 = 32'd1826
; 
32'd138889: dataIn1 = 32'd3017
; 
32'd138890: dataIn1 = 32'd3018
; 
32'd138891: dataIn1 = 32'd3019
; 
32'd138892: dataIn1 = 32'd3395
; 
32'd138893: dataIn1 = 32'd11188
; 
32'd138894: dataIn1 = 32'd11189
; 
32'd138895: dataIn1 = 32'd1825
; 
32'd138896: dataIn1 = 32'd3017
; 
32'd138897: dataIn1 = 32'd3018
; 
32'd138898: dataIn1 = 32'd3019
; 
32'd138899: dataIn1 = 32'd3368
; 
32'd138900: dataIn1 = 32'd11187
; 
32'd138901: dataIn1 = 32'd11188
; 
32'd138902: dataIn1 = 32'd1825
; 
32'd138903: dataIn1 = 32'd1826
; 
32'd138904: dataIn1 = 32'd3017
; 
32'd138905: dataIn1 = 32'd3018
; 
32'd138906: dataIn1 = 32'd3019
; 
32'd138907: dataIn1 = 32'd3020
; 
32'd138908: dataIn1 = 32'd3021
; 
32'd138909: dataIn1 = 32'd192
; 
32'd138910: dataIn1 = 32'd1826
; 
32'd138911: dataIn1 = 32'd3019
; 
32'd138912: dataIn1 = 32'd3020
; 
32'd138913: dataIn1 = 32'd3021
; 
32'd138914: dataIn1 = 32'd3393
; 
32'd138915: dataIn1 = 32'd3397
; 
32'd138916: dataIn1 = 32'd192
; 
32'd138917: dataIn1 = 32'd1825
; 
32'd138918: dataIn1 = 32'd3019
; 
32'd138919: dataIn1 = 32'd3020
; 
32'd138920: dataIn1 = 32'd3021
; 
32'd138921: dataIn1 = 32'd3365
; 
32'd138922: dataIn1 = 32'd3369
; 
32'd138923: dataIn1 = 32'd1827
; 
32'd138924: dataIn1 = 32'd1828
; 
32'd138925: dataIn1 = 32'd3022
; 
32'd138926: dataIn1 = 32'd3023
; 
32'd138927: dataIn1 = 32'd3024
; 
32'd138928: dataIn1 = 32'd3025
; 
32'd138929: dataIn1 = 32'd3026
; 
32'd138930: dataIn1 = 32'd1828
; 
32'd138931: dataIn1 = 32'd3022
; 
32'd138932: dataIn1 = 32'd3023
; 
32'd138933: dataIn1 = 32'd3024
; 
32'd138934: dataIn1 = 32'd3441
; 
32'd138935: dataIn1 = 32'd11195
; 
32'd138936: dataIn1 = 32'd11196
; 
32'd138937: dataIn1 = 32'd11197
; 
32'd138938: dataIn1 = 32'd1827
; 
32'd138939: dataIn1 = 32'd3022
; 
32'd138940: dataIn1 = 32'd3023
; 
32'd138941: dataIn1 = 32'd3024
; 
32'd138942: dataIn1 = 32'd3403
; 
32'd138943: dataIn1 = 32'd11195
; 
32'd138944: dataIn1 = 32'd193
; 
32'd138945: dataIn1 = 32'd1828
; 
32'd138946: dataIn1 = 32'd3022
; 
32'd138947: dataIn1 = 32'd3025
; 
32'd138948: dataIn1 = 32'd3026
; 
32'd138949: dataIn1 = 32'd193
; 
32'd138950: dataIn1 = 32'd1827
; 
32'd138951: dataIn1 = 32'd3022
; 
32'd138952: dataIn1 = 32'd3025
; 
32'd138953: dataIn1 = 32'd3026
; 
32'd138954: dataIn1 = 32'd3398
; 
32'd138955: dataIn1 = 32'd3401
; 
32'd138956: dataIn1 = 32'd747
; 
32'd138957: dataIn1 = 32'd1425
; 
32'd138958: dataIn1 = 32'd1854
; 
32'd138959: dataIn1 = 32'd3027
; 
32'd138960: dataIn1 = 32'd3028
; 
32'd138961: dataIn1 = 32'd3029
; 
32'd138962: dataIn1 = 32'd3442
; 
32'd138963: dataIn1 = 32'd1853
; 
32'd138964: dataIn1 = 32'd1854
; 
32'd138965: dataIn1 = 32'd3027
; 
32'd138966: dataIn1 = 32'd3028
; 
32'd138967: dataIn1 = 32'd3029
; 
32'd138968: dataIn1 = 32'd3030
; 
32'd138969: dataIn1 = 32'd3031
; 
32'd138970: dataIn1 = 32'd747
; 
32'd138971: dataIn1 = 32'd1426
; 
32'd138972: dataIn1 = 32'd1853
; 
32'd138973: dataIn1 = 32'd3027
; 
32'd138974: dataIn1 = 32'd3028
; 
32'd138975: dataIn1 = 32'd3029
; 
32'd138976: dataIn1 = 32'd3410
; 
32'd138977: dataIn1 = 32'd391
; 
32'd138978: dataIn1 = 32'd1854
; 
32'd138979: dataIn1 = 32'd3028
; 
32'd138980: dataIn1 = 32'd3030
; 
32'd138981: dataIn1 = 32'd3031
; 
32'd138982: dataIn1 = 32'd10256
; 
32'd138983: dataIn1 = 32'd10257
; 
32'd138984: dataIn1 = 32'd391
; 
32'd138985: dataIn1 = 32'd1853
; 
32'd138986: dataIn1 = 32'd3028
; 
32'd138987: dataIn1 = 32'd3030
; 
32'd138988: dataIn1 = 32'd3031
; 
32'd138989: dataIn1 = 32'd3406
; 
32'd138990: dataIn1 = 32'd3408
; 
32'd138991: dataIn1 = 32'd755
; 
32'd138992: dataIn1 = 32'd1439
; 
32'd138993: dataIn1 = 32'd1857
; 
32'd138994: dataIn1 = 32'd3032
; 
32'd138995: dataIn1 = 32'd3033
; 
32'd138996: dataIn1 = 32'd3034
; 
32'd138997: dataIn1 = 32'd3413
; 
32'd138998: dataIn1 = 32'd755
; 
32'd138999: dataIn1 = 32'd1440
; 
32'd139000: dataIn1 = 32'd1856
; 
32'd139001: dataIn1 = 32'd3032
; 
32'd139002: dataIn1 = 32'd3033
; 
32'd139003: dataIn1 = 32'd3034
; 
32'd139004: dataIn1 = 32'd3414
; 
32'd139005: dataIn1 = 32'd393
; 
32'd139006: dataIn1 = 32'd1856
; 
32'd139007: dataIn1 = 32'd1857
; 
32'd139008: dataIn1 = 32'd3032
; 
32'd139009: dataIn1 = 32'd3033
; 
32'd139010: dataIn1 = 32'd3034
; 
32'd139011: dataIn1 = 32'd795
; 
32'd139012: dataIn1 = 32'd1501
; 
32'd139013: dataIn1 = 32'd1869
; 
32'd139014: dataIn1 = 32'd3035
; 
32'd139015: dataIn1 = 32'd3036
; 
32'd139016: dataIn1 = 32'd3037
; 
32'd139017: dataIn1 = 32'd3444
; 
32'd139018: dataIn1 = 32'd795
; 
32'd139019: dataIn1 = 32'd1502
; 
32'd139020: dataIn1 = 32'd1868
; 
32'd139021: dataIn1 = 32'd3035
; 
32'd139022: dataIn1 = 32'd3036
; 
32'd139023: dataIn1 = 32'd3037
; 
32'd139024: dataIn1 = 32'd3443
; 
32'd139025: dataIn1 = 32'd1868
; 
32'd139026: dataIn1 = 32'd1869
; 
32'd139027: dataIn1 = 32'd3035
; 
32'd139028: dataIn1 = 32'd3036
; 
32'd139029: dataIn1 = 32'd3037
; 
32'd139030: dataIn1 = 32'd3038
; 
32'd139031: dataIn1 = 32'd3039
; 
32'd139032: dataIn1 = 32'd980
; 
32'd139033: dataIn1 = 32'd1869
; 
32'd139034: dataIn1 = 32'd3037
; 
32'd139035: dataIn1 = 32'd3038
; 
32'd139036: dataIn1 = 32'd3039
; 
32'd139037: dataIn1 = 32'd3417
; 
32'd139038: dataIn1 = 32'd3418
; 
32'd139039: dataIn1 = 32'd980
; 
32'd139040: dataIn1 = 32'd1868
; 
32'd139041: dataIn1 = 32'd2049
; 
32'd139042: dataIn1 = 32'd3037
; 
32'd139043: dataIn1 = 32'd3038
; 
32'd139044: dataIn1 = 32'd3039
; 
32'd139045: dataIn1 = 32'd414
; 
32'd139046: dataIn1 = 32'd800
; 
32'd139047: dataIn1 = 32'd1872
; 
32'd139048: dataIn1 = 32'd2759
; 
32'd139049: dataIn1 = 32'd3040
; 
32'd139050: dataIn1 = 32'd3440
; 
32'd139051: dataIn1 = 32'd3445
; 
32'd139052: dataIn1 = 32'd1724
; 
32'd139053: dataIn1 = 32'd1977
; 
32'd139054: dataIn1 = 32'd2764
; 
32'd139055: dataIn1 = 32'd3041
; 
32'd139056: dataIn1 = 32'd3042
; 
32'd139057: dataIn1 = 32'd3043
; 
32'd139058: dataIn1 = 32'd3044
; 
32'd139059: dataIn1 = 32'd1724
; 
32'd139060: dataIn1 = 32'd1729
; 
32'd139061: dataIn1 = 32'd3041
; 
32'd139062: dataIn1 = 32'd3042
; 
32'd139063: dataIn1 = 32'd3043
; 
32'd139064: dataIn1 = 32'd3045
; 
32'd139065: dataIn1 = 32'd3046
; 
32'd139066: dataIn1 = 32'd1729
; 
32'd139067: dataIn1 = 32'd1977
; 
32'd139068: dataIn1 = 32'd2781
; 
32'd139069: dataIn1 = 32'd3041
; 
32'd139070: dataIn1 = 32'd3042
; 
32'd139071: dataIn1 = 32'd3043
; 
32'd139072: dataIn1 = 32'd3047
; 
32'd139073: dataIn1 = 32'd279
; 
32'd139074: dataIn1 = 32'd1977
; 
32'd139075: dataIn1 = 32'd2764
; 
32'd139076: dataIn1 = 32'd3041
; 
32'd139077: dataIn1 = 32'd3044
; 
32'd139078: dataIn1 = 32'd3989
; 
32'd139079: dataIn1 = 32'd3998
; 
32'd139080: dataIn1 = 32'd1724
; 
32'd139081: dataIn1 = 32'd2762
; 
32'd139082: dataIn1 = 32'd3042
; 
32'd139083: dataIn1 = 32'd3045
; 
32'd139084: dataIn1 = 32'd3046
; 
32'd139085: dataIn1 = 32'd10992
; 
32'd139086: dataIn1 = 32'd10993
; 
32'd139087: dataIn1 = 32'd1729
; 
32'd139088: dataIn1 = 32'd2778
; 
32'd139089: dataIn1 = 32'd3042
; 
32'd139090: dataIn1 = 32'd3045
; 
32'd139091: dataIn1 = 32'd3046
; 
32'd139092: dataIn1 = 32'd10993
; 
32'd139093: dataIn1 = 32'd10994
; 
32'd139094: dataIn1 = 32'd155
; 
32'd139095: dataIn1 = 32'd1977
; 
32'd139096: dataIn1 = 32'd2781
; 
32'd139097: dataIn1 = 32'd3043
; 
32'd139098: dataIn1 = 32'd3047
; 
32'd139099: dataIn1 = 32'd4000
; 
32'd139100: dataIn1 = 32'd4009
; 
32'd139101: dataIn1 = 32'd1723
; 
32'd139102: dataIn1 = 32'd1978
; 
32'd139103: dataIn1 = 32'd2765
; 
32'd139104: dataIn1 = 32'd3048
; 
32'd139105: dataIn1 = 32'd3049
; 
32'd139106: dataIn1 = 32'd3050
; 
32'd139107: dataIn1 = 32'd3051
; 
32'd139108: dataIn1 = 32'd1725
; 
32'd139109: dataIn1 = 32'd1978
; 
32'd139110: dataIn1 = 32'd2771
; 
32'd139111: dataIn1 = 32'd3048
; 
32'd139112: dataIn1 = 32'd3049
; 
32'd139113: dataIn1 = 32'd3050
; 
32'd139114: dataIn1 = 32'd3052
; 
32'd139115: dataIn1 = 32'd1723
; 
32'd139116: dataIn1 = 32'd1725
; 
32'd139117: dataIn1 = 32'd3048
; 
32'd139118: dataIn1 = 32'd3049
; 
32'd139119: dataIn1 = 32'd3050
; 
32'd139120: dataIn1 = 32'd3053
; 
32'd139121: dataIn1 = 32'd3054
; 
32'd139122: dataIn1 = 32'd279
; 
32'd139123: dataIn1 = 32'd1978
; 
32'd139124: dataIn1 = 32'd2765
; 
32'd139125: dataIn1 = 32'd3048
; 
32'd139126: dataIn1 = 32'd3051
; 
32'd139127: dataIn1 = 32'd3990
; 
32'd139128: dataIn1 = 32'd3995
; 
32'd139129: dataIn1 = 32'd154
; 
32'd139130: dataIn1 = 32'd1978
; 
32'd139131: dataIn1 = 32'd2771
; 
32'd139132: dataIn1 = 32'd3049
; 
32'd139133: dataIn1 = 32'd3052
; 
32'd139134: dataIn1 = 32'd3960
; 
32'd139135: dataIn1 = 32'd3996
; 
32'd139136: dataIn1 = 32'd1723
; 
32'd139137: dataIn1 = 32'd2763
; 
32'd139138: dataIn1 = 32'd3050
; 
32'd139139: dataIn1 = 32'd3053
; 
32'd139140: dataIn1 = 32'd3054
; 
32'd139141: dataIn1 = 32'd10989
; 
32'd139142: dataIn1 = 32'd10990
; 
32'd139143: dataIn1 = 32'd1299
; 
32'd139144: dataIn1 = 32'd1725
; 
32'd139145: dataIn1 = 32'd2768
; 
32'd139146: dataIn1 = 32'd3050
; 
32'd139147: dataIn1 = 32'd3053
; 
32'd139148: dataIn1 = 32'd3054
; 
32'd139149: dataIn1 = 32'd10989
; 
32'd139150: dataIn1 = 32'd1728
; 
32'd139151: dataIn1 = 32'd1730
; 
32'd139152: dataIn1 = 32'd3055
; 
32'd139153: dataIn1 = 32'd3056
; 
32'd139154: dataIn1 = 32'd3057
; 
32'd139155: dataIn1 = 32'd3058
; 
32'd139156: dataIn1 = 32'd3059
; 
32'd139157: dataIn1 = 32'd1728
; 
32'd139158: dataIn1 = 32'd1979
; 
32'd139159: dataIn1 = 32'd2775
; 
32'd139160: dataIn1 = 32'd3055
; 
32'd139161: dataIn1 = 32'd3056
; 
32'd139162: dataIn1 = 32'd3057
; 
32'd139163: dataIn1 = 32'd3060
; 
32'd139164: dataIn1 = 32'd1730
; 
32'd139165: dataIn1 = 32'd1979
; 
32'd139166: dataIn1 = 32'd2780
; 
32'd139167: dataIn1 = 32'd3055
; 
32'd139168: dataIn1 = 32'd3056
; 
32'd139169: dataIn1 = 32'd3057
; 
32'd139170: dataIn1 = 32'd3061
; 
32'd139171: dataIn1 = 32'd1728
; 
32'd139172: dataIn1 = 32'd2772
; 
32'd139173: dataIn1 = 32'd3055
; 
32'd139174: dataIn1 = 32'd3058
; 
32'd139175: dataIn1 = 32'd3059
; 
32'd139176: dataIn1 = 32'd10997
; 
32'd139177: dataIn1 = 32'd10998
; 
32'd139178: dataIn1 = 32'd1730
; 
32'd139179: dataIn1 = 32'd2777
; 
32'd139180: dataIn1 = 32'd3055
; 
32'd139181: dataIn1 = 32'd3058
; 
32'd139182: dataIn1 = 32'd3059
; 
32'd139183: dataIn1 = 32'd10996
; 
32'd139184: dataIn1 = 32'd10997
; 
32'd139185: dataIn1 = 32'd286
; 
32'd139186: dataIn1 = 32'd1979
; 
32'd139187: dataIn1 = 32'd2775
; 
32'd139188: dataIn1 = 32'd3056
; 
32'd139189: dataIn1 = 32'd3060
; 
32'd139190: dataIn1 = 32'd4015
; 
32'd139191: dataIn1 = 32'd4024
; 
32'd139192: dataIn1 = 32'd155
; 
32'd139193: dataIn1 = 32'd1979
; 
32'd139194: dataIn1 = 32'd2780
; 
32'd139195: dataIn1 = 32'd3057
; 
32'd139196: dataIn1 = 32'd3061
; 
32'd139197: dataIn1 = 32'd4008
; 
32'd139198: dataIn1 = 32'd4025
; 
32'd139199: dataIn1 = 32'd1731
; 
32'd139200: dataIn1 = 32'd1980
; 
32'd139201: dataIn1 = 32'd2786
; 
32'd139202: dataIn1 = 32'd3062
; 
32'd139203: dataIn1 = 32'd3063
; 
32'd139204: dataIn1 = 32'd3064
; 
32'd139205: dataIn1 = 32'd3065
; 
32'd139206: dataIn1 = 32'd1727
; 
32'd139207: dataIn1 = 32'd1980
; 
32'd139208: dataIn1 = 32'd2776
; 
32'd139209: dataIn1 = 32'd3062
; 
32'd139210: dataIn1 = 32'd3063
; 
32'd139211: dataIn1 = 32'd3064
; 
32'd139212: dataIn1 = 32'd3066
; 
32'd139213: dataIn1 = 32'd1727
; 
32'd139214: dataIn1 = 32'd1731
; 
32'd139215: dataIn1 = 32'd3062
; 
32'd139216: dataIn1 = 32'd3063
; 
32'd139217: dataIn1 = 32'd3064
; 
32'd139218: dataIn1 = 32'd3067
; 
32'd139219: dataIn1 = 32'd3068
; 
32'd139220: dataIn1 = 32'd157
; 
32'd139221: dataIn1 = 32'd1980
; 
32'd139222: dataIn1 = 32'd2786
; 
32'd139223: dataIn1 = 32'd3062
; 
32'd139224: dataIn1 = 32'd3065
; 
32'd139225: dataIn1 = 32'd4019
; 
32'd139226: dataIn1 = 32'd4029
; 
32'd139227: dataIn1 = 32'd286
; 
32'd139228: dataIn1 = 32'd1980
; 
32'd139229: dataIn1 = 32'd2776
; 
32'd139230: dataIn1 = 32'd3063
; 
32'd139231: dataIn1 = 32'd3066
; 
32'd139232: dataIn1 = 32'd4016
; 
32'd139233: dataIn1 = 32'd4020
; 
32'd139234: dataIn1 = 32'd1731
; 
32'd139235: dataIn1 = 32'd2784
; 
32'd139236: dataIn1 = 32'd3064
; 
32'd139237: dataIn1 = 32'd3067
; 
32'd139238: dataIn1 = 32'd3068
; 
32'd139239: dataIn1 = 32'd11001
; 
32'd139240: dataIn1 = 32'd11002
; 
32'd139241: dataIn1 = 32'd1727
; 
32'd139242: dataIn1 = 32'd2774
; 
32'd139243: dataIn1 = 32'd3064
; 
32'd139244: dataIn1 = 32'd3067
; 
32'd139245: dataIn1 = 32'd3068
; 
32'd139246: dataIn1 = 32'd11000
; 
32'd139247: dataIn1 = 32'd11001
; 
32'd139248: dataIn1 = 32'd1732
; 
32'd139249: dataIn1 = 32'd1981
; 
32'd139250: dataIn1 = 32'd2785
; 
32'd139251: dataIn1 = 32'd3069
; 
32'd139252: dataIn1 = 32'd3070
; 
32'd139253: dataIn1 = 32'd3071
; 
32'd139254: dataIn1 = 32'd3072
; 
32'd139255: dataIn1 = 32'd1733
; 
32'd139256: dataIn1 = 32'd1981
; 
32'd139257: dataIn1 = 32'd2791
; 
32'd139258: dataIn1 = 32'd3069
; 
32'd139259: dataIn1 = 32'd3070
; 
32'd139260: dataIn1 = 32'd3071
; 
32'd139261: dataIn1 = 32'd3073
; 
32'd139262: dataIn1 = 32'd1732
; 
32'd139263: dataIn1 = 32'd1733
; 
32'd139264: dataIn1 = 32'd3069
; 
32'd139265: dataIn1 = 32'd3070
; 
32'd139266: dataIn1 = 32'd3071
; 
32'd139267: dataIn1 = 32'd3074
; 
32'd139268: dataIn1 = 32'd3075
; 
32'd139269: dataIn1 = 32'd157
; 
32'd139270: dataIn1 = 32'd1981
; 
32'd139271: dataIn1 = 32'd2785
; 
32'd139272: dataIn1 = 32'd3069
; 
32'd139273: dataIn1 = 32'd3072
; 
32'd139274: dataIn1 = 32'd4030
; 
32'd139275: dataIn1 = 32'd4043
; 
32'd139276: dataIn1 = 32'd293
; 
32'd139277: dataIn1 = 32'd1981
; 
32'd139278: dataIn1 = 32'd2791
; 
32'd139279: dataIn1 = 32'd3070
; 
32'd139280: dataIn1 = 32'd3073
; 
32'd139281: dataIn1 = 32'd4040
; 
32'd139282: dataIn1 = 32'd4044
; 
32'd139283: dataIn1 = 32'd1732
; 
32'd139284: dataIn1 = 32'd2783
; 
32'd139285: dataIn1 = 32'd3071
; 
32'd139286: dataIn1 = 32'd3074
; 
32'd139287: dataIn1 = 32'd3075
; 
32'd139288: dataIn1 = 32'd11004
; 
32'd139289: dataIn1 = 32'd11005
; 
32'd139290: dataIn1 = 32'd1733
; 
32'd139291: dataIn1 = 32'd2789
; 
32'd139292: dataIn1 = 32'd3071
; 
32'd139293: dataIn1 = 32'd3074
; 
32'd139294: dataIn1 = 32'd3075
; 
32'd139295: dataIn1 = 32'd11005
; 
32'd139296: dataIn1 = 32'd11006
; 
32'd139297: dataIn1 = 32'd1734
; 
32'd139298: dataIn1 = 32'd1741
; 
32'd139299: dataIn1 = 32'd3076
; 
32'd139300: dataIn1 = 32'd3077
; 
32'd139301: dataIn1 = 32'd3078
; 
32'd139302: dataIn1 = 32'd3079
; 
32'd139303: dataIn1 = 32'd3080
; 
32'd139304: dataIn1 = 32'd1734
; 
32'd139305: dataIn1 = 32'd1982
; 
32'd139306: dataIn1 = 32'd2790
; 
32'd139307: dataIn1 = 32'd3076
; 
32'd139308: dataIn1 = 32'd3077
; 
32'd139309: dataIn1 = 32'd3078
; 
32'd139310: dataIn1 = 32'd3081
; 
32'd139311: dataIn1 = 32'd1741
; 
32'd139312: dataIn1 = 32'd1982
; 
32'd139313: dataIn1 = 32'd2811
; 
32'd139314: dataIn1 = 32'd3076
; 
32'd139315: dataIn1 = 32'd3077
; 
32'd139316: dataIn1 = 32'd3078
; 
32'd139317: dataIn1 = 32'd3082
; 
32'd139318: dataIn1 = 32'd1734
; 
32'd139319: dataIn1 = 32'd2787
; 
32'd139320: dataIn1 = 32'd3076
; 
32'd139321: dataIn1 = 32'd3079
; 
32'd139322: dataIn1 = 32'd3080
; 
32'd139323: dataIn1 = 32'd11008
; 
32'd139324: dataIn1 = 32'd11009
; 
32'd139325: dataIn1 = 32'd1741
; 
32'd139326: dataIn1 = 32'd2809
; 
32'd139327: dataIn1 = 32'd3076
; 
32'd139328: dataIn1 = 32'd3079
; 
32'd139329: dataIn1 = 32'd3080
; 
32'd139330: dataIn1 = 32'd11009
; 
32'd139331: dataIn1 = 32'd11010
; 
32'd139332: dataIn1 = 32'd293
; 
32'd139333: dataIn1 = 32'd1982
; 
32'd139334: dataIn1 = 32'd2790
; 
32'd139335: dataIn1 = 32'd3077
; 
32'd139336: dataIn1 = 32'd3081
; 
32'd139337: dataIn1 = 32'd4039
; 
32'd139338: dataIn1 = 32'd4047
; 
32'd139339: dataIn1 = 32'd159
; 
32'd139340: dataIn1 = 32'd1982
; 
32'd139341: dataIn1 = 32'd2811
; 
32'd139342: dataIn1 = 32'd3078
; 
32'd139343: dataIn1 = 32'd3082
; 
32'd139344: dataIn1 = 32'd4048
; 
32'd139345: dataIn1 = 32'd4056
; 
32'd139346: dataIn1 = 32'd1736
; 
32'd139347: dataIn1 = 32'd1983
; 
32'd139348: dataIn1 = 32'd2795
; 
32'd139349: dataIn1 = 32'd3083
; 
32'd139350: dataIn1 = 32'd3084
; 
32'd139351: dataIn1 = 32'd3085
; 
32'd139352: dataIn1 = 32'd3086
; 
32'd139353: dataIn1 = 32'd1736
; 
32'd139354: dataIn1 = 32'd1745
; 
32'd139355: dataIn1 = 32'd3083
; 
32'd139356: dataIn1 = 32'd3084
; 
32'd139357: dataIn1 = 32'd3085
; 
32'd139358: dataIn1 = 32'd3087
; 
32'd139359: dataIn1 = 32'd3088
; 
32'd139360: dataIn1 = 32'd1745
; 
32'd139361: dataIn1 = 32'd1983
; 
32'd139362: dataIn1 = 32'd2821
; 
32'd139363: dataIn1 = 32'd3083
; 
32'd139364: dataIn1 = 32'd3084
; 
32'd139365: dataIn1 = 32'd3085
; 
32'd139366: dataIn1 = 32'd3089
; 
32'd139367: dataIn1 = 32'd295
; 
32'd139368: dataIn1 = 32'd1983
; 
32'd139369: dataIn1 = 32'd2795
; 
32'd139370: dataIn1 = 32'd3083
; 
32'd139371: dataIn1 = 32'd3086
; 
32'd139372: dataIn1 = 32'd4085
; 
32'd139373: dataIn1 = 32'd4094
; 
32'd139374: dataIn1 = 32'd1736
; 
32'd139375: dataIn1 = 32'd2793
; 
32'd139376: dataIn1 = 32'd3084
; 
32'd139377: dataIn1 = 32'd3087
; 
32'd139378: dataIn1 = 32'd3088
; 
32'd139379: dataIn1 = 32'd11024
; 
32'd139380: dataIn1 = 32'd11025
; 
32'd139381: dataIn1 = 32'd1745
; 
32'd139382: dataIn1 = 32'd2818
; 
32'd139383: dataIn1 = 32'd3084
; 
32'd139384: dataIn1 = 32'd3087
; 
32'd139385: dataIn1 = 32'd3088
; 
32'd139386: dataIn1 = 32'd11025
; 
32'd139387: dataIn1 = 32'd11026
; 
32'd139388: dataIn1 = 32'd162
; 
32'd139389: dataIn1 = 32'd1983
; 
32'd139390: dataIn1 = 32'd2821
; 
32'd139391: dataIn1 = 32'd3085
; 
32'd139392: dataIn1 = 32'd3089
; 
32'd139393: dataIn1 = 32'd4096
; 
32'd139394: dataIn1 = 32'd4105
; 
32'd139395: dataIn1 = 32'd1735
; 
32'd139396: dataIn1 = 32'd1984
; 
32'd139397: dataIn1 = 32'd2796
; 
32'd139398: dataIn1 = 32'd3090
; 
32'd139399: dataIn1 = 32'd3091
; 
32'd139400: dataIn1 = 32'd3092
; 
32'd139401: dataIn1 = 32'd3093
; 
32'd139402: dataIn1 = 32'd1739
; 
32'd139403: dataIn1 = 32'd1984
; 
32'd139404: dataIn1 = 32'd2806
; 
32'd139405: dataIn1 = 32'd3090
; 
32'd139406: dataIn1 = 32'd3091
; 
32'd139407: dataIn1 = 32'd3092
; 
32'd139408: dataIn1 = 32'd3094
; 
32'd139409: dataIn1 = 32'd1735
; 
32'd139410: dataIn1 = 32'd1739
; 
32'd139411: dataIn1 = 32'd3090
; 
32'd139412: dataIn1 = 32'd3091
; 
32'd139413: dataIn1 = 32'd3092
; 
32'd139414: dataIn1 = 32'd3095
; 
32'd139415: dataIn1 = 32'd3096
; 
32'd139416: dataIn1 = 32'd295
; 
32'd139417: dataIn1 = 32'd1984
; 
32'd139418: dataIn1 = 32'd2796
; 
32'd139419: dataIn1 = 32'd3090
; 
32'd139420: dataIn1 = 32'd3093
; 
32'd139421: dataIn1 = 32'd4086
; 
32'd139422: dataIn1 = 32'd4091
; 
32'd139423: dataIn1 = 32'd161
; 
32'd139424: dataIn1 = 32'd1984
; 
32'd139425: dataIn1 = 32'd2806
; 
32'd139426: dataIn1 = 32'd3091
; 
32'd139427: dataIn1 = 32'd3094
; 
32'd139428: dataIn1 = 32'd4079
; 
32'd139429: dataIn1 = 32'd4092
; 
32'd139430: dataIn1 = 32'd1735
; 
32'd139431: dataIn1 = 32'd2794
; 
32'd139432: dataIn1 = 32'd3092
; 
32'd139433: dataIn1 = 32'd3095
; 
32'd139434: dataIn1 = 32'd3096
; 
32'd139435: dataIn1 = 32'd11021
; 
32'd139436: dataIn1 = 32'd11022
; 
32'd139437: dataIn1 = 32'd1739
; 
32'd139438: dataIn1 = 32'd2804
; 
32'd139439: dataIn1 = 32'd3092
; 
32'd139440: dataIn1 = 32'd3095
; 
32'd139441: dataIn1 = 32'd3096
; 
32'd139442: dataIn1 = 32'd11020
; 
32'd139443: dataIn1 = 32'd11021
; 
32'd139444: dataIn1 = 32'd1738
; 
32'd139445: dataIn1 = 32'd1740
; 
32'd139446: dataIn1 = 32'd3097
; 
32'd139447: dataIn1 = 32'd3098
; 
32'd139448: dataIn1 = 32'd3099
; 
32'd139449: dataIn1 = 32'd3100
; 
32'd139450: dataIn1 = 32'd3101
; 
32'd139451: dataIn1 = 32'd1740
; 
32'd139452: dataIn1 = 32'd1985
; 
32'd139453: dataIn1 = 32'd2805
; 
32'd139454: dataIn1 = 32'd3097
; 
32'd139455: dataIn1 = 32'd3098
; 
32'd139456: dataIn1 = 32'd3099
; 
32'd139457: dataIn1 = 32'd3102
; 
32'd139458: dataIn1 = 32'd1738
; 
32'd139459: dataIn1 = 32'd1985
; 
32'd139460: dataIn1 = 32'd2800
; 
32'd139461: dataIn1 = 32'd3097
; 
32'd139462: dataIn1 = 32'd3098
; 
32'd139463: dataIn1 = 32'd3099
; 
32'd139464: dataIn1 = 32'd3103
; 
32'd139465: dataIn1 = 32'd1740
; 
32'd139466: dataIn1 = 32'd2802
; 
32'd139467: dataIn1 = 32'd3097
; 
32'd139468: dataIn1 = 32'd3100
; 
32'd139469: dataIn1 = 32'd3101
; 
32'd139470: dataIn1 = 32'd11017
; 
32'd139471: dataIn1 = 32'd11018
; 
32'd139472: dataIn1 = 32'd1738
; 
32'd139473: dataIn1 = 32'd2797
; 
32'd139474: dataIn1 = 32'd3097
; 
32'd139475: dataIn1 = 32'd3100
; 
32'd139476: dataIn1 = 32'd3101
; 
32'd139477: dataIn1 = 32'd11016
; 
32'd139478: dataIn1 = 32'd11017
; 
32'd139479: dataIn1 = 32'd161
; 
32'd139480: dataIn1 = 32'd1985
; 
32'd139481: dataIn1 = 32'd2805
; 
32'd139482: dataIn1 = 32'd3098
; 
32'd139483: dataIn1 = 32'd3102
; 
32'd139484: dataIn1 = 32'd4071
; 
32'd139485: dataIn1 = 32'd4078
; 
32'd139486: dataIn1 = 32'd301
; 
32'd139487: dataIn1 = 32'd1985
; 
32'd139488: dataIn1 = 32'd2800
; 
32'd139489: dataIn1 = 32'd3099
; 
32'd139490: dataIn1 = 32'd3103
; 
32'd139491: dataIn1 = 32'd4065
; 
32'd139492: dataIn1 = 32'd4072
; 
32'd139493: dataIn1 = 32'd1742
; 
32'd139494: dataIn1 = 32'd1986
; 
32'd139495: dataIn1 = 32'd2810
; 
32'd139496: dataIn1 = 32'd3104
; 
32'd139497: dataIn1 = 32'd3105
; 
32'd139498: dataIn1 = 32'd3106
; 
32'd139499: dataIn1 = 32'd3107
; 
32'd139500: dataIn1 = 32'd1737
; 
32'd139501: dataIn1 = 32'd1742
; 
32'd139502: dataIn1 = 32'd3104
; 
32'd139503: dataIn1 = 32'd3105
; 
32'd139504: dataIn1 = 32'd3106
; 
32'd139505: dataIn1 = 32'd3108
; 
32'd139506: dataIn1 = 32'd3109
; 
32'd139507: dataIn1 = 32'd1737
; 
32'd139508: dataIn1 = 32'd1986
; 
32'd139509: dataIn1 = 32'd2801
; 
32'd139510: dataIn1 = 32'd3104
; 
32'd139511: dataIn1 = 32'd3105
; 
32'd139512: dataIn1 = 32'd3106
; 
32'd139513: dataIn1 = 32'd3110
; 
32'd139514: dataIn1 = 32'd159
; 
32'd139515: dataIn1 = 32'd1986
; 
32'd139516: dataIn1 = 32'd2810
; 
32'd139517: dataIn1 = 32'd3104
; 
32'd139518: dataIn1 = 32'd3107
; 
32'd139519: dataIn1 = 32'd4057
; 
32'd139520: dataIn1 = 32'd4067
; 
32'd139521: dataIn1 = 32'd1742
; 
32'd139522: dataIn1 = 32'd2808
; 
32'd139523: dataIn1 = 32'd3105
; 
32'd139524: dataIn1 = 32'd3108
; 
32'd139525: dataIn1 = 32'd3109
; 
32'd139526: dataIn1 = 32'd11012
; 
32'd139527: dataIn1 = 32'd11013
; 
32'd139528: dataIn1 = 32'd1737
; 
32'd139529: dataIn1 = 32'd2798
; 
32'd139530: dataIn1 = 32'd3105
; 
32'd139531: dataIn1 = 32'd3108
; 
32'd139532: dataIn1 = 32'd3109
; 
32'd139533: dataIn1 = 32'd11013
; 
32'd139534: dataIn1 = 32'd11014
; 
32'd139535: dataIn1 = 32'd301
; 
32'd139536: dataIn1 = 32'd1986
; 
32'd139537: dataIn1 = 32'd2801
; 
32'd139538: dataIn1 = 32'd3106
; 
32'd139539: dataIn1 = 32'd3110
; 
32'd139540: dataIn1 = 32'd4066
; 
32'd139541: dataIn1 = 32'd4069
; 
32'd139542: dataIn1 = 32'd1744
; 
32'd139543: dataIn1 = 32'd1746
; 
32'd139544: dataIn1 = 32'd3111
; 
32'd139545: dataIn1 = 32'd3112
; 
32'd139546: dataIn1 = 32'd3113
; 
32'd139547: dataIn1 = 32'd3114
; 
32'd139548: dataIn1 = 32'd3115
; 
32'd139549: dataIn1 = 32'd1744
; 
32'd139550: dataIn1 = 32'd1987
; 
32'd139551: dataIn1 = 32'd2815
; 
32'd139552: dataIn1 = 32'd3111
; 
32'd139553: dataIn1 = 32'd3112
; 
32'd139554: dataIn1 = 32'd3113
; 
32'd139555: dataIn1 = 32'd3116
; 
32'd139556: dataIn1 = 32'd1746
; 
32'd139557: dataIn1 = 32'd1987
; 
32'd139558: dataIn1 = 32'd2820
; 
32'd139559: dataIn1 = 32'd3111
; 
32'd139560: dataIn1 = 32'd3112
; 
32'd139561: dataIn1 = 32'd3113
; 
32'd139562: dataIn1 = 32'd3117
; 
32'd139563: dataIn1 = 32'd1744
; 
32'd139564: dataIn1 = 32'd2812
; 
32'd139565: dataIn1 = 32'd3111
; 
32'd139566: dataIn1 = 32'd3114
; 
32'd139567: dataIn1 = 32'd3115
; 
32'd139568: dataIn1 = 32'd11029
; 
32'd139569: dataIn1 = 32'd11030
; 
32'd139570: dataIn1 = 32'd1746
; 
32'd139571: dataIn1 = 32'd2817
; 
32'd139572: dataIn1 = 32'd3111
; 
32'd139573: dataIn1 = 32'd3114
; 
32'd139574: dataIn1 = 32'd3115
; 
32'd139575: dataIn1 = 32'd11028
; 
32'd139576: dataIn1 = 32'd11029
; 
32'd139577: dataIn1 = 32'd302
; 
32'd139578: dataIn1 = 32'd1987
; 
32'd139579: dataIn1 = 32'd2815
; 
32'd139580: dataIn1 = 32'd3112
; 
32'd139581: dataIn1 = 32'd3116
; 
32'd139582: dataIn1 = 32'd4111
; 
32'd139583: dataIn1 = 32'd4120
; 
32'd139584: dataIn1 = 32'd162
; 
32'd139585: dataIn1 = 32'd1987
; 
32'd139586: dataIn1 = 32'd2820
; 
32'd139587: dataIn1 = 32'd3113
; 
32'd139588: dataIn1 = 32'd3117
; 
32'd139589: dataIn1 = 32'd4104
; 
32'd139590: dataIn1 = 32'd4121
; 
32'd139591: dataIn1 = 32'd1747
; 
32'd139592: dataIn1 = 32'd1988
; 
32'd139593: dataIn1 = 32'd2826
; 
32'd139594: dataIn1 = 32'd3118
; 
32'd139595: dataIn1 = 32'd3119
; 
32'd139596: dataIn1 = 32'd3120
; 
32'd139597: dataIn1 = 32'd3121
; 
32'd139598: dataIn1 = 32'd1743
; 
32'd139599: dataIn1 = 32'd1988
; 
32'd139600: dataIn1 = 32'd2816
; 
32'd139601: dataIn1 = 32'd3118
; 
32'd139602: dataIn1 = 32'd3119
; 
32'd139603: dataIn1 = 32'd3120
; 
32'd139604: dataIn1 = 32'd3122
; 
32'd139605: dataIn1 = 32'd1743
; 
32'd139606: dataIn1 = 32'd1747
; 
32'd139607: dataIn1 = 32'd3118
; 
32'd139608: dataIn1 = 32'd3119
; 
32'd139609: dataIn1 = 32'd3120
; 
32'd139610: dataIn1 = 32'd3123
; 
32'd139611: dataIn1 = 32'd3124
; 
32'd139612: dataIn1 = 32'd163
; 
32'd139613: dataIn1 = 32'd1988
; 
32'd139614: dataIn1 = 32'd2826
; 
32'd139615: dataIn1 = 32'd3118
; 
32'd139616: dataIn1 = 32'd3121
; 
32'd139617: dataIn1 = 32'd4115
; 
32'd139618: dataIn1 = 32'd4125
; 
32'd139619: dataIn1 = 32'd302
; 
32'd139620: dataIn1 = 32'd1988
; 
32'd139621: dataIn1 = 32'd2816
; 
32'd139622: dataIn1 = 32'd3119
; 
32'd139623: dataIn1 = 32'd3122
; 
32'd139624: dataIn1 = 32'd4112
; 
32'd139625: dataIn1 = 32'd4116
; 
32'd139626: dataIn1 = 32'd1747
; 
32'd139627: dataIn1 = 32'd2824
; 
32'd139628: dataIn1 = 32'd3120
; 
32'd139629: dataIn1 = 32'd3123
; 
32'd139630: dataIn1 = 32'd3124
; 
32'd139631: dataIn1 = 32'd11033
; 
32'd139632: dataIn1 = 32'd11034
; 
32'd139633: dataIn1 = 32'd1743
; 
32'd139634: dataIn1 = 32'd2814
; 
32'd139635: dataIn1 = 32'd3120
; 
32'd139636: dataIn1 = 32'd3123
; 
32'd139637: dataIn1 = 32'd3124
; 
32'd139638: dataIn1 = 32'd11032
; 
32'd139639: dataIn1 = 32'd11033
; 
32'd139640: dataIn1 = 32'd1748
; 
32'd139641: dataIn1 = 32'd1989
; 
32'd139642: dataIn1 = 32'd2825
; 
32'd139643: dataIn1 = 32'd3125
; 
32'd139644: dataIn1 = 32'd3126
; 
32'd139645: dataIn1 = 32'd3127
; 
32'd139646: dataIn1 = 32'd3128
; 
32'd139647: dataIn1 = 32'd1749
; 
32'd139648: dataIn1 = 32'd1989
; 
32'd139649: dataIn1 = 32'd2831
; 
32'd139650: dataIn1 = 32'd3125
; 
32'd139651: dataIn1 = 32'd3126
; 
32'd139652: dataIn1 = 32'd3127
; 
32'd139653: dataIn1 = 32'd3129
; 
32'd139654: dataIn1 = 32'd1748
; 
32'd139655: dataIn1 = 32'd1749
; 
32'd139656: dataIn1 = 32'd3125
; 
32'd139657: dataIn1 = 32'd3126
; 
32'd139658: dataIn1 = 32'd3127
; 
32'd139659: dataIn1 = 32'd3130
; 
32'd139660: dataIn1 = 32'd3131
; 
32'd139661: dataIn1 = 32'd163
; 
32'd139662: dataIn1 = 32'd1989
; 
32'd139663: dataIn1 = 32'd2825
; 
32'd139664: dataIn1 = 32'd3125
; 
32'd139665: dataIn1 = 32'd3128
; 
32'd139666: dataIn1 = 32'd4126
; 
32'd139667: dataIn1 = 32'd4139
; 
32'd139668: dataIn1 = 32'd309
; 
32'd139669: dataIn1 = 32'd1989
; 
32'd139670: dataIn1 = 32'd2831
; 
32'd139671: dataIn1 = 32'd3126
; 
32'd139672: dataIn1 = 32'd3129
; 
32'd139673: dataIn1 = 32'd4136
; 
32'd139674: dataIn1 = 32'd4140
; 
32'd139675: dataIn1 = 32'd1748
; 
32'd139676: dataIn1 = 32'd2823
; 
32'd139677: dataIn1 = 32'd3127
; 
32'd139678: dataIn1 = 32'd3130
; 
32'd139679: dataIn1 = 32'd3131
; 
32'd139680: dataIn1 = 32'd11036
; 
32'd139681: dataIn1 = 32'd11037
; 
32'd139682: dataIn1 = 32'd1749
; 
32'd139683: dataIn1 = 32'd2829
; 
32'd139684: dataIn1 = 32'd3127
; 
32'd139685: dataIn1 = 32'd3130
; 
32'd139686: dataIn1 = 32'd3131
; 
32'd139687: dataIn1 = 32'd11037
; 
32'd139688: dataIn1 = 32'd11038
; 
32'd139689: dataIn1 = 32'd1750
; 
32'd139690: dataIn1 = 32'd1757
; 
32'd139691: dataIn1 = 32'd3132
; 
32'd139692: dataIn1 = 32'd3133
; 
32'd139693: dataIn1 = 32'd3134
; 
32'd139694: dataIn1 = 32'd3135
; 
32'd139695: dataIn1 = 32'd3136
; 
32'd139696: dataIn1 = 32'd1750
; 
32'd139697: dataIn1 = 32'd1990
; 
32'd139698: dataIn1 = 32'd2830
; 
32'd139699: dataIn1 = 32'd3132
; 
32'd139700: dataIn1 = 32'd3133
; 
32'd139701: dataIn1 = 32'd3134
; 
32'd139702: dataIn1 = 32'd3137
; 
32'd139703: dataIn1 = 32'd1757
; 
32'd139704: dataIn1 = 32'd1990
; 
32'd139705: dataIn1 = 32'd2851
; 
32'd139706: dataIn1 = 32'd3132
; 
32'd139707: dataIn1 = 32'd3133
; 
32'd139708: dataIn1 = 32'd3134
; 
32'd139709: dataIn1 = 32'd3138
; 
32'd139710: dataIn1 = 32'd1750
; 
32'd139711: dataIn1 = 32'd2827
; 
32'd139712: dataIn1 = 32'd3132
; 
32'd139713: dataIn1 = 32'd3135
; 
32'd139714: dataIn1 = 32'd3136
; 
32'd139715: dataIn1 = 32'd11040
; 
32'd139716: dataIn1 = 32'd11041
; 
32'd139717: dataIn1 = 32'd1757
; 
32'd139718: dataIn1 = 32'd2849
; 
32'd139719: dataIn1 = 32'd3132
; 
32'd139720: dataIn1 = 32'd3135
; 
32'd139721: dataIn1 = 32'd3136
; 
32'd139722: dataIn1 = 32'd11041
; 
32'd139723: dataIn1 = 32'd11042
; 
32'd139724: dataIn1 = 32'd309
; 
32'd139725: dataIn1 = 32'd1990
; 
32'd139726: dataIn1 = 32'd2830
; 
32'd139727: dataIn1 = 32'd3133
; 
32'd139728: dataIn1 = 32'd3137
; 
32'd139729: dataIn1 = 32'd4135
; 
32'd139730: dataIn1 = 32'd4143
; 
32'd139731: dataIn1 = 32'd165
; 
32'd139732: dataIn1 = 32'd1990
; 
32'd139733: dataIn1 = 32'd2851
; 
32'd139734: dataIn1 = 32'd3134
; 
32'd139735: dataIn1 = 32'd3138
; 
32'd139736: dataIn1 = 32'd4144
; 
32'd139737: dataIn1 = 32'd4152
; 
32'd139738: dataIn1 = 32'd1752
; 
32'd139739: dataIn1 = 32'd1991
; 
32'd139740: dataIn1 = 32'd2835
; 
32'd139741: dataIn1 = 32'd3139
; 
32'd139742: dataIn1 = 32'd3140
; 
32'd139743: dataIn1 = 32'd3141
; 
32'd139744: dataIn1 = 32'd3142
; 
32'd139745: dataIn1 = 32'd1752
; 
32'd139746: dataIn1 = 32'd1761
; 
32'd139747: dataIn1 = 32'd3139
; 
32'd139748: dataIn1 = 32'd3140
; 
32'd139749: dataIn1 = 32'd3141
; 
32'd139750: dataIn1 = 32'd3143
; 
32'd139751: dataIn1 = 32'd3144
; 
32'd139752: dataIn1 = 32'd1761
; 
32'd139753: dataIn1 = 32'd1991
; 
32'd139754: dataIn1 = 32'd2861
; 
32'd139755: dataIn1 = 32'd3139
; 
32'd139756: dataIn1 = 32'd3140
; 
32'd139757: dataIn1 = 32'd3141
; 
32'd139758: dataIn1 = 32'd3145
; 
32'd139759: dataIn1 = 32'd311
; 
32'd139760: dataIn1 = 32'd1991
; 
32'd139761: dataIn1 = 32'd2835
; 
32'd139762: dataIn1 = 32'd3139
; 
32'd139763: dataIn1 = 32'd3142
; 
32'd139764: dataIn1 = 32'd4181
; 
32'd139765: dataIn1 = 32'd4190
; 
32'd139766: dataIn1 = 32'd1752
; 
32'd139767: dataIn1 = 32'd2833
; 
32'd139768: dataIn1 = 32'd3140
; 
32'd139769: dataIn1 = 32'd3143
; 
32'd139770: dataIn1 = 32'd3144
; 
32'd139771: dataIn1 = 32'd11056
; 
32'd139772: dataIn1 = 32'd11057
; 
32'd139773: dataIn1 = 32'd1761
; 
32'd139774: dataIn1 = 32'd2858
; 
32'd139775: dataIn1 = 32'd3140
; 
32'd139776: dataIn1 = 32'd3143
; 
32'd139777: dataIn1 = 32'd3144
; 
32'd139778: dataIn1 = 32'd11057
; 
32'd139779: dataIn1 = 32'd11058
; 
32'd139780: dataIn1 = 32'd168
; 
32'd139781: dataIn1 = 32'd1991
; 
32'd139782: dataIn1 = 32'd2861
; 
32'd139783: dataIn1 = 32'd3141
; 
32'd139784: dataIn1 = 32'd3145
; 
32'd139785: dataIn1 = 32'd4192
; 
32'd139786: dataIn1 = 32'd4201
; 
32'd139787: dataIn1 = 32'd1751
; 
32'd139788: dataIn1 = 32'd1992
; 
32'd139789: dataIn1 = 32'd2836
; 
32'd139790: dataIn1 = 32'd3146
; 
32'd139791: dataIn1 = 32'd3147
; 
32'd139792: dataIn1 = 32'd3148
; 
32'd139793: dataIn1 = 32'd3149
; 
32'd139794: dataIn1 = 32'd1755
; 
32'd139795: dataIn1 = 32'd1992
; 
32'd139796: dataIn1 = 32'd2846
; 
32'd139797: dataIn1 = 32'd3146
; 
32'd139798: dataIn1 = 32'd3147
; 
32'd139799: dataIn1 = 32'd3148
; 
32'd139800: dataIn1 = 32'd3150
; 
32'd139801: dataIn1 = 32'd1751
; 
32'd139802: dataIn1 = 32'd1755
; 
32'd139803: dataIn1 = 32'd3146
; 
32'd139804: dataIn1 = 32'd3147
; 
32'd139805: dataIn1 = 32'd3148
; 
32'd139806: dataIn1 = 32'd3151
; 
32'd139807: dataIn1 = 32'd3152
; 
32'd139808: dataIn1 = 32'd311
; 
32'd139809: dataIn1 = 32'd1992
; 
32'd139810: dataIn1 = 32'd2836
; 
32'd139811: dataIn1 = 32'd3146
; 
32'd139812: dataIn1 = 32'd3149
; 
32'd139813: dataIn1 = 32'd4182
; 
32'd139814: dataIn1 = 32'd4187
; 
32'd139815: dataIn1 = 32'd167
; 
32'd139816: dataIn1 = 32'd1992
; 
32'd139817: dataIn1 = 32'd2846
; 
32'd139818: dataIn1 = 32'd3147
; 
32'd139819: dataIn1 = 32'd3150
; 
32'd139820: dataIn1 = 32'd4175
; 
32'd139821: dataIn1 = 32'd4188
; 
32'd139822: dataIn1 = 32'd1751
; 
32'd139823: dataIn1 = 32'd2834
; 
32'd139824: dataIn1 = 32'd3148
; 
32'd139825: dataIn1 = 32'd3151
; 
32'd139826: dataIn1 = 32'd3152
; 
32'd139827: dataIn1 = 32'd11053
; 
32'd139828: dataIn1 = 32'd11054
; 
32'd139829: dataIn1 = 32'd1755
; 
32'd139830: dataIn1 = 32'd2844
; 
32'd139831: dataIn1 = 32'd3148
; 
32'd139832: dataIn1 = 32'd3151
; 
32'd139833: dataIn1 = 32'd3152
; 
32'd139834: dataIn1 = 32'd11052
; 
32'd139835: dataIn1 = 32'd11053
; 
32'd139836: dataIn1 = 32'd1754
; 
32'd139837: dataIn1 = 32'd1756
; 
32'd139838: dataIn1 = 32'd3153
; 
32'd139839: dataIn1 = 32'd3154
; 
32'd139840: dataIn1 = 32'd3155
; 
32'd139841: dataIn1 = 32'd3156
; 
32'd139842: dataIn1 = 32'd3157
; 
32'd139843: dataIn1 = 32'd1756
; 
32'd139844: dataIn1 = 32'd1993
; 
32'd139845: dataIn1 = 32'd2845
; 
32'd139846: dataIn1 = 32'd3153
; 
32'd139847: dataIn1 = 32'd3154
; 
32'd139848: dataIn1 = 32'd3155
; 
32'd139849: dataIn1 = 32'd3158
; 
32'd139850: dataIn1 = 32'd1754
; 
32'd139851: dataIn1 = 32'd1993
; 
32'd139852: dataIn1 = 32'd2840
; 
32'd139853: dataIn1 = 32'd3153
; 
32'd139854: dataIn1 = 32'd3154
; 
32'd139855: dataIn1 = 32'd3155
; 
32'd139856: dataIn1 = 32'd3159
; 
32'd139857: dataIn1 = 32'd1756
; 
32'd139858: dataIn1 = 32'd2842
; 
32'd139859: dataIn1 = 32'd3153
; 
32'd139860: dataIn1 = 32'd3156
; 
32'd139861: dataIn1 = 32'd3157
; 
32'd139862: dataIn1 = 32'd11049
; 
32'd139863: dataIn1 = 32'd11050
; 
32'd139864: dataIn1 = 32'd1754
; 
32'd139865: dataIn1 = 32'd2837
; 
32'd139866: dataIn1 = 32'd3153
; 
32'd139867: dataIn1 = 32'd3156
; 
32'd139868: dataIn1 = 32'd3157
; 
32'd139869: dataIn1 = 32'd11048
; 
32'd139870: dataIn1 = 32'd11049
; 
32'd139871: dataIn1 = 32'd167
; 
32'd139872: dataIn1 = 32'd1993
; 
32'd139873: dataIn1 = 32'd2845
; 
32'd139874: dataIn1 = 32'd3154
; 
32'd139875: dataIn1 = 32'd3158
; 
32'd139876: dataIn1 = 32'd4167
; 
32'd139877: dataIn1 = 32'd4174
; 
32'd139878: dataIn1 = 32'd317
; 
32'd139879: dataIn1 = 32'd1993
; 
32'd139880: dataIn1 = 32'd2840
; 
32'd139881: dataIn1 = 32'd3155
; 
32'd139882: dataIn1 = 32'd3159
; 
32'd139883: dataIn1 = 32'd4161
; 
32'd139884: dataIn1 = 32'd4168
; 
32'd139885: dataIn1 = 32'd1758
; 
32'd139886: dataIn1 = 32'd1994
; 
32'd139887: dataIn1 = 32'd2850
; 
32'd139888: dataIn1 = 32'd3160
; 
32'd139889: dataIn1 = 32'd3161
; 
32'd139890: dataIn1 = 32'd3162
; 
32'd139891: dataIn1 = 32'd3163
; 
32'd139892: dataIn1 = 32'd1753
; 
32'd139893: dataIn1 = 32'd1758
; 
32'd139894: dataIn1 = 32'd3160
; 
32'd139895: dataIn1 = 32'd3161
; 
32'd139896: dataIn1 = 32'd3162
; 
32'd139897: dataIn1 = 32'd3164
; 
32'd139898: dataIn1 = 32'd3165
; 
32'd139899: dataIn1 = 32'd1753
; 
32'd139900: dataIn1 = 32'd1994
; 
32'd139901: dataIn1 = 32'd2841
; 
32'd139902: dataIn1 = 32'd3160
; 
32'd139903: dataIn1 = 32'd3161
; 
32'd139904: dataIn1 = 32'd3162
; 
32'd139905: dataIn1 = 32'd3166
; 
32'd139906: dataIn1 = 32'd165
; 
32'd139907: dataIn1 = 32'd1994
; 
32'd139908: dataIn1 = 32'd2850
; 
32'd139909: dataIn1 = 32'd3160
; 
32'd139910: dataIn1 = 32'd3163
; 
32'd139911: dataIn1 = 32'd4153
; 
32'd139912: dataIn1 = 32'd4163
; 
32'd139913: dataIn1 = 32'd1758
; 
32'd139914: dataIn1 = 32'd2848
; 
32'd139915: dataIn1 = 32'd3161
; 
32'd139916: dataIn1 = 32'd3164
; 
32'd139917: dataIn1 = 32'd3165
; 
32'd139918: dataIn1 = 32'd11044
; 
32'd139919: dataIn1 = 32'd11045
; 
32'd139920: dataIn1 = 32'd1753
; 
32'd139921: dataIn1 = 32'd2838
; 
32'd139922: dataIn1 = 32'd3161
; 
32'd139923: dataIn1 = 32'd3164
; 
32'd139924: dataIn1 = 32'd3165
; 
32'd139925: dataIn1 = 32'd11045
; 
32'd139926: dataIn1 = 32'd11046
; 
32'd139927: dataIn1 = 32'd317
; 
32'd139928: dataIn1 = 32'd1994
; 
32'd139929: dataIn1 = 32'd2841
; 
32'd139930: dataIn1 = 32'd3162
; 
32'd139931: dataIn1 = 32'd3166
; 
32'd139932: dataIn1 = 32'd4162
; 
32'd139933: dataIn1 = 32'd4165
; 
32'd139934: dataIn1 = 32'd1760
; 
32'd139935: dataIn1 = 32'd1762
; 
32'd139936: dataIn1 = 32'd3167
; 
32'd139937: dataIn1 = 32'd3168
; 
32'd139938: dataIn1 = 32'd3169
; 
32'd139939: dataIn1 = 32'd3170
; 
32'd139940: dataIn1 = 32'd3171
; 
32'd139941: dataIn1 = 32'd1760
; 
32'd139942: dataIn1 = 32'd1995
; 
32'd139943: dataIn1 = 32'd2855
; 
32'd139944: dataIn1 = 32'd3167
; 
32'd139945: dataIn1 = 32'd3168
; 
32'd139946: dataIn1 = 32'd3169
; 
32'd139947: dataIn1 = 32'd3172
; 
32'd139948: dataIn1 = 32'd1762
; 
32'd139949: dataIn1 = 32'd1995
; 
32'd139950: dataIn1 = 32'd2860
; 
32'd139951: dataIn1 = 32'd3167
; 
32'd139952: dataIn1 = 32'd3168
; 
32'd139953: dataIn1 = 32'd3169
; 
32'd139954: dataIn1 = 32'd3173
; 
32'd139955: dataIn1 = 32'd1760
; 
32'd139956: dataIn1 = 32'd2852
; 
32'd139957: dataIn1 = 32'd3167
; 
32'd139958: dataIn1 = 32'd3170
; 
32'd139959: dataIn1 = 32'd3171
; 
32'd139960: dataIn1 = 32'd11061
; 
32'd139961: dataIn1 = 32'd11062
; 
32'd139962: dataIn1 = 32'd1762
; 
32'd139963: dataIn1 = 32'd2857
; 
32'd139964: dataIn1 = 32'd3167
; 
32'd139965: dataIn1 = 32'd3170
; 
32'd139966: dataIn1 = 32'd3171
; 
32'd139967: dataIn1 = 32'd11060
; 
32'd139968: dataIn1 = 32'd11061
; 
32'd139969: dataIn1 = 32'd318
; 
32'd139970: dataIn1 = 32'd1995
; 
32'd139971: dataIn1 = 32'd2855
; 
32'd139972: dataIn1 = 32'd3168
; 
32'd139973: dataIn1 = 32'd3172
; 
32'd139974: dataIn1 = 32'd4207
; 
32'd139975: dataIn1 = 32'd4216
; 
32'd139976: dataIn1 = 32'd168
; 
32'd139977: dataIn1 = 32'd1995
; 
32'd139978: dataIn1 = 32'd2860
; 
32'd139979: dataIn1 = 32'd3169
; 
32'd139980: dataIn1 = 32'd3173
; 
32'd139981: dataIn1 = 32'd4200
; 
32'd139982: dataIn1 = 32'd4217
; 
32'd139983: dataIn1 = 32'd1763
; 
32'd139984: dataIn1 = 32'd1996
; 
32'd139985: dataIn1 = 32'd2866
; 
32'd139986: dataIn1 = 32'd3174
; 
32'd139987: dataIn1 = 32'd3175
; 
32'd139988: dataIn1 = 32'd3176
; 
32'd139989: dataIn1 = 32'd3177
; 
32'd139990: dataIn1 = 32'd1759
; 
32'd139991: dataIn1 = 32'd1996
; 
32'd139992: dataIn1 = 32'd2856
; 
32'd139993: dataIn1 = 32'd3174
; 
32'd139994: dataIn1 = 32'd3175
; 
32'd139995: dataIn1 = 32'd3176
; 
32'd139996: dataIn1 = 32'd3178
; 
32'd139997: dataIn1 = 32'd1759
; 
32'd139998: dataIn1 = 32'd1763
; 
32'd139999: dataIn1 = 32'd3174
; 
32'd140000: dataIn1 = 32'd3175
; 
32'd140001: dataIn1 = 32'd3176
; 
32'd140002: dataIn1 = 32'd3179
; 
32'd140003: dataIn1 = 32'd3180
; 
32'd140004: dataIn1 = 32'd169
; 
32'd140005: dataIn1 = 32'd1996
; 
32'd140006: dataIn1 = 32'd2866
; 
32'd140007: dataIn1 = 32'd3174
; 
32'd140008: dataIn1 = 32'd3177
; 
32'd140009: dataIn1 = 32'd4211
; 
32'd140010: dataIn1 = 32'd4221
; 
32'd140011: dataIn1 = 32'd318
; 
32'd140012: dataIn1 = 32'd1996
; 
32'd140013: dataIn1 = 32'd2856
; 
32'd140014: dataIn1 = 32'd3175
; 
32'd140015: dataIn1 = 32'd3178
; 
32'd140016: dataIn1 = 32'd4208
; 
32'd140017: dataIn1 = 32'd4212
; 
32'd140018: dataIn1 = 32'd1763
; 
32'd140019: dataIn1 = 32'd2864
; 
32'd140020: dataIn1 = 32'd3176
; 
32'd140021: dataIn1 = 32'd3179
; 
32'd140022: dataIn1 = 32'd3180
; 
32'd140023: dataIn1 = 32'd11065
; 
32'd140024: dataIn1 = 32'd11066
; 
32'd140025: dataIn1 = 32'd1759
; 
32'd140026: dataIn1 = 32'd2854
; 
32'd140027: dataIn1 = 32'd3176
; 
32'd140028: dataIn1 = 32'd3179
; 
32'd140029: dataIn1 = 32'd3180
; 
32'd140030: dataIn1 = 32'd11064
; 
32'd140031: dataIn1 = 32'd11065
; 
32'd140032: dataIn1 = 32'd1764
; 
32'd140033: dataIn1 = 32'd1997
; 
32'd140034: dataIn1 = 32'd2865
; 
32'd140035: dataIn1 = 32'd3181
; 
32'd140036: dataIn1 = 32'd3182
; 
32'd140037: dataIn1 = 32'd3183
; 
32'd140038: dataIn1 = 32'd3184
; 
32'd140039: dataIn1 = 32'd1765
; 
32'd140040: dataIn1 = 32'd1997
; 
32'd140041: dataIn1 = 32'd2871
; 
32'd140042: dataIn1 = 32'd3181
; 
32'd140043: dataIn1 = 32'd3182
; 
32'd140044: dataIn1 = 32'd3183
; 
32'd140045: dataIn1 = 32'd3185
; 
32'd140046: dataIn1 = 32'd1764
; 
32'd140047: dataIn1 = 32'd1765
; 
32'd140048: dataIn1 = 32'd3181
; 
32'd140049: dataIn1 = 32'd3182
; 
32'd140050: dataIn1 = 32'd3183
; 
32'd140051: dataIn1 = 32'd3186
; 
32'd140052: dataIn1 = 32'd3187
; 
32'd140053: dataIn1 = 32'd169
; 
32'd140054: dataIn1 = 32'd1997
; 
32'd140055: dataIn1 = 32'd2865
; 
32'd140056: dataIn1 = 32'd3181
; 
32'd140057: dataIn1 = 32'd3184
; 
32'd140058: dataIn1 = 32'd4222
; 
32'd140059: dataIn1 = 32'd4235
; 
32'd140060: dataIn1 = 32'd325
; 
32'd140061: dataIn1 = 32'd1997
; 
32'd140062: dataIn1 = 32'd2871
; 
32'd140063: dataIn1 = 32'd3182
; 
32'd140064: dataIn1 = 32'd3185
; 
32'd140065: dataIn1 = 32'd4232
; 
32'd140066: dataIn1 = 32'd4236
; 
32'd140067: dataIn1 = 32'd1764
; 
32'd140068: dataIn1 = 32'd2863
; 
32'd140069: dataIn1 = 32'd3183
; 
32'd140070: dataIn1 = 32'd3186
; 
32'd140071: dataIn1 = 32'd3187
; 
32'd140072: dataIn1 = 32'd11068
; 
32'd140073: dataIn1 = 32'd11069
; 
32'd140074: dataIn1 = 32'd1765
; 
32'd140075: dataIn1 = 32'd2869
; 
32'd140076: dataIn1 = 32'd3183
; 
32'd140077: dataIn1 = 32'd3186
; 
32'd140078: dataIn1 = 32'd3187
; 
32'd140079: dataIn1 = 32'd11069
; 
32'd140080: dataIn1 = 32'd11070
; 
32'd140081: dataIn1 = 32'd1766
; 
32'd140082: dataIn1 = 32'd1773
; 
32'd140083: dataIn1 = 32'd3188
; 
32'd140084: dataIn1 = 32'd3189
; 
32'd140085: dataIn1 = 32'd3190
; 
32'd140086: dataIn1 = 32'd3191
; 
32'd140087: dataIn1 = 32'd3192
; 
32'd140088: dataIn1 = 32'd1766
; 
32'd140089: dataIn1 = 32'd1998
; 
32'd140090: dataIn1 = 32'd2870
; 
32'd140091: dataIn1 = 32'd3188
; 
32'd140092: dataIn1 = 32'd3189
; 
32'd140093: dataIn1 = 32'd3190
; 
32'd140094: dataIn1 = 32'd3193
; 
32'd140095: dataIn1 = 32'd1773
; 
32'd140096: dataIn1 = 32'd1998
; 
32'd140097: dataIn1 = 32'd2891
; 
32'd140098: dataIn1 = 32'd3188
; 
32'd140099: dataIn1 = 32'd3189
; 
32'd140100: dataIn1 = 32'd3190
; 
32'd140101: dataIn1 = 32'd3194
; 
32'd140102: dataIn1 = 32'd1766
; 
32'd140103: dataIn1 = 32'd2867
; 
32'd140104: dataIn1 = 32'd3188
; 
32'd140105: dataIn1 = 32'd3191
; 
32'd140106: dataIn1 = 32'd3192
; 
32'd140107: dataIn1 = 32'd11072
; 
32'd140108: dataIn1 = 32'd11073
; 
32'd140109: dataIn1 = 32'd1773
; 
32'd140110: dataIn1 = 32'd2889
; 
32'd140111: dataIn1 = 32'd3188
; 
32'd140112: dataIn1 = 32'd3191
; 
32'd140113: dataIn1 = 32'd3192
; 
32'd140114: dataIn1 = 32'd11073
; 
32'd140115: dataIn1 = 32'd11074
; 
32'd140116: dataIn1 = 32'd325
; 
32'd140117: dataIn1 = 32'd1998
; 
32'd140118: dataIn1 = 32'd2870
; 
32'd140119: dataIn1 = 32'd3189
; 
32'd140120: dataIn1 = 32'd3193
; 
32'd140121: dataIn1 = 32'd4231
; 
32'd140122: dataIn1 = 32'd4239
; 
32'd140123: dataIn1 = 32'd171
; 
32'd140124: dataIn1 = 32'd1998
; 
32'd140125: dataIn1 = 32'd2891
; 
32'd140126: dataIn1 = 32'd3190
; 
32'd140127: dataIn1 = 32'd3194
; 
32'd140128: dataIn1 = 32'd4240
; 
32'd140129: dataIn1 = 32'd4248
; 
32'd140130: dataIn1 = 32'd1768
; 
32'd140131: dataIn1 = 32'd1999
; 
32'd140132: dataIn1 = 32'd2875
; 
32'd140133: dataIn1 = 32'd3195
; 
32'd140134: dataIn1 = 32'd3196
; 
32'd140135: dataIn1 = 32'd3197
; 
32'd140136: dataIn1 = 32'd3198
; 
32'd140137: dataIn1 = 32'd1768
; 
32'd140138: dataIn1 = 32'd1777
; 
32'd140139: dataIn1 = 32'd3195
; 
32'd140140: dataIn1 = 32'd3196
; 
32'd140141: dataIn1 = 32'd3197
; 
32'd140142: dataIn1 = 32'd3199
; 
32'd140143: dataIn1 = 32'd3200
; 
32'd140144: dataIn1 = 32'd1777
; 
32'd140145: dataIn1 = 32'd1999
; 
32'd140146: dataIn1 = 32'd2901
; 
32'd140147: dataIn1 = 32'd3195
; 
32'd140148: dataIn1 = 32'd3196
; 
32'd140149: dataIn1 = 32'd3197
; 
32'd140150: dataIn1 = 32'd3201
; 
32'd140151: dataIn1 = 32'd327
; 
32'd140152: dataIn1 = 32'd1999
; 
32'd140153: dataIn1 = 32'd2875
; 
32'd140154: dataIn1 = 32'd3195
; 
32'd140155: dataIn1 = 32'd3198
; 
32'd140156: dataIn1 = 32'd4277
; 
32'd140157: dataIn1 = 32'd4286
; 
32'd140158: dataIn1 = 32'd1768
; 
32'd140159: dataIn1 = 32'd2873
; 
32'd140160: dataIn1 = 32'd3196
; 
32'd140161: dataIn1 = 32'd3199
; 
32'd140162: dataIn1 = 32'd3200
; 
32'd140163: dataIn1 = 32'd11088
; 
32'd140164: dataIn1 = 32'd11089
; 
32'd140165: dataIn1 = 32'd1777
; 
32'd140166: dataIn1 = 32'd2898
; 
32'd140167: dataIn1 = 32'd3196
; 
32'd140168: dataIn1 = 32'd3199
; 
32'd140169: dataIn1 = 32'd3200
; 
32'd140170: dataIn1 = 32'd11089
; 
32'd140171: dataIn1 = 32'd11090
; 
32'd140172: dataIn1 = 32'd174
; 
32'd140173: dataIn1 = 32'd1999
; 
32'd140174: dataIn1 = 32'd2901
; 
32'd140175: dataIn1 = 32'd3197
; 
32'd140176: dataIn1 = 32'd3201
; 
32'd140177: dataIn1 = 32'd4288
; 
32'd140178: dataIn1 = 32'd4297
; 
32'd140179: dataIn1 = 32'd1767
; 
32'd140180: dataIn1 = 32'd2000
; 
32'd140181: dataIn1 = 32'd2876
; 
32'd140182: dataIn1 = 32'd3202
; 
32'd140183: dataIn1 = 32'd3203
; 
32'd140184: dataIn1 = 32'd3204
; 
32'd140185: dataIn1 = 32'd3205
; 
32'd140186: dataIn1 = 32'd1771
; 
32'd140187: dataIn1 = 32'd2000
; 
32'd140188: dataIn1 = 32'd2886
; 
32'd140189: dataIn1 = 32'd3202
; 
32'd140190: dataIn1 = 32'd3203
; 
32'd140191: dataIn1 = 32'd3204
; 
32'd140192: dataIn1 = 32'd3206
; 
32'd140193: dataIn1 = 32'd1767
; 
32'd140194: dataIn1 = 32'd1771
; 
32'd140195: dataIn1 = 32'd3202
; 
32'd140196: dataIn1 = 32'd3203
; 
32'd140197: dataIn1 = 32'd3204
; 
32'd140198: dataIn1 = 32'd3207
; 
32'd140199: dataIn1 = 32'd3208
; 
32'd140200: dataIn1 = 32'd327
; 
32'd140201: dataIn1 = 32'd2000
; 
32'd140202: dataIn1 = 32'd2876
; 
32'd140203: dataIn1 = 32'd3202
; 
32'd140204: dataIn1 = 32'd3205
; 
32'd140205: dataIn1 = 32'd4278
; 
32'd140206: dataIn1 = 32'd4283
; 
32'd140207: dataIn1 = 32'd173
; 
32'd140208: dataIn1 = 32'd2000
; 
32'd140209: dataIn1 = 32'd2886
; 
32'd140210: dataIn1 = 32'd3203
; 
32'd140211: dataIn1 = 32'd3206
; 
32'd140212: dataIn1 = 32'd4271
; 
32'd140213: dataIn1 = 32'd4284
; 
32'd140214: dataIn1 = 32'd1767
; 
32'd140215: dataIn1 = 32'd2874
; 
32'd140216: dataIn1 = 32'd3204
; 
32'd140217: dataIn1 = 32'd3207
; 
32'd140218: dataIn1 = 32'd3208
; 
32'd140219: dataIn1 = 32'd11085
; 
32'd140220: dataIn1 = 32'd11086
; 
32'd140221: dataIn1 = 32'd1771
; 
32'd140222: dataIn1 = 32'd2884
; 
32'd140223: dataIn1 = 32'd3204
; 
32'd140224: dataIn1 = 32'd3207
; 
32'd140225: dataIn1 = 32'd3208
; 
32'd140226: dataIn1 = 32'd11084
; 
32'd140227: dataIn1 = 32'd11085
; 
32'd140228: dataIn1 = 32'd1770
; 
32'd140229: dataIn1 = 32'd1772
; 
32'd140230: dataIn1 = 32'd3209
; 
32'd140231: dataIn1 = 32'd3210
; 
32'd140232: dataIn1 = 32'd3211
; 
32'd140233: dataIn1 = 32'd3212
; 
32'd140234: dataIn1 = 32'd3213
; 
32'd140235: dataIn1 = 32'd1772
; 
32'd140236: dataIn1 = 32'd2001
; 
32'd140237: dataIn1 = 32'd2885
; 
32'd140238: dataIn1 = 32'd3209
; 
32'd140239: dataIn1 = 32'd3210
; 
32'd140240: dataIn1 = 32'd3211
; 
32'd140241: dataIn1 = 32'd3214
; 
32'd140242: dataIn1 = 32'd1770
; 
32'd140243: dataIn1 = 32'd2001
; 
32'd140244: dataIn1 = 32'd2880
; 
32'd140245: dataIn1 = 32'd3209
; 
32'd140246: dataIn1 = 32'd3210
; 
32'd140247: dataIn1 = 32'd3211
; 
32'd140248: dataIn1 = 32'd3215
; 
32'd140249: dataIn1 = 32'd1772
; 
32'd140250: dataIn1 = 32'd2882
; 
32'd140251: dataIn1 = 32'd3209
; 
32'd140252: dataIn1 = 32'd3212
; 
32'd140253: dataIn1 = 32'd3213
; 
32'd140254: dataIn1 = 32'd11081
; 
32'd140255: dataIn1 = 32'd11082
; 
32'd140256: dataIn1 = 32'd1770
; 
32'd140257: dataIn1 = 32'd2877
; 
32'd140258: dataIn1 = 32'd3209
; 
32'd140259: dataIn1 = 32'd3212
; 
32'd140260: dataIn1 = 32'd3213
; 
32'd140261: dataIn1 = 32'd11080
; 
32'd140262: dataIn1 = 32'd11081
; 
32'd140263: dataIn1 = 32'd173
; 
32'd140264: dataIn1 = 32'd2001
; 
32'd140265: dataIn1 = 32'd2885
; 
32'd140266: dataIn1 = 32'd3210
; 
32'd140267: dataIn1 = 32'd3214
; 
32'd140268: dataIn1 = 32'd4263
; 
32'd140269: dataIn1 = 32'd4270
; 
32'd140270: dataIn1 = 32'd333
; 
32'd140271: dataIn1 = 32'd2001
; 
32'd140272: dataIn1 = 32'd2880
; 
32'd140273: dataIn1 = 32'd3211
; 
32'd140274: dataIn1 = 32'd3215
; 
32'd140275: dataIn1 = 32'd4257
; 
32'd140276: dataIn1 = 32'd4264
; 
32'd140277: dataIn1 = 32'd1774
; 
32'd140278: dataIn1 = 32'd2002
; 
32'd140279: dataIn1 = 32'd2890
; 
32'd140280: dataIn1 = 32'd3216
; 
32'd140281: dataIn1 = 32'd3217
; 
32'd140282: dataIn1 = 32'd3218
; 
32'd140283: dataIn1 = 32'd3219
; 
32'd140284: dataIn1 = 32'd1769
; 
32'd140285: dataIn1 = 32'd1774
; 
32'd140286: dataIn1 = 32'd3216
; 
32'd140287: dataIn1 = 32'd3217
; 
32'd140288: dataIn1 = 32'd3218
; 
32'd140289: dataIn1 = 32'd3220
; 
32'd140290: dataIn1 = 32'd3221
; 
32'd140291: dataIn1 = 32'd1769
; 
32'd140292: dataIn1 = 32'd2002
; 
32'd140293: dataIn1 = 32'd2881
; 
32'd140294: dataIn1 = 32'd3216
; 
32'd140295: dataIn1 = 32'd3217
; 
32'd140296: dataIn1 = 32'd3218
; 
32'd140297: dataIn1 = 32'd3222
; 
32'd140298: dataIn1 = 32'd171
; 
32'd140299: dataIn1 = 32'd2002
; 
32'd140300: dataIn1 = 32'd2890
; 
32'd140301: dataIn1 = 32'd3216
; 
32'd140302: dataIn1 = 32'd3219
; 
32'd140303: dataIn1 = 32'd4249
; 
32'd140304: dataIn1 = 32'd4259
; 
32'd140305: dataIn1 = 32'd1774
; 
32'd140306: dataIn1 = 32'd2888
; 
32'd140307: dataIn1 = 32'd3217
; 
32'd140308: dataIn1 = 32'd3220
; 
32'd140309: dataIn1 = 32'd3221
; 
32'd140310: dataIn1 = 32'd11076
; 
32'd140311: dataIn1 = 32'd11077
; 
32'd140312: dataIn1 = 32'd1769
; 
32'd140313: dataIn1 = 32'd2878
; 
32'd140314: dataIn1 = 32'd3217
; 
32'd140315: dataIn1 = 32'd3220
; 
32'd140316: dataIn1 = 32'd3221
; 
32'd140317: dataIn1 = 32'd11077
; 
32'd140318: dataIn1 = 32'd11078
; 
32'd140319: dataIn1 = 32'd333
; 
32'd140320: dataIn1 = 32'd2002
; 
32'd140321: dataIn1 = 32'd2881
; 
32'd140322: dataIn1 = 32'd3218
; 
32'd140323: dataIn1 = 32'd3222
; 
32'd140324: dataIn1 = 32'd4258
; 
32'd140325: dataIn1 = 32'd4261
; 
32'd140326: dataIn1 = 32'd1776
; 
32'd140327: dataIn1 = 32'd1778
; 
32'd140328: dataIn1 = 32'd3223
; 
32'd140329: dataIn1 = 32'd3224
; 
32'd140330: dataIn1 = 32'd3225
; 
32'd140331: dataIn1 = 32'd3226
; 
32'd140332: dataIn1 = 32'd3227
; 
32'd140333: dataIn1 = 32'd1776
; 
32'd140334: dataIn1 = 32'd2003
; 
32'd140335: dataIn1 = 32'd2895
; 
32'd140336: dataIn1 = 32'd3223
; 
32'd140337: dataIn1 = 32'd3224
; 
32'd140338: dataIn1 = 32'd3225
; 
32'd140339: dataIn1 = 32'd3228
; 
32'd140340: dataIn1 = 32'd1778
; 
32'd140341: dataIn1 = 32'd2003
; 
32'd140342: dataIn1 = 32'd2900
; 
32'd140343: dataIn1 = 32'd3223
; 
32'd140344: dataIn1 = 32'd3224
; 
32'd140345: dataIn1 = 32'd3225
; 
32'd140346: dataIn1 = 32'd3229
; 
32'd140347: dataIn1 = 32'd1776
; 
32'd140348: dataIn1 = 32'd2892
; 
32'd140349: dataIn1 = 32'd3223
; 
32'd140350: dataIn1 = 32'd3226
; 
32'd140351: dataIn1 = 32'd3227
; 
32'd140352: dataIn1 = 32'd11093
; 
32'd140353: dataIn1 = 32'd11094
; 
32'd140354: dataIn1 = 32'd1778
; 
32'd140355: dataIn1 = 32'd2897
; 
32'd140356: dataIn1 = 32'd3223
; 
32'd140357: dataIn1 = 32'd3226
; 
32'd140358: dataIn1 = 32'd3227
; 
32'd140359: dataIn1 = 32'd11092
; 
32'd140360: dataIn1 = 32'd11093
; 
32'd140361: dataIn1 = 32'd334
; 
32'd140362: dataIn1 = 32'd2003
; 
32'd140363: dataIn1 = 32'd2895
; 
32'd140364: dataIn1 = 32'd3224
; 
32'd140365: dataIn1 = 32'd3228
; 
32'd140366: dataIn1 = 32'd4303
; 
32'd140367: dataIn1 = 32'd4312
; 
32'd140368: dataIn1 = 32'd174
; 
32'd140369: dataIn1 = 32'd2003
; 
32'd140370: dataIn1 = 32'd2900
; 
32'd140371: dataIn1 = 32'd3225
; 
32'd140372: dataIn1 = 32'd3229
; 
32'd140373: dataIn1 = 32'd4296
; 
32'd140374: dataIn1 = 32'd4313
; 
32'd140375: dataIn1 = 32'd1779
; 
32'd140376: dataIn1 = 32'd2004
; 
32'd140377: dataIn1 = 32'd2906
; 
32'd140378: dataIn1 = 32'd3230
; 
32'd140379: dataIn1 = 32'd3231
; 
32'd140380: dataIn1 = 32'd3232
; 
32'd140381: dataIn1 = 32'd3233
; 
32'd140382: dataIn1 = 32'd1775
; 
32'd140383: dataIn1 = 32'd2004
; 
32'd140384: dataIn1 = 32'd2896
; 
32'd140385: dataIn1 = 32'd3230
; 
32'd140386: dataIn1 = 32'd3231
; 
32'd140387: dataIn1 = 32'd3232
; 
32'd140388: dataIn1 = 32'd3234
; 
32'd140389: dataIn1 = 32'd1775
; 
32'd140390: dataIn1 = 32'd1779
; 
32'd140391: dataIn1 = 32'd3230
; 
32'd140392: dataIn1 = 32'd3231
; 
32'd140393: dataIn1 = 32'd3232
; 
32'd140394: dataIn1 = 32'd3235
; 
32'd140395: dataIn1 = 32'd3236
; 
32'd140396: dataIn1 = 32'd175
; 
32'd140397: dataIn1 = 32'd2004
; 
32'd140398: dataIn1 = 32'd2906
; 
32'd140399: dataIn1 = 32'd3230
; 
32'd140400: dataIn1 = 32'd3233
; 
32'd140401: dataIn1 = 32'd4307
; 
32'd140402: dataIn1 = 32'd4317
; 
32'd140403: dataIn1 = 32'd334
; 
32'd140404: dataIn1 = 32'd2004
; 
32'd140405: dataIn1 = 32'd2896
; 
32'd140406: dataIn1 = 32'd3231
; 
32'd140407: dataIn1 = 32'd3234
; 
32'd140408: dataIn1 = 32'd4304
; 
32'd140409: dataIn1 = 32'd4308
; 
32'd140410: dataIn1 = 32'd1779
; 
32'd140411: dataIn1 = 32'd2904
; 
32'd140412: dataIn1 = 32'd3232
; 
32'd140413: dataIn1 = 32'd3235
; 
32'd140414: dataIn1 = 32'd3236
; 
32'd140415: dataIn1 = 32'd11097
; 
32'd140416: dataIn1 = 32'd11098
; 
32'd140417: dataIn1 = 32'd1775
; 
32'd140418: dataIn1 = 32'd2894
; 
32'd140419: dataIn1 = 32'd3232
; 
32'd140420: dataIn1 = 32'd3235
; 
32'd140421: dataIn1 = 32'd3236
; 
32'd140422: dataIn1 = 32'd11096
; 
32'd140423: dataIn1 = 32'd11097
; 
32'd140424: dataIn1 = 32'd1780
; 
32'd140425: dataIn1 = 32'd2005
; 
32'd140426: dataIn1 = 32'd2905
; 
32'd140427: dataIn1 = 32'd3237
; 
32'd140428: dataIn1 = 32'd3238
; 
32'd140429: dataIn1 = 32'd3239
; 
32'd140430: dataIn1 = 32'd3240
; 
32'd140431: dataIn1 = 32'd1781
; 
32'd140432: dataIn1 = 32'd2005
; 
32'd140433: dataIn1 = 32'd2911
; 
32'd140434: dataIn1 = 32'd3237
; 
32'd140435: dataIn1 = 32'd3238
; 
32'd140436: dataIn1 = 32'd3239
; 
32'd140437: dataIn1 = 32'd3241
; 
32'd140438: dataIn1 = 32'd1780
; 
32'd140439: dataIn1 = 32'd1781
; 
32'd140440: dataIn1 = 32'd3237
; 
32'd140441: dataIn1 = 32'd3238
; 
32'd140442: dataIn1 = 32'd3239
; 
32'd140443: dataIn1 = 32'd3242
; 
32'd140444: dataIn1 = 32'd3243
; 
32'd140445: dataIn1 = 32'd175
; 
32'd140446: dataIn1 = 32'd2005
; 
32'd140447: dataIn1 = 32'd2905
; 
32'd140448: dataIn1 = 32'd3237
; 
32'd140449: dataIn1 = 32'd3240
; 
32'd140450: dataIn1 = 32'd4318
; 
32'd140451: dataIn1 = 32'd4331
; 
32'd140452: dataIn1 = 32'd341
; 
32'd140453: dataIn1 = 32'd2005
; 
32'd140454: dataIn1 = 32'd2911
; 
32'd140455: dataIn1 = 32'd3238
; 
32'd140456: dataIn1 = 32'd3241
; 
32'd140457: dataIn1 = 32'd4328
; 
32'd140458: dataIn1 = 32'd4332
; 
32'd140459: dataIn1 = 32'd1780
; 
32'd140460: dataIn1 = 32'd2903
; 
32'd140461: dataIn1 = 32'd3239
; 
32'd140462: dataIn1 = 32'd3242
; 
32'd140463: dataIn1 = 32'd3243
; 
32'd140464: dataIn1 = 32'd11100
; 
32'd140465: dataIn1 = 32'd11101
; 
32'd140466: dataIn1 = 32'd1781
; 
32'd140467: dataIn1 = 32'd2909
; 
32'd140468: dataIn1 = 32'd3239
; 
32'd140469: dataIn1 = 32'd3242
; 
32'd140470: dataIn1 = 32'd3243
; 
32'd140471: dataIn1 = 32'd11101
; 
32'd140472: dataIn1 = 32'd11102
; 
32'd140473: dataIn1 = 32'd1782
; 
32'd140474: dataIn1 = 32'd1789
; 
32'd140475: dataIn1 = 32'd3244
; 
32'd140476: dataIn1 = 32'd3245
; 
32'd140477: dataIn1 = 32'd3246
; 
32'd140478: dataIn1 = 32'd3247
; 
32'd140479: dataIn1 = 32'd3248
; 
32'd140480: dataIn1 = 32'd1782
; 
32'd140481: dataIn1 = 32'd2006
; 
32'd140482: dataIn1 = 32'd2910
; 
32'd140483: dataIn1 = 32'd3244
; 
32'd140484: dataIn1 = 32'd3245
; 
32'd140485: dataIn1 = 32'd3246
; 
32'd140486: dataIn1 = 32'd3249
; 
32'd140487: dataIn1 = 32'd1789
; 
32'd140488: dataIn1 = 32'd2006
; 
32'd140489: dataIn1 = 32'd2931
; 
32'd140490: dataIn1 = 32'd3244
; 
32'd140491: dataIn1 = 32'd3245
; 
32'd140492: dataIn1 = 32'd3246
; 
32'd140493: dataIn1 = 32'd3250
; 
32'd140494: dataIn1 = 32'd1782
; 
32'd140495: dataIn1 = 32'd2907
; 
32'd140496: dataIn1 = 32'd3244
; 
32'd140497: dataIn1 = 32'd3247
; 
32'd140498: dataIn1 = 32'd3248
; 
32'd140499: dataIn1 = 32'd11104
; 
32'd140500: dataIn1 = 32'd11105
; 
32'd140501: dataIn1 = 32'd1789
; 
32'd140502: dataIn1 = 32'd2929
; 
32'd140503: dataIn1 = 32'd3244
; 
32'd140504: dataIn1 = 32'd3247
; 
32'd140505: dataIn1 = 32'd3248
; 
32'd140506: dataIn1 = 32'd11105
; 
32'd140507: dataIn1 = 32'd11106
; 
32'd140508: dataIn1 = 32'd341
; 
32'd140509: dataIn1 = 32'd2006
; 
32'd140510: dataIn1 = 32'd2910
; 
32'd140511: dataIn1 = 32'd3245
; 
32'd140512: dataIn1 = 32'd3249
; 
32'd140513: dataIn1 = 32'd4327
; 
32'd140514: dataIn1 = 32'd4335
; 
32'd140515: dataIn1 = 32'd177
; 
32'd140516: dataIn1 = 32'd2006
; 
32'd140517: dataIn1 = 32'd2931
; 
32'd140518: dataIn1 = 32'd3246
; 
32'd140519: dataIn1 = 32'd3250
; 
32'd140520: dataIn1 = 32'd4336
; 
32'd140521: dataIn1 = 32'd4344
; 
32'd140522: dataIn1 = 32'd1784
; 
32'd140523: dataIn1 = 32'd2007
; 
32'd140524: dataIn1 = 32'd2915
; 
32'd140525: dataIn1 = 32'd3251
; 
32'd140526: dataIn1 = 32'd3252
; 
32'd140527: dataIn1 = 32'd3253
; 
32'd140528: dataIn1 = 32'd3254
; 
32'd140529: dataIn1 = 32'd1784
; 
32'd140530: dataIn1 = 32'd1793
; 
32'd140531: dataIn1 = 32'd3251
; 
32'd140532: dataIn1 = 32'd3252
; 
32'd140533: dataIn1 = 32'd3253
; 
32'd140534: dataIn1 = 32'd3255
; 
32'd140535: dataIn1 = 32'd3256
; 
32'd140536: dataIn1 = 32'd1793
; 
32'd140537: dataIn1 = 32'd2007
; 
32'd140538: dataIn1 = 32'd2941
; 
32'd140539: dataIn1 = 32'd3251
; 
32'd140540: dataIn1 = 32'd3252
; 
32'd140541: dataIn1 = 32'd3253
; 
32'd140542: dataIn1 = 32'd3257
; 
32'd140543: dataIn1 = 32'd343
; 
32'd140544: dataIn1 = 32'd2007
; 
32'd140545: dataIn1 = 32'd2915
; 
32'd140546: dataIn1 = 32'd3251
; 
32'd140547: dataIn1 = 32'd3254
; 
32'd140548: dataIn1 = 32'd4373
; 
32'd140549: dataIn1 = 32'd4382
; 
32'd140550: dataIn1 = 32'd1784
; 
32'd140551: dataIn1 = 32'd2913
; 
32'd140552: dataIn1 = 32'd3252
; 
32'd140553: dataIn1 = 32'd3255
; 
32'd140554: dataIn1 = 32'd3256
; 
32'd140555: dataIn1 = 32'd11120
; 
32'd140556: dataIn1 = 32'd11121
; 
32'd140557: dataIn1 = 32'd1793
; 
32'd140558: dataIn1 = 32'd2938
; 
32'd140559: dataIn1 = 32'd3252
; 
32'd140560: dataIn1 = 32'd3255
; 
32'd140561: dataIn1 = 32'd3256
; 
32'd140562: dataIn1 = 32'd11121
; 
32'd140563: dataIn1 = 32'd11122
; 
32'd140564: dataIn1 = 32'd180
; 
32'd140565: dataIn1 = 32'd2007
; 
32'd140566: dataIn1 = 32'd2941
; 
32'd140567: dataIn1 = 32'd3253
; 
32'd140568: dataIn1 = 32'd3257
; 
32'd140569: dataIn1 = 32'd4384
; 
32'd140570: dataIn1 = 32'd4393
; 
32'd140571: dataIn1 = 32'd1783
; 
32'd140572: dataIn1 = 32'd2008
; 
32'd140573: dataIn1 = 32'd2916
; 
32'd140574: dataIn1 = 32'd3258
; 
32'd140575: dataIn1 = 32'd3259
; 
32'd140576: dataIn1 = 32'd3260
; 
32'd140577: dataIn1 = 32'd3261
; 
32'd140578: dataIn1 = 32'd1787
; 
32'd140579: dataIn1 = 32'd2008
; 
32'd140580: dataIn1 = 32'd2926
; 
32'd140581: dataIn1 = 32'd3258
; 
32'd140582: dataIn1 = 32'd3259
; 
32'd140583: dataIn1 = 32'd3260
; 
32'd140584: dataIn1 = 32'd3262
; 
32'd140585: dataIn1 = 32'd1783
; 
32'd140586: dataIn1 = 32'd1787
; 
32'd140587: dataIn1 = 32'd3258
; 
32'd140588: dataIn1 = 32'd3259
; 
32'd140589: dataIn1 = 32'd3260
; 
32'd140590: dataIn1 = 32'd3263
; 
32'd140591: dataIn1 = 32'd3264
; 
32'd140592: dataIn1 = 32'd343
; 
32'd140593: dataIn1 = 32'd2008
; 
32'd140594: dataIn1 = 32'd2916
; 
32'd140595: dataIn1 = 32'd3258
; 
32'd140596: dataIn1 = 32'd3261
; 
32'd140597: dataIn1 = 32'd4374
; 
32'd140598: dataIn1 = 32'd4379
; 
32'd140599: dataIn1 = 32'd179
; 
32'd140600: dataIn1 = 32'd2008
; 
32'd140601: dataIn1 = 32'd2926
; 
32'd140602: dataIn1 = 32'd3259
; 
32'd140603: dataIn1 = 32'd3262
; 
32'd140604: dataIn1 = 32'd4367
; 
32'd140605: dataIn1 = 32'd4380
; 
32'd140606: dataIn1 = 32'd1783
; 
32'd140607: dataIn1 = 32'd2914
; 
32'd140608: dataIn1 = 32'd3260
; 
32'd140609: dataIn1 = 32'd3263
; 
32'd140610: dataIn1 = 32'd3264
; 
32'd140611: dataIn1 = 32'd11117
; 
32'd140612: dataIn1 = 32'd11118
; 
32'd140613: dataIn1 = 32'd1787
; 
32'd140614: dataIn1 = 32'd2924
; 
32'd140615: dataIn1 = 32'd3260
; 
32'd140616: dataIn1 = 32'd3263
; 
32'd140617: dataIn1 = 32'd3264
; 
32'd140618: dataIn1 = 32'd11116
; 
32'd140619: dataIn1 = 32'd11117
; 
32'd140620: dataIn1 = 32'd1786
; 
32'd140621: dataIn1 = 32'd1788
; 
32'd140622: dataIn1 = 32'd3265
; 
32'd140623: dataIn1 = 32'd3266
; 
32'd140624: dataIn1 = 32'd3267
; 
32'd140625: dataIn1 = 32'd3268
; 
32'd140626: dataIn1 = 32'd3269
; 
32'd140627: dataIn1 = 32'd1788
; 
32'd140628: dataIn1 = 32'd2009
; 
32'd140629: dataIn1 = 32'd2925
; 
32'd140630: dataIn1 = 32'd3265
; 
32'd140631: dataIn1 = 32'd3266
; 
32'd140632: dataIn1 = 32'd3267
; 
32'd140633: dataIn1 = 32'd3270
; 
32'd140634: dataIn1 = 32'd1786
; 
32'd140635: dataIn1 = 32'd2009
; 
32'd140636: dataIn1 = 32'd2920
; 
32'd140637: dataIn1 = 32'd3265
; 
32'd140638: dataIn1 = 32'd3266
; 
32'd140639: dataIn1 = 32'd3267
; 
32'd140640: dataIn1 = 32'd3271
; 
32'd140641: dataIn1 = 32'd1788
; 
32'd140642: dataIn1 = 32'd2922
; 
32'd140643: dataIn1 = 32'd3265
; 
32'd140644: dataIn1 = 32'd3268
; 
32'd140645: dataIn1 = 32'd3269
; 
32'd140646: dataIn1 = 32'd11113
; 
32'd140647: dataIn1 = 32'd11114
; 
32'd140648: dataIn1 = 32'd1786
; 
32'd140649: dataIn1 = 32'd2917
; 
32'd140650: dataIn1 = 32'd3265
; 
32'd140651: dataIn1 = 32'd3268
; 
32'd140652: dataIn1 = 32'd3269
; 
32'd140653: dataIn1 = 32'd11112
; 
32'd140654: dataIn1 = 32'd11113
; 
32'd140655: dataIn1 = 32'd179
; 
32'd140656: dataIn1 = 32'd2009
; 
32'd140657: dataIn1 = 32'd2925
; 
32'd140658: dataIn1 = 32'd3266
; 
32'd140659: dataIn1 = 32'd3270
; 
32'd140660: dataIn1 = 32'd4359
; 
32'd140661: dataIn1 = 32'd4366
; 
32'd140662: dataIn1 = 32'd349
; 
32'd140663: dataIn1 = 32'd2009
; 
32'd140664: dataIn1 = 32'd2920
; 
32'd140665: dataIn1 = 32'd3267
; 
32'd140666: dataIn1 = 32'd3271
; 
32'd140667: dataIn1 = 32'd4353
; 
32'd140668: dataIn1 = 32'd4360
; 
32'd140669: dataIn1 = 32'd1790
; 
32'd140670: dataIn1 = 32'd2010
; 
32'd140671: dataIn1 = 32'd2930
; 
32'd140672: dataIn1 = 32'd3272
; 
32'd140673: dataIn1 = 32'd3273
; 
32'd140674: dataIn1 = 32'd3274
; 
32'd140675: dataIn1 = 32'd3275
; 
32'd140676: dataIn1 = 32'd1785
; 
32'd140677: dataIn1 = 32'd1790
; 
32'd140678: dataIn1 = 32'd3272
; 
32'd140679: dataIn1 = 32'd3273
; 
32'd140680: dataIn1 = 32'd3274
; 
32'd140681: dataIn1 = 32'd3276
; 
32'd140682: dataIn1 = 32'd3277
; 
32'd140683: dataIn1 = 32'd1785
; 
32'd140684: dataIn1 = 32'd2010
; 
32'd140685: dataIn1 = 32'd2921
; 
32'd140686: dataIn1 = 32'd3272
; 
32'd140687: dataIn1 = 32'd3273
; 
32'd140688: dataIn1 = 32'd3274
; 
32'd140689: dataIn1 = 32'd3278
; 
32'd140690: dataIn1 = 32'd177
; 
32'd140691: dataIn1 = 32'd2010
; 
32'd140692: dataIn1 = 32'd2930
; 
32'd140693: dataIn1 = 32'd3272
; 
32'd140694: dataIn1 = 32'd3275
; 
32'd140695: dataIn1 = 32'd4345
; 
32'd140696: dataIn1 = 32'd4355
; 
32'd140697: dataIn1 = 32'd1790
; 
32'd140698: dataIn1 = 32'd2928
; 
32'd140699: dataIn1 = 32'd3273
; 
32'd140700: dataIn1 = 32'd3276
; 
32'd140701: dataIn1 = 32'd3277
; 
32'd140702: dataIn1 = 32'd11108
; 
32'd140703: dataIn1 = 32'd11109
; 
32'd140704: dataIn1 = 32'd1785
; 
32'd140705: dataIn1 = 32'd2918
; 
32'd140706: dataIn1 = 32'd3273
; 
32'd140707: dataIn1 = 32'd3276
; 
32'd140708: dataIn1 = 32'd3277
; 
32'd140709: dataIn1 = 32'd11109
; 
32'd140710: dataIn1 = 32'd11110
; 
32'd140711: dataIn1 = 32'd349
; 
32'd140712: dataIn1 = 32'd2010
; 
32'd140713: dataIn1 = 32'd2921
; 
32'd140714: dataIn1 = 32'd3274
; 
32'd140715: dataIn1 = 32'd3278
; 
32'd140716: dataIn1 = 32'd4354
; 
32'd140717: dataIn1 = 32'd4357
; 
32'd140718: dataIn1 = 32'd1792
; 
32'd140719: dataIn1 = 32'd1794
; 
32'd140720: dataIn1 = 32'd3279
; 
32'd140721: dataIn1 = 32'd3280
; 
32'd140722: dataIn1 = 32'd3281
; 
32'd140723: dataIn1 = 32'd3282
; 
32'd140724: dataIn1 = 32'd3283
; 
32'd140725: dataIn1 = 32'd1792
; 
32'd140726: dataIn1 = 32'd2011
; 
32'd140727: dataIn1 = 32'd2935
; 
32'd140728: dataIn1 = 32'd3279
; 
32'd140729: dataIn1 = 32'd3280
; 
32'd140730: dataIn1 = 32'd3281
; 
32'd140731: dataIn1 = 32'd3284
; 
32'd140732: dataIn1 = 32'd1794
; 
32'd140733: dataIn1 = 32'd2011
; 
32'd140734: dataIn1 = 32'd2940
; 
32'd140735: dataIn1 = 32'd3279
; 
32'd140736: dataIn1 = 32'd3280
; 
32'd140737: dataIn1 = 32'd3281
; 
32'd140738: dataIn1 = 32'd3285
; 
32'd140739: dataIn1 = 32'd1792
; 
32'd140740: dataIn1 = 32'd2932
; 
32'd140741: dataIn1 = 32'd3279
; 
32'd140742: dataIn1 = 32'd3282
; 
32'd140743: dataIn1 = 32'd3283
; 
32'd140744: dataIn1 = 32'd11125
; 
32'd140745: dataIn1 = 32'd11126
; 
32'd140746: dataIn1 = 32'd1794
; 
32'd140747: dataIn1 = 32'd2937
; 
32'd140748: dataIn1 = 32'd3279
; 
32'd140749: dataIn1 = 32'd3282
; 
32'd140750: dataIn1 = 32'd3283
; 
32'd140751: dataIn1 = 32'd11124
; 
32'd140752: dataIn1 = 32'd11125
; 
32'd140753: dataIn1 = 32'd350
; 
32'd140754: dataIn1 = 32'd2011
; 
32'd140755: dataIn1 = 32'd2935
; 
32'd140756: dataIn1 = 32'd3280
; 
32'd140757: dataIn1 = 32'd3284
; 
32'd140758: dataIn1 = 32'd4399
; 
32'd140759: dataIn1 = 32'd4408
; 
32'd140760: dataIn1 = 32'd180
; 
32'd140761: dataIn1 = 32'd2011
; 
32'd140762: dataIn1 = 32'd2940
; 
32'd140763: dataIn1 = 32'd3281
; 
32'd140764: dataIn1 = 32'd3285
; 
32'd140765: dataIn1 = 32'd4392
; 
32'd140766: dataIn1 = 32'd4409
; 
32'd140767: dataIn1 = 32'd1795
; 
32'd140768: dataIn1 = 32'd2012
; 
32'd140769: dataIn1 = 32'd2946
; 
32'd140770: dataIn1 = 32'd3286
; 
32'd140771: dataIn1 = 32'd3287
; 
32'd140772: dataIn1 = 32'd3288
; 
32'd140773: dataIn1 = 32'd3289
; 
32'd140774: dataIn1 = 32'd1791
; 
32'd140775: dataIn1 = 32'd2012
; 
32'd140776: dataIn1 = 32'd2936
; 
32'd140777: dataIn1 = 32'd3286
; 
32'd140778: dataIn1 = 32'd3287
; 
32'd140779: dataIn1 = 32'd3288
; 
32'd140780: dataIn1 = 32'd3290
; 
32'd140781: dataIn1 = 32'd1791
; 
32'd140782: dataIn1 = 32'd1795
; 
32'd140783: dataIn1 = 32'd3286
; 
32'd140784: dataIn1 = 32'd3287
; 
32'd140785: dataIn1 = 32'd3288
; 
32'd140786: dataIn1 = 32'd3291
; 
32'd140787: dataIn1 = 32'd3292
; 
32'd140788: dataIn1 = 32'd181
; 
32'd140789: dataIn1 = 32'd2012
; 
32'd140790: dataIn1 = 32'd2946
; 
32'd140791: dataIn1 = 32'd3286
; 
32'd140792: dataIn1 = 32'd3289
; 
32'd140793: dataIn1 = 32'd4403
; 
32'd140794: dataIn1 = 32'd4413
; 
32'd140795: dataIn1 = 32'd350
; 
32'd140796: dataIn1 = 32'd2012
; 
32'd140797: dataIn1 = 32'd2936
; 
32'd140798: dataIn1 = 32'd3287
; 
32'd140799: dataIn1 = 32'd3290
; 
32'd140800: dataIn1 = 32'd4400
; 
32'd140801: dataIn1 = 32'd4404
; 
32'd140802: dataIn1 = 32'd1795
; 
32'd140803: dataIn1 = 32'd2944
; 
32'd140804: dataIn1 = 32'd3288
; 
32'd140805: dataIn1 = 32'd3291
; 
32'd140806: dataIn1 = 32'd3292
; 
32'd140807: dataIn1 = 32'd11129
; 
32'd140808: dataIn1 = 32'd11130
; 
32'd140809: dataIn1 = 32'd1791
; 
32'd140810: dataIn1 = 32'd2934
; 
32'd140811: dataIn1 = 32'd3288
; 
32'd140812: dataIn1 = 32'd3291
; 
32'd140813: dataIn1 = 32'd3292
; 
32'd140814: dataIn1 = 32'd11128
; 
32'd140815: dataIn1 = 32'd11129
; 
32'd140816: dataIn1 = 32'd1796
; 
32'd140817: dataIn1 = 32'd2013
; 
32'd140818: dataIn1 = 32'd2945
; 
32'd140819: dataIn1 = 32'd3293
; 
32'd140820: dataIn1 = 32'd3294
; 
32'd140821: dataIn1 = 32'd3295
; 
32'd140822: dataIn1 = 32'd3296
; 
32'd140823: dataIn1 = 32'd1797
; 
32'd140824: dataIn1 = 32'd2013
; 
32'd140825: dataIn1 = 32'd2951
; 
32'd140826: dataIn1 = 32'd3293
; 
32'd140827: dataIn1 = 32'd3294
; 
32'd140828: dataIn1 = 32'd3295
; 
32'd140829: dataIn1 = 32'd3297
; 
32'd140830: dataIn1 = 32'd1796
; 
32'd140831: dataIn1 = 32'd1797
; 
32'd140832: dataIn1 = 32'd3293
; 
32'd140833: dataIn1 = 32'd3294
; 
32'd140834: dataIn1 = 32'd3295
; 
32'd140835: dataIn1 = 32'd3298
; 
32'd140836: dataIn1 = 32'd3299
; 
32'd140837: dataIn1 = 32'd181
; 
32'd140838: dataIn1 = 32'd2013
; 
32'd140839: dataIn1 = 32'd2945
; 
32'd140840: dataIn1 = 32'd3293
; 
32'd140841: dataIn1 = 32'd3296
; 
32'd140842: dataIn1 = 32'd4414
; 
32'd140843: dataIn1 = 32'd4427
; 
32'd140844: dataIn1 = 32'd357
; 
32'd140845: dataIn1 = 32'd2013
; 
32'd140846: dataIn1 = 32'd2951
; 
32'd140847: dataIn1 = 32'd3294
; 
32'd140848: dataIn1 = 32'd3297
; 
32'd140849: dataIn1 = 32'd4424
; 
32'd140850: dataIn1 = 32'd4428
; 
32'd140851: dataIn1 = 32'd1796
; 
32'd140852: dataIn1 = 32'd2943
; 
32'd140853: dataIn1 = 32'd3295
; 
32'd140854: dataIn1 = 32'd3298
; 
32'd140855: dataIn1 = 32'd3299
; 
32'd140856: dataIn1 = 32'd11132
; 
32'd140857: dataIn1 = 32'd11133
; 
32'd140858: dataIn1 = 32'd1797
; 
32'd140859: dataIn1 = 32'd2949
; 
32'd140860: dataIn1 = 32'd3295
; 
32'd140861: dataIn1 = 32'd3298
; 
32'd140862: dataIn1 = 32'd3299
; 
32'd140863: dataIn1 = 32'd11133
; 
32'd140864: dataIn1 = 32'd11134
; 
32'd140865: dataIn1 = 32'd1798
; 
32'd140866: dataIn1 = 32'd1805
; 
32'd140867: dataIn1 = 32'd3300
; 
32'd140868: dataIn1 = 32'd3301
; 
32'd140869: dataIn1 = 32'd3302
; 
32'd140870: dataIn1 = 32'd3303
; 
32'd140871: dataIn1 = 32'd3304
; 
32'd140872: dataIn1 = 32'd1798
; 
32'd140873: dataIn1 = 32'd2014
; 
32'd140874: dataIn1 = 32'd2950
; 
32'd140875: dataIn1 = 32'd3300
; 
32'd140876: dataIn1 = 32'd3301
; 
32'd140877: dataIn1 = 32'd3302
; 
32'd140878: dataIn1 = 32'd3305
; 
32'd140879: dataIn1 = 32'd1805
; 
32'd140880: dataIn1 = 32'd2014
; 
32'd140881: dataIn1 = 32'd2971
; 
32'd140882: dataIn1 = 32'd3300
; 
32'd140883: dataIn1 = 32'd3301
; 
32'd140884: dataIn1 = 32'd3302
; 
32'd140885: dataIn1 = 32'd3306
; 
32'd140886: dataIn1 = 32'd1798
; 
32'd140887: dataIn1 = 32'd2947
; 
32'd140888: dataIn1 = 32'd3300
; 
32'd140889: dataIn1 = 32'd3303
; 
32'd140890: dataIn1 = 32'd3304
; 
32'd140891: dataIn1 = 32'd11136
; 
32'd140892: dataIn1 = 32'd11137
; 
32'd140893: dataIn1 = 32'd1805
; 
32'd140894: dataIn1 = 32'd2969
; 
32'd140895: dataIn1 = 32'd3300
; 
32'd140896: dataIn1 = 32'd3303
; 
32'd140897: dataIn1 = 32'd3304
; 
32'd140898: dataIn1 = 32'd11137
; 
32'd140899: dataIn1 = 32'd11138
; 
32'd140900: dataIn1 = 32'd357
; 
32'd140901: dataIn1 = 32'd2014
; 
32'd140902: dataIn1 = 32'd2950
; 
32'd140903: dataIn1 = 32'd3301
; 
32'd140904: dataIn1 = 32'd3305
; 
32'd140905: dataIn1 = 32'd4423
; 
32'd140906: dataIn1 = 32'd4431
; 
32'd140907: dataIn1 = 32'd183
; 
32'd140908: dataIn1 = 32'd2014
; 
32'd140909: dataIn1 = 32'd2971
; 
32'd140910: dataIn1 = 32'd3302
; 
32'd140911: dataIn1 = 32'd3306
; 
32'd140912: dataIn1 = 32'd4432
; 
32'd140913: dataIn1 = 32'd4440
; 
32'd140914: dataIn1 = 32'd1800
; 
32'd140915: dataIn1 = 32'd2015
; 
32'd140916: dataIn1 = 32'd2955
; 
32'd140917: dataIn1 = 32'd3307
; 
32'd140918: dataIn1 = 32'd3308
; 
32'd140919: dataIn1 = 32'd3309
; 
32'd140920: dataIn1 = 32'd3310
; 
32'd140921: dataIn1 = 32'd1800
; 
32'd140922: dataIn1 = 32'd1809
; 
32'd140923: dataIn1 = 32'd3307
; 
32'd140924: dataIn1 = 32'd3308
; 
32'd140925: dataIn1 = 32'd3309
; 
32'd140926: dataIn1 = 32'd3311
; 
32'd140927: dataIn1 = 32'd3312
; 
32'd140928: dataIn1 = 32'd1809
; 
32'd140929: dataIn1 = 32'd2015
; 
32'd140930: dataIn1 = 32'd2981
; 
32'd140931: dataIn1 = 32'd3307
; 
32'd140932: dataIn1 = 32'd3308
; 
32'd140933: dataIn1 = 32'd3309
; 
32'd140934: dataIn1 = 32'd3313
; 
32'd140935: dataIn1 = 32'd359
; 
32'd140936: dataIn1 = 32'd2015
; 
32'd140937: dataIn1 = 32'd2955
; 
32'd140938: dataIn1 = 32'd3307
; 
32'd140939: dataIn1 = 32'd3310
; 
32'd140940: dataIn1 = 32'd4469
; 
32'd140941: dataIn1 = 32'd4478
; 
32'd140942: dataIn1 = 32'd1800
; 
32'd140943: dataIn1 = 32'd2953
; 
32'd140944: dataIn1 = 32'd3308
; 
32'd140945: dataIn1 = 32'd3311
; 
32'd140946: dataIn1 = 32'd3312
; 
32'd140947: dataIn1 = 32'd11152
; 
32'd140948: dataIn1 = 32'd11153
; 
32'd140949: dataIn1 = 32'd1809
; 
32'd140950: dataIn1 = 32'd2978
; 
32'd140951: dataIn1 = 32'd3308
; 
32'd140952: dataIn1 = 32'd3311
; 
32'd140953: dataIn1 = 32'd3312
; 
32'd140954: dataIn1 = 32'd11153
; 
32'd140955: dataIn1 = 32'd11154
; 
32'd140956: dataIn1 = 32'd186
; 
32'd140957: dataIn1 = 32'd2015
; 
32'd140958: dataIn1 = 32'd2981
; 
32'd140959: dataIn1 = 32'd3309
; 
32'd140960: dataIn1 = 32'd3313
; 
32'd140961: dataIn1 = 32'd4480
; 
32'd140962: dataIn1 = 32'd4489
; 
32'd140963: dataIn1 = 32'd1799
; 
32'd140964: dataIn1 = 32'd2016
; 
32'd140965: dataIn1 = 32'd2956
; 
32'd140966: dataIn1 = 32'd3314
; 
32'd140967: dataIn1 = 32'd3315
; 
32'd140968: dataIn1 = 32'd3316
; 
32'd140969: dataIn1 = 32'd3317
; 
32'd140970: dataIn1 = 32'd1803
; 
32'd140971: dataIn1 = 32'd2016
; 
32'd140972: dataIn1 = 32'd2966
; 
32'd140973: dataIn1 = 32'd3314
; 
32'd140974: dataIn1 = 32'd3315
; 
32'd140975: dataIn1 = 32'd3316
; 
32'd140976: dataIn1 = 32'd3318
; 
32'd140977: dataIn1 = 32'd1799
; 
32'd140978: dataIn1 = 32'd1803
; 
32'd140979: dataIn1 = 32'd3314
; 
32'd140980: dataIn1 = 32'd3315
; 
32'd140981: dataIn1 = 32'd3316
; 
32'd140982: dataIn1 = 32'd3319
; 
32'd140983: dataIn1 = 32'd3320
; 
32'd140984: dataIn1 = 32'd359
; 
32'd140985: dataIn1 = 32'd2016
; 
32'd140986: dataIn1 = 32'd2956
; 
32'd140987: dataIn1 = 32'd3314
; 
32'd140988: dataIn1 = 32'd3317
; 
32'd140989: dataIn1 = 32'd4470
; 
32'd140990: dataIn1 = 32'd4475
; 
32'd140991: dataIn1 = 32'd185
; 
32'd140992: dataIn1 = 32'd2016
; 
32'd140993: dataIn1 = 32'd2966
; 
32'd140994: dataIn1 = 32'd3315
; 
32'd140995: dataIn1 = 32'd3318
; 
32'd140996: dataIn1 = 32'd4463
; 
32'd140997: dataIn1 = 32'd4476
; 
32'd140998: dataIn1 = 32'd1799
; 
32'd140999: dataIn1 = 32'd2954
; 
32'd141000: dataIn1 = 32'd3316
; 
32'd141001: dataIn1 = 32'd3319
; 
32'd141002: dataIn1 = 32'd3320
; 
32'd141003: dataIn1 = 32'd11149
; 
32'd141004: dataIn1 = 32'd11150
; 
32'd141005: dataIn1 = 32'd1803
; 
32'd141006: dataIn1 = 32'd2964
; 
32'd141007: dataIn1 = 32'd3316
; 
32'd141008: dataIn1 = 32'd3319
; 
32'd141009: dataIn1 = 32'd3320
; 
32'd141010: dataIn1 = 32'd11148
; 
32'd141011: dataIn1 = 32'd11149
; 
32'd141012: dataIn1 = 32'd1802
; 
32'd141013: dataIn1 = 32'd1804
; 
32'd141014: dataIn1 = 32'd3321
; 
32'd141015: dataIn1 = 32'd3322
; 
32'd141016: dataIn1 = 32'd3323
; 
32'd141017: dataIn1 = 32'd3324
; 
32'd141018: dataIn1 = 32'd3325
; 
32'd141019: dataIn1 = 32'd1804
; 
32'd141020: dataIn1 = 32'd2017
; 
32'd141021: dataIn1 = 32'd2965
; 
32'd141022: dataIn1 = 32'd3321
; 
32'd141023: dataIn1 = 32'd3322
; 
32'd141024: dataIn1 = 32'd3323
; 
32'd141025: dataIn1 = 32'd3326
; 
32'd141026: dataIn1 = 32'd1802
; 
32'd141027: dataIn1 = 32'd2017
; 
32'd141028: dataIn1 = 32'd2960
; 
32'd141029: dataIn1 = 32'd3321
; 
32'd141030: dataIn1 = 32'd3322
; 
32'd141031: dataIn1 = 32'd3323
; 
32'd141032: dataIn1 = 32'd3327
; 
32'd141033: dataIn1 = 32'd1804
; 
32'd141034: dataIn1 = 32'd2962
; 
32'd141035: dataIn1 = 32'd3321
; 
32'd141036: dataIn1 = 32'd3324
; 
32'd141037: dataIn1 = 32'd3325
; 
32'd141038: dataIn1 = 32'd11145
; 
32'd141039: dataIn1 = 32'd11146
; 
32'd141040: dataIn1 = 32'd1802
; 
32'd141041: dataIn1 = 32'd2957
; 
32'd141042: dataIn1 = 32'd3321
; 
32'd141043: dataIn1 = 32'd3324
; 
32'd141044: dataIn1 = 32'd3325
; 
32'd141045: dataIn1 = 32'd11144
; 
32'd141046: dataIn1 = 32'd11145
; 
32'd141047: dataIn1 = 32'd185
; 
32'd141048: dataIn1 = 32'd2017
; 
32'd141049: dataIn1 = 32'd2965
; 
32'd141050: dataIn1 = 32'd3322
; 
32'd141051: dataIn1 = 32'd3326
; 
32'd141052: dataIn1 = 32'd4455
; 
32'd141053: dataIn1 = 32'd4462
; 
32'd141054: dataIn1 = 32'd365
; 
32'd141055: dataIn1 = 32'd2017
; 
32'd141056: dataIn1 = 32'd2960
; 
32'd141057: dataIn1 = 32'd3323
; 
32'd141058: dataIn1 = 32'd3327
; 
32'd141059: dataIn1 = 32'd4449
; 
32'd141060: dataIn1 = 32'd4456
; 
32'd141061: dataIn1 = 32'd1806
; 
32'd141062: dataIn1 = 32'd2018
; 
32'd141063: dataIn1 = 32'd2970
; 
32'd141064: dataIn1 = 32'd3328
; 
32'd141065: dataIn1 = 32'd3329
; 
32'd141066: dataIn1 = 32'd3330
; 
32'd141067: dataIn1 = 32'd3331
; 
32'd141068: dataIn1 = 32'd1801
; 
32'd141069: dataIn1 = 32'd1806
; 
32'd141070: dataIn1 = 32'd3328
; 
32'd141071: dataIn1 = 32'd3329
; 
32'd141072: dataIn1 = 32'd3330
; 
32'd141073: dataIn1 = 32'd3332
; 
32'd141074: dataIn1 = 32'd3333
; 
32'd141075: dataIn1 = 32'd1801
; 
32'd141076: dataIn1 = 32'd2018
; 
32'd141077: dataIn1 = 32'd2961
; 
32'd141078: dataIn1 = 32'd3328
; 
32'd141079: dataIn1 = 32'd3329
; 
32'd141080: dataIn1 = 32'd3330
; 
32'd141081: dataIn1 = 32'd3334
; 
32'd141082: dataIn1 = 32'd183
; 
32'd141083: dataIn1 = 32'd2018
; 
32'd141084: dataIn1 = 32'd2970
; 
32'd141085: dataIn1 = 32'd3328
; 
32'd141086: dataIn1 = 32'd3331
; 
32'd141087: dataIn1 = 32'd4441
; 
32'd141088: dataIn1 = 32'd4451
; 
32'd141089: dataIn1 = 32'd1806
; 
32'd141090: dataIn1 = 32'd2968
; 
32'd141091: dataIn1 = 32'd3329
; 
32'd141092: dataIn1 = 32'd3332
; 
32'd141093: dataIn1 = 32'd3333
; 
32'd141094: dataIn1 = 32'd11140
; 
32'd141095: dataIn1 = 32'd11141
; 
32'd141096: dataIn1 = 32'd1801
; 
32'd141097: dataIn1 = 32'd2958
; 
32'd141098: dataIn1 = 32'd3329
; 
32'd141099: dataIn1 = 32'd3332
; 
32'd141100: dataIn1 = 32'd3333
; 
32'd141101: dataIn1 = 32'd11141
; 
32'd141102: dataIn1 = 32'd11142
; 
32'd141103: dataIn1 = 32'd365
; 
32'd141104: dataIn1 = 32'd2018
; 
32'd141105: dataIn1 = 32'd2961
; 
32'd141106: dataIn1 = 32'd3330
; 
32'd141107: dataIn1 = 32'd3334
; 
32'd141108: dataIn1 = 32'd4450
; 
32'd141109: dataIn1 = 32'd4453
; 
32'd141110: dataIn1 = 32'd1808
; 
32'd141111: dataIn1 = 32'd1810
; 
32'd141112: dataIn1 = 32'd3335
; 
32'd141113: dataIn1 = 32'd3336
; 
32'd141114: dataIn1 = 32'd3337
; 
32'd141115: dataIn1 = 32'd3338
; 
32'd141116: dataIn1 = 32'd3339
; 
32'd141117: dataIn1 = 32'd1808
; 
32'd141118: dataIn1 = 32'd2019
; 
32'd141119: dataIn1 = 32'd2975
; 
32'd141120: dataIn1 = 32'd3335
; 
32'd141121: dataIn1 = 32'd3336
; 
32'd141122: dataIn1 = 32'd3337
; 
32'd141123: dataIn1 = 32'd3340
; 
32'd141124: dataIn1 = 32'd1810
; 
32'd141125: dataIn1 = 32'd2019
; 
32'd141126: dataIn1 = 32'd2980
; 
32'd141127: dataIn1 = 32'd3335
; 
32'd141128: dataIn1 = 32'd3336
; 
32'd141129: dataIn1 = 32'd3337
; 
32'd141130: dataIn1 = 32'd3341
; 
32'd141131: dataIn1 = 32'd1808
; 
32'd141132: dataIn1 = 32'd2972
; 
32'd141133: dataIn1 = 32'd3335
; 
32'd141134: dataIn1 = 32'd3338
; 
32'd141135: dataIn1 = 32'd3339
; 
32'd141136: dataIn1 = 32'd11157
; 
32'd141137: dataIn1 = 32'd11158
; 
32'd141138: dataIn1 = 32'd1810
; 
32'd141139: dataIn1 = 32'd2977
; 
32'd141140: dataIn1 = 32'd3335
; 
32'd141141: dataIn1 = 32'd3338
; 
32'd141142: dataIn1 = 32'd3339
; 
32'd141143: dataIn1 = 32'd11156
; 
32'd141144: dataIn1 = 32'd11157
; 
32'd141145: dataIn1 = 32'd366
; 
32'd141146: dataIn1 = 32'd2019
; 
32'd141147: dataIn1 = 32'd2975
; 
32'd141148: dataIn1 = 32'd3336
; 
32'd141149: dataIn1 = 32'd3340
; 
32'd141150: dataIn1 = 32'd4495
; 
32'd141151: dataIn1 = 32'd4504
; 
32'd141152: dataIn1 = 32'd186
; 
32'd141153: dataIn1 = 32'd2019
; 
32'd141154: dataIn1 = 32'd2980
; 
32'd141155: dataIn1 = 32'd3337
; 
32'd141156: dataIn1 = 32'd3341
; 
32'd141157: dataIn1 = 32'd4488
; 
32'd141158: dataIn1 = 32'd4505
; 
32'd141159: dataIn1 = 32'd1811
; 
32'd141160: dataIn1 = 32'd2020
; 
32'd141161: dataIn1 = 32'd2986
; 
32'd141162: dataIn1 = 32'd3342
; 
32'd141163: dataIn1 = 32'd3343
; 
32'd141164: dataIn1 = 32'd3344
; 
32'd141165: dataIn1 = 32'd3345
; 
32'd141166: dataIn1 = 32'd1807
; 
32'd141167: dataIn1 = 32'd2020
; 
32'd141168: dataIn1 = 32'd2976
; 
32'd141169: dataIn1 = 32'd3342
; 
32'd141170: dataIn1 = 32'd3343
; 
32'd141171: dataIn1 = 32'd3344
; 
32'd141172: dataIn1 = 32'd3346
; 
32'd141173: dataIn1 = 32'd1807
; 
32'd141174: dataIn1 = 32'd1811
; 
32'd141175: dataIn1 = 32'd3342
; 
32'd141176: dataIn1 = 32'd3343
; 
32'd141177: dataIn1 = 32'd3344
; 
32'd141178: dataIn1 = 32'd3347
; 
32'd141179: dataIn1 = 32'd3348
; 
32'd141180: dataIn1 = 32'd187
; 
32'd141181: dataIn1 = 32'd2020
; 
32'd141182: dataIn1 = 32'd2986
; 
32'd141183: dataIn1 = 32'd3342
; 
32'd141184: dataIn1 = 32'd3345
; 
32'd141185: dataIn1 = 32'd4499
; 
32'd141186: dataIn1 = 32'd4509
; 
32'd141187: dataIn1 = 32'd366
; 
32'd141188: dataIn1 = 32'd2020
; 
32'd141189: dataIn1 = 32'd2976
; 
32'd141190: dataIn1 = 32'd3343
; 
32'd141191: dataIn1 = 32'd3346
; 
32'd141192: dataIn1 = 32'd4496
; 
32'd141193: dataIn1 = 32'd4500
; 
32'd141194: dataIn1 = 32'd1811
; 
32'd141195: dataIn1 = 32'd2984
; 
32'd141196: dataIn1 = 32'd3344
; 
32'd141197: dataIn1 = 32'd3347
; 
32'd141198: dataIn1 = 32'd3348
; 
32'd141199: dataIn1 = 32'd11161
; 
32'd141200: dataIn1 = 32'd11162
; 
32'd141201: dataIn1 = 32'd1807
; 
32'd141202: dataIn1 = 32'd2974
; 
32'd141203: dataIn1 = 32'd3344
; 
32'd141204: dataIn1 = 32'd3347
; 
32'd141205: dataIn1 = 32'd3348
; 
32'd141206: dataIn1 = 32'd11160
; 
32'd141207: dataIn1 = 32'd11161
; 
32'd141208: dataIn1 = 32'd1812
; 
32'd141209: dataIn1 = 32'd2021
; 
32'd141210: dataIn1 = 32'd2985
; 
32'd141211: dataIn1 = 32'd3349
; 
32'd141212: dataIn1 = 32'd3350
; 
32'd141213: dataIn1 = 32'd3351
; 
32'd141214: dataIn1 = 32'd3352
; 
32'd141215: dataIn1 = 32'd1813
; 
32'd141216: dataIn1 = 32'd2021
; 
32'd141217: dataIn1 = 32'd2991
; 
32'd141218: dataIn1 = 32'd3349
; 
32'd141219: dataIn1 = 32'd3350
; 
32'd141220: dataIn1 = 32'd3351
; 
32'd141221: dataIn1 = 32'd3353
; 
32'd141222: dataIn1 = 32'd1812
; 
32'd141223: dataIn1 = 32'd1813
; 
32'd141224: dataIn1 = 32'd3349
; 
32'd141225: dataIn1 = 32'd3350
; 
32'd141226: dataIn1 = 32'd3351
; 
32'd141227: dataIn1 = 32'd3354
; 
32'd141228: dataIn1 = 32'd3355
; 
32'd141229: dataIn1 = 32'd187
; 
32'd141230: dataIn1 = 32'd2021
; 
32'd141231: dataIn1 = 32'd2985
; 
32'd141232: dataIn1 = 32'd3349
; 
32'd141233: dataIn1 = 32'd3352
; 
32'd141234: dataIn1 = 32'd4510
; 
32'd141235: dataIn1 = 32'd4523
; 
32'd141236: dataIn1 = 32'd373
; 
32'd141237: dataIn1 = 32'd2021
; 
32'd141238: dataIn1 = 32'd2991
; 
32'd141239: dataIn1 = 32'd3350
; 
32'd141240: dataIn1 = 32'd3353
; 
32'd141241: dataIn1 = 32'd4520
; 
32'd141242: dataIn1 = 32'd4524
; 
32'd141243: dataIn1 = 32'd1812
; 
32'd141244: dataIn1 = 32'd2983
; 
32'd141245: dataIn1 = 32'd3351
; 
32'd141246: dataIn1 = 32'd3354
; 
32'd141247: dataIn1 = 32'd3355
; 
32'd141248: dataIn1 = 32'd11164
; 
32'd141249: dataIn1 = 32'd11165
; 
32'd141250: dataIn1 = 32'd1813
; 
32'd141251: dataIn1 = 32'd2989
; 
32'd141252: dataIn1 = 32'd3351
; 
32'd141253: dataIn1 = 32'd3354
; 
32'd141254: dataIn1 = 32'd3355
; 
32'd141255: dataIn1 = 32'd11165
; 
32'd141256: dataIn1 = 32'd11166
; 
32'd141257: dataIn1 = 32'd1814
; 
32'd141258: dataIn1 = 32'd1821
; 
32'd141259: dataIn1 = 32'd3356
; 
32'd141260: dataIn1 = 32'd3357
; 
32'd141261: dataIn1 = 32'd3358
; 
32'd141262: dataIn1 = 32'd3359
; 
32'd141263: dataIn1 = 32'd3360
; 
32'd141264: dataIn1 = 32'd1814
; 
32'd141265: dataIn1 = 32'd2022
; 
32'd141266: dataIn1 = 32'd2990
; 
32'd141267: dataIn1 = 32'd3356
; 
32'd141268: dataIn1 = 32'd3357
; 
32'd141269: dataIn1 = 32'd3358
; 
32'd141270: dataIn1 = 32'd3361
; 
32'd141271: dataIn1 = 32'd1821
; 
32'd141272: dataIn1 = 32'd2022
; 
32'd141273: dataIn1 = 32'd3011
; 
32'd141274: dataIn1 = 32'd3356
; 
32'd141275: dataIn1 = 32'd3357
; 
32'd141276: dataIn1 = 32'd3358
; 
32'd141277: dataIn1 = 32'd3362
; 
32'd141278: dataIn1 = 32'd1814
; 
32'd141279: dataIn1 = 32'd2987
; 
32'd141280: dataIn1 = 32'd3356
; 
32'd141281: dataIn1 = 32'd3359
; 
32'd141282: dataIn1 = 32'd3360
; 
32'd141283: dataIn1 = 32'd11168
; 
32'd141284: dataIn1 = 32'd11169
; 
32'd141285: dataIn1 = 32'd1821
; 
32'd141286: dataIn1 = 32'd3009
; 
32'd141287: dataIn1 = 32'd3356
; 
32'd141288: dataIn1 = 32'd3359
; 
32'd141289: dataIn1 = 32'd3360
; 
32'd141290: dataIn1 = 32'd11169
; 
32'd141291: dataIn1 = 32'd11170
; 
32'd141292: dataIn1 = 32'd11171
; 
32'd141293: dataIn1 = 32'd373
; 
32'd141294: dataIn1 = 32'd2022
; 
32'd141295: dataIn1 = 32'd2990
; 
32'd141296: dataIn1 = 32'd3357
; 
32'd141297: dataIn1 = 32'd3361
; 
32'd141298: dataIn1 = 32'd4519
; 
32'd141299: dataIn1 = 32'd4527
; 
32'd141300: dataIn1 = 32'd189
; 
32'd141301: dataIn1 = 32'd2022
; 
32'd141302: dataIn1 = 32'd3011
; 
32'd141303: dataIn1 = 32'd3358
; 
32'd141304: dataIn1 = 32'd3362
; 
32'd141305: dataIn1 = 32'd4528
; 
32'd141306: dataIn1 = 32'd4536
; 
32'd141307: dataIn1 = 32'd1816
; 
32'd141308: dataIn1 = 32'd2023
; 
32'd141309: dataIn1 = 32'd2995
; 
32'd141310: dataIn1 = 32'd3363
; 
32'd141311: dataIn1 = 32'd3364
; 
32'd141312: dataIn1 = 32'd3365
; 
32'd141313: dataIn1 = 32'd3366
; 
32'd141314: dataIn1 = 32'd1816
; 
32'd141315: dataIn1 = 32'd1825
; 
32'd141316: dataIn1 = 32'd3363
; 
32'd141317: dataIn1 = 32'd3364
; 
32'd141318: dataIn1 = 32'd3365
; 
32'd141319: dataIn1 = 32'd3367
; 
32'd141320: dataIn1 = 32'd3368
; 
32'd141321: dataIn1 = 32'd1825
; 
32'd141322: dataIn1 = 32'd2023
; 
32'd141323: dataIn1 = 32'd3021
; 
32'd141324: dataIn1 = 32'd3363
; 
32'd141325: dataIn1 = 32'd3364
; 
32'd141326: dataIn1 = 32'd3365
; 
32'd141327: dataIn1 = 32'd3369
; 
32'd141328: dataIn1 = 32'd375
; 
32'd141329: dataIn1 = 32'd2023
; 
32'd141330: dataIn1 = 32'd2995
; 
32'd141331: dataIn1 = 32'd3363
; 
32'd141332: dataIn1 = 32'd3366
; 
32'd141333: dataIn1 = 32'd4565
; 
32'd141334: dataIn1 = 32'd4574
; 
32'd141335: dataIn1 = 32'd1816
; 
32'd141336: dataIn1 = 32'd2993
; 
32'd141337: dataIn1 = 32'd3364
; 
32'd141338: dataIn1 = 32'd3367
; 
32'd141339: dataIn1 = 32'd3368
; 
32'd141340: dataIn1 = 32'd11185
; 
32'd141341: dataIn1 = 32'd11186
; 
32'd141342: dataIn1 = 32'd1825
; 
32'd141343: dataIn1 = 32'd3018
; 
32'd141344: dataIn1 = 32'd3364
; 
32'd141345: dataIn1 = 32'd3367
; 
32'd141346: dataIn1 = 32'd3368
; 
32'd141347: dataIn1 = 32'd11186
; 
32'd141348: dataIn1 = 32'd11187
; 
32'd141349: dataIn1 = 32'd192
; 
32'd141350: dataIn1 = 32'd2023
; 
32'd141351: dataIn1 = 32'd3021
; 
32'd141352: dataIn1 = 32'd3365
; 
32'd141353: dataIn1 = 32'd3369
; 
32'd141354: dataIn1 = 32'd4576
; 
32'd141355: dataIn1 = 32'd4585
; 
32'd141356: dataIn1 = 32'd1815
; 
32'd141357: dataIn1 = 32'd2024
; 
32'd141358: dataIn1 = 32'd2996
; 
32'd141359: dataIn1 = 32'd3370
; 
32'd141360: dataIn1 = 32'd3371
; 
32'd141361: dataIn1 = 32'd3372
; 
32'd141362: dataIn1 = 32'd3373
; 
32'd141363: dataIn1 = 32'd1819
; 
32'd141364: dataIn1 = 32'd2024
; 
32'd141365: dataIn1 = 32'd3006
; 
32'd141366: dataIn1 = 32'd3370
; 
32'd141367: dataIn1 = 32'd3371
; 
32'd141368: dataIn1 = 32'd3372
; 
32'd141369: dataIn1 = 32'd3374
; 
32'd141370: dataIn1 = 32'd1815
; 
32'd141371: dataIn1 = 32'd1819
; 
32'd141372: dataIn1 = 32'd3370
; 
32'd141373: dataIn1 = 32'd3371
; 
32'd141374: dataIn1 = 32'd3372
; 
32'd141375: dataIn1 = 32'd3375
; 
32'd141376: dataIn1 = 32'd3376
; 
32'd141377: dataIn1 = 32'd375
; 
32'd141378: dataIn1 = 32'd2024
; 
32'd141379: dataIn1 = 32'd2996
; 
32'd141380: dataIn1 = 32'd3370
; 
32'd141381: dataIn1 = 32'd3373
; 
32'd141382: dataIn1 = 32'd4566
; 
32'd141383: dataIn1 = 32'd4571
; 
32'd141384: dataIn1 = 32'd191
; 
32'd141385: dataIn1 = 32'd2024
; 
32'd141386: dataIn1 = 32'd3006
; 
32'd141387: dataIn1 = 32'd3371
; 
32'd141388: dataIn1 = 32'd3374
; 
32'd141389: dataIn1 = 32'd4559
; 
32'd141390: dataIn1 = 32'd4572
; 
32'd141391: dataIn1 = 32'd1815
; 
32'd141392: dataIn1 = 32'd2994
; 
32'd141393: dataIn1 = 32'd3372
; 
32'd141394: dataIn1 = 32'd3375
; 
32'd141395: dataIn1 = 32'd3376
; 
32'd141396: dataIn1 = 32'd11182
; 
32'd141397: dataIn1 = 32'd11183
; 
32'd141398: dataIn1 = 32'd1819
; 
32'd141399: dataIn1 = 32'd3004
; 
32'd141400: dataIn1 = 32'd3372
; 
32'd141401: dataIn1 = 32'd3375
; 
32'd141402: dataIn1 = 32'd3376
; 
32'd141403: dataIn1 = 32'd11181
; 
32'd141404: dataIn1 = 32'd11182
; 
32'd141405: dataIn1 = 32'd1818
; 
32'd141406: dataIn1 = 32'd1820
; 
32'd141407: dataIn1 = 32'd3377
; 
32'd141408: dataIn1 = 32'd3378
; 
32'd141409: dataIn1 = 32'd3379
; 
32'd141410: dataIn1 = 32'd3380
; 
32'd141411: dataIn1 = 32'd3381
; 
32'd141412: dataIn1 = 32'd1820
; 
32'd141413: dataIn1 = 32'd2025
; 
32'd141414: dataIn1 = 32'd3005
; 
32'd141415: dataIn1 = 32'd3377
; 
32'd141416: dataIn1 = 32'd3378
; 
32'd141417: dataIn1 = 32'd3379
; 
32'd141418: dataIn1 = 32'd3382
; 
32'd141419: dataIn1 = 32'd1818
; 
32'd141420: dataIn1 = 32'd2025
; 
32'd141421: dataIn1 = 32'd3000
; 
32'd141422: dataIn1 = 32'd3377
; 
32'd141423: dataIn1 = 32'd3378
; 
32'd141424: dataIn1 = 32'd3379
; 
32'd141425: dataIn1 = 32'd3383
; 
32'd141426: dataIn1 = 32'd1820
; 
32'd141427: dataIn1 = 32'd3002
; 
32'd141428: dataIn1 = 32'd3377
; 
32'd141429: dataIn1 = 32'd3380
; 
32'd141430: dataIn1 = 32'd3381
; 
32'd141431: dataIn1 = 32'd11177
; 
32'd141432: dataIn1 = 32'd11178
; 
32'd141433: dataIn1 = 32'd1818
; 
32'd141434: dataIn1 = 32'd2997
; 
32'd141435: dataIn1 = 32'd3377
; 
32'd141436: dataIn1 = 32'd3380
; 
32'd141437: dataIn1 = 32'd3381
; 
32'd141438: dataIn1 = 32'd11176
; 
32'd141439: dataIn1 = 32'd11177
; 
32'd141440: dataIn1 = 32'd191
; 
32'd141441: dataIn1 = 32'd2025
; 
32'd141442: dataIn1 = 32'd3005
; 
32'd141443: dataIn1 = 32'd3378
; 
32'd141444: dataIn1 = 32'd3382
; 
32'd141445: dataIn1 = 32'd4551
; 
32'd141446: dataIn1 = 32'd4558
; 
32'd141447: dataIn1 = 32'd381
; 
32'd141448: dataIn1 = 32'd2025
; 
32'd141449: dataIn1 = 32'd3000
; 
32'd141450: dataIn1 = 32'd3379
; 
32'd141451: dataIn1 = 32'd3383
; 
32'd141452: dataIn1 = 32'd4545
; 
32'd141453: dataIn1 = 32'd4552
; 
32'd141454: dataIn1 = 32'd1822
; 
32'd141455: dataIn1 = 32'd2026
; 
32'd141456: dataIn1 = 32'd3010
; 
32'd141457: dataIn1 = 32'd3384
; 
32'd141458: dataIn1 = 32'd3385
; 
32'd141459: dataIn1 = 32'd3386
; 
32'd141460: dataIn1 = 32'd3387
; 
32'd141461: dataIn1 = 32'd1817
; 
32'd141462: dataIn1 = 32'd1822
; 
32'd141463: dataIn1 = 32'd3384
; 
32'd141464: dataIn1 = 32'd3385
; 
32'd141465: dataIn1 = 32'd3386
; 
32'd141466: dataIn1 = 32'd3388
; 
32'd141467: dataIn1 = 32'd3389
; 
32'd141468: dataIn1 = 32'd1817
; 
32'd141469: dataIn1 = 32'd2026
; 
32'd141470: dataIn1 = 32'd3001
; 
32'd141471: dataIn1 = 32'd3384
; 
32'd141472: dataIn1 = 32'd3385
; 
32'd141473: dataIn1 = 32'd3386
; 
32'd141474: dataIn1 = 32'd3390
; 
32'd141475: dataIn1 = 32'd189
; 
32'd141476: dataIn1 = 32'd2026
; 
32'd141477: dataIn1 = 32'd3010
; 
32'd141478: dataIn1 = 32'd3384
; 
32'd141479: dataIn1 = 32'd3387
; 
32'd141480: dataIn1 = 32'd4537
; 
32'd141481: dataIn1 = 32'd4547
; 
32'd141482: dataIn1 = 32'd1822
; 
32'd141483: dataIn1 = 32'd3008
; 
32'd141484: dataIn1 = 32'd3385
; 
32'd141485: dataIn1 = 32'd3388
; 
32'd141486: dataIn1 = 32'd3389
; 
32'd141487: dataIn1 = 32'd11172
; 
32'd141488: dataIn1 = 32'd11173
; 
32'd141489: dataIn1 = 32'd1817
; 
32'd141490: dataIn1 = 32'd2998
; 
32'd141491: dataIn1 = 32'd3385
; 
32'd141492: dataIn1 = 32'd3388
; 
32'd141493: dataIn1 = 32'd3389
; 
32'd141494: dataIn1 = 32'd11173
; 
32'd141495: dataIn1 = 32'd11174
; 
32'd141496: dataIn1 = 32'd381
; 
32'd141497: dataIn1 = 32'd2026
; 
32'd141498: dataIn1 = 32'd3001
; 
32'd141499: dataIn1 = 32'd3386
; 
32'd141500: dataIn1 = 32'd3390
; 
32'd141501: dataIn1 = 32'd4546
; 
32'd141502: dataIn1 = 32'd4549
; 
32'd141503: dataIn1 = 32'd1824
; 
32'd141504: dataIn1 = 32'd1826
; 
32'd141505: dataIn1 = 32'd3391
; 
32'd141506: dataIn1 = 32'd3392
; 
32'd141507: dataIn1 = 32'd3393
; 
32'd141508: dataIn1 = 32'd3394
; 
32'd141509: dataIn1 = 32'd3395
; 
32'd141510: dataIn1 = 32'd1824
; 
32'd141511: dataIn1 = 32'd2027
; 
32'd141512: dataIn1 = 32'd3015
; 
32'd141513: dataIn1 = 32'd3391
; 
32'd141514: dataIn1 = 32'd3392
; 
32'd141515: dataIn1 = 32'd3393
; 
32'd141516: dataIn1 = 32'd3396
; 
32'd141517: dataIn1 = 32'd1826
; 
32'd141518: dataIn1 = 32'd2027
; 
32'd141519: dataIn1 = 32'd3020
; 
32'd141520: dataIn1 = 32'd3391
; 
32'd141521: dataIn1 = 32'd3392
; 
32'd141522: dataIn1 = 32'd3393
; 
32'd141523: dataIn1 = 32'd3397
; 
32'd141524: dataIn1 = 32'd1824
; 
32'd141525: dataIn1 = 32'd3012
; 
32'd141526: dataIn1 = 32'd3391
; 
32'd141527: dataIn1 = 32'd3394
; 
32'd141528: dataIn1 = 32'd3395
; 
32'd141529: dataIn1 = 32'd11190
; 
32'd141530: dataIn1 = 32'd11191
; 
32'd141531: dataIn1 = 32'd1826
; 
32'd141532: dataIn1 = 32'd3017
; 
32'd141533: dataIn1 = 32'd3391
; 
32'd141534: dataIn1 = 32'd3394
; 
32'd141535: dataIn1 = 32'd3395
; 
32'd141536: dataIn1 = 32'd11189
; 
32'd141537: dataIn1 = 32'd11190
; 
32'd141538: dataIn1 = 32'd382
; 
32'd141539: dataIn1 = 32'd2027
; 
32'd141540: dataIn1 = 32'd3015
; 
32'd141541: dataIn1 = 32'd3392
; 
32'd141542: dataIn1 = 32'd3396
; 
32'd141543: dataIn1 = 32'd4591
; 
32'd141544: dataIn1 = 32'd4600
; 
32'd141545: dataIn1 = 32'd192
; 
32'd141546: dataIn1 = 32'd2027
; 
32'd141547: dataIn1 = 32'd3020
; 
32'd141548: dataIn1 = 32'd3393
; 
32'd141549: dataIn1 = 32'd3397
; 
32'd141550: dataIn1 = 32'd4584
; 
32'd141551: dataIn1 = 32'd4601
; 
32'd141552: dataIn1 = 32'd1827
; 
32'd141553: dataIn1 = 32'd2028
; 
32'd141554: dataIn1 = 32'd3026
; 
32'd141555: dataIn1 = 32'd3398
; 
32'd141556: dataIn1 = 32'd3399
; 
32'd141557: dataIn1 = 32'd3400
; 
32'd141558: dataIn1 = 32'd3401
; 
32'd141559: dataIn1 = 32'd1823
; 
32'd141560: dataIn1 = 32'd2028
; 
32'd141561: dataIn1 = 32'd3016
; 
32'd141562: dataIn1 = 32'd3398
; 
32'd141563: dataIn1 = 32'd3399
; 
32'd141564: dataIn1 = 32'd3400
; 
32'd141565: dataIn1 = 32'd3402
; 
32'd141566: dataIn1 = 32'd1823
; 
32'd141567: dataIn1 = 32'd1827
; 
32'd141568: dataIn1 = 32'd3398
; 
32'd141569: dataIn1 = 32'd3399
; 
32'd141570: dataIn1 = 32'd3400
; 
32'd141571: dataIn1 = 32'd3403
; 
32'd141572: dataIn1 = 32'd3404
; 
32'd141573: dataIn1 = 32'd193
; 
32'd141574: dataIn1 = 32'd2028
; 
32'd141575: dataIn1 = 32'd3026
; 
32'd141576: dataIn1 = 32'd3398
; 
32'd141577: dataIn1 = 32'd3401
; 
32'd141578: dataIn1 = 32'd4595
; 
32'd141579: dataIn1 = 32'd5305
; 
32'd141580: dataIn1 = 32'd382
; 
32'd141581: dataIn1 = 32'd2028
; 
32'd141582: dataIn1 = 32'd3016
; 
32'd141583: dataIn1 = 32'd3399
; 
32'd141584: dataIn1 = 32'd3402
; 
32'd141585: dataIn1 = 32'd4592
; 
32'd141586: dataIn1 = 32'd4596
; 
32'd141587: dataIn1 = 32'd1827
; 
32'd141588: dataIn1 = 32'd3024
; 
32'd141589: dataIn1 = 32'd3400
; 
32'd141590: dataIn1 = 32'd3403
; 
32'd141591: dataIn1 = 32'd3404
; 
32'd141592: dataIn1 = 32'd11194
; 
32'd141593: dataIn1 = 32'd11195
; 
32'd141594: dataIn1 = 32'd1823
; 
32'd141595: dataIn1 = 32'd3014
; 
32'd141596: dataIn1 = 32'd3400
; 
32'd141597: dataIn1 = 32'd3403
; 
32'd141598: dataIn1 = 32'd3404
; 
32'd141599: dataIn1 = 32'd11193
; 
32'd141600: dataIn1 = 32'd11194
; 
32'd141601: dataIn1 = 32'd969
; 
32'd141602: dataIn1 = 32'd1847
; 
32'd141603: dataIn1 = 32'd2039
; 
32'd141604: dataIn1 = 32'd3405
; 
32'd141605: dataIn1 = 32'd3406
; 
32'd141606: dataIn1 = 32'd3407
; 
32'd141607: dataIn1 = 32'd1853
; 
32'd141608: dataIn1 = 32'd2039
; 
32'd141609: dataIn1 = 32'd3031
; 
32'd141610: dataIn1 = 32'd3405
; 
32'd141611: dataIn1 = 32'd3406
; 
32'd141612: dataIn1 = 32'd3407
; 
32'd141613: dataIn1 = 32'd3408
; 
32'd141614: dataIn1 = 32'd1847
; 
32'd141615: dataIn1 = 32'd1853
; 
32'd141616: dataIn1 = 32'd3405
; 
32'd141617: dataIn1 = 32'd3406
; 
32'd141618: dataIn1 = 32'd3407
; 
32'd141619: dataIn1 = 32'd3409
; 
32'd141620: dataIn1 = 32'd3410
; 
32'd141621: dataIn1 = 32'd391
; 
32'd141622: dataIn1 = 32'd2039
; 
32'd141623: dataIn1 = 32'd3031
; 
32'd141624: dataIn1 = 32'd3406
; 
32'd141625: dataIn1 = 32'd3408
; 
32'd141626: dataIn1 = 32'd4612
; 
32'd141627: dataIn1 = 32'd5306
; 
32'd141628: dataIn1 = 32'd203
; 
32'd141629: dataIn1 = 32'd1416
; 
32'd141630: dataIn1 = 32'd1847
; 
32'd141631: dataIn1 = 32'd3407
; 
32'd141632: dataIn1 = 32'd3409
; 
32'd141633: dataIn1 = 32'd3410
; 
32'd141634: dataIn1 = 32'd3446
; 
32'd141635: dataIn1 = 32'd203
; 
32'd141636: dataIn1 = 32'd1426
; 
32'd141637: dataIn1 = 32'd1853
; 
32'd141638: dataIn1 = 32'd3029
; 
32'd141639: dataIn1 = 32'd3407
; 
32'd141640: dataIn1 = 32'd3409
; 
32'd141641: dataIn1 = 32'd3410
; 
32'd141642: dataIn1 = 32'd758
; 
32'd141643: dataIn1 = 32'd1857
; 
32'd141644: dataIn1 = 32'd3411
; 
32'd141645: dataIn1 = 32'd3412
; 
32'd141646: dataIn1 = 32'd3413
; 
32'd141647: dataIn1 = 32'd10258
; 
32'd141648: dataIn1 = 32'd10270
; 
32'd141649: dataIn1 = 32'd394
; 
32'd141650: dataIn1 = 32'd758
; 
32'd141651: dataIn1 = 32'd1445
; 
32'd141652: dataIn1 = 32'd3411
; 
32'd141653: dataIn1 = 32'd3412
; 
32'd141654: dataIn1 = 32'd3413
; 
32'd141655: dataIn1 = 32'd3447
; 
32'd141656: dataIn1 = 32'd394
; 
32'd141657: dataIn1 = 32'd1439
; 
32'd141658: dataIn1 = 32'd1857
; 
32'd141659: dataIn1 = 32'd3032
; 
32'd141660: dataIn1 = 32'd3411
; 
32'd141661: dataIn1 = 32'd3412
; 
32'd141662: dataIn1 = 32'd3413
; 
32'd141663: dataIn1 = 32'd204
; 
32'd141664: dataIn1 = 32'd1440
; 
32'd141665: dataIn1 = 32'd1856
; 
32'd141666: dataIn1 = 32'd3033
; 
32'd141667: dataIn1 = 32'd3414
; 
32'd141668: dataIn1 = 32'd3415
; 
32'd141669: dataIn1 = 32'd3416
; 
32'd141670: dataIn1 = 32'd745
; 
32'd141671: dataIn1 = 32'd1856
; 
32'd141672: dataIn1 = 32'd2041
; 
32'd141673: dataIn1 = 32'd3414
; 
32'd141674: dataIn1 = 32'd3415
; 
32'd141675: dataIn1 = 32'd3416
; 
32'd141676: dataIn1 = 32'd204
; 
32'd141677: dataIn1 = 32'd745
; 
32'd141678: dataIn1 = 32'd1430
; 
32'd141679: dataIn1 = 32'd3414
; 
32'd141680: dataIn1 = 32'd3415
; 
32'd141681: dataIn1 = 32'd3416
; 
32'd141682: dataIn1 = 32'd3448
; 
32'd141683: dataIn1 = 32'd980
; 
32'd141684: dataIn1 = 32'd2048
; 
32'd141685: dataIn1 = 32'd3038
; 
32'd141686: dataIn1 = 32'd3417
; 
32'd141687: dataIn1 = 32'd3418
; 
32'd141688: dataIn1 = 32'd4625
; 
32'd141689: dataIn1 = 32'd5307
; 
32'd141690: dataIn1 = 32'd1869
; 
32'd141691: dataIn1 = 32'd2048
; 
32'd141692: dataIn1 = 32'd3038
; 
32'd141693: dataIn1 = 32'd3417
; 
32'd141694: dataIn1 = 32'd3418
; 
32'd141695: dataIn1 = 32'd10260
; 
32'd141696: dataIn1 = 32'd10261
; 
32'd141697: dataIn1 = 32'd17
; 
32'd141698: dataIn1 = 32'd27
; 
32'd141699: dataIn1 = 32'd1137
; 
32'd141700: dataIn1 = 32'd2138
; 
32'd141701: dataIn1 = 32'd2748
; 
32'd141702: dataIn1 = 32'd3419
; 
32'd141703: dataIn1 = 32'd3437
; 
32'd141704: dataIn1 = 32'd5515
; 
32'd141705: dataIn1 = 32'd156
; 
32'd141706: dataIn1 = 32'd442
; 
32'd141707: dataIn1 = 32'd586
; 
32'd141708: dataIn1 = 32'd2486
; 
32'd141709: dataIn1 = 32'd3420
; 
32'd141710: dataIn1 = 32'd3421
; 
32'd141711: dataIn1 = 32'd3454
; 
32'd141712: dataIn1 = 32'd3464
; 
32'd141713: dataIn1 = 32'd285
; 
32'd141714: dataIn1 = 32'd442
; 
32'd141715: dataIn1 = 32'd586
; 
32'd141716: dataIn1 = 32'd2295
; 
32'd141717: dataIn1 = 32'd2485
; 
32'd141718: dataIn1 = 32'd3420
; 
32'd141719: dataIn1 = 32'd3421
; 
32'd141720: dataIn1 = 32'd3449
; 
32'd141721: dataIn1 = 32'd5304
; 
32'd141722: dataIn1 = 32'd151
; 
32'd141723: dataIn1 = 32'd408
; 
32'd141724: dataIn1 = 32'd775
; 
32'd141725: dataIn1 = 32'd2495
; 
32'd141726: dataIn1 = 32'd3422
; 
32'd141727: dataIn1 = 32'd3423
; 
32'd141728: dataIn1 = 32'd3424
; 
32'd141729: dataIn1 = 32'd3451
; 
32'd141730: dataIn1 = 32'd151
; 
32'd141731: dataIn1 = 32'd407
; 
32'd141732: dataIn1 = 32'd775
; 
32'd141733: dataIn1 = 32'd976
; 
32'd141734: dataIn1 = 32'd2493
; 
32'd141735: dataIn1 = 32'd3422
; 
32'd141736: dataIn1 = 32'd3423
; 
32'd141737: dataIn1 = 32'd3450
; 
32'd141738: dataIn1 = 32'd271
; 
32'd141739: dataIn1 = 32'd408
; 
32'd141740: dataIn1 = 32'd784
; 
32'd141741: dataIn1 = 32'd2503
; 
32'd141742: dataIn1 = 32'd3422
; 
32'd141743: dataIn1 = 32'd3424
; 
32'd141744: dataIn1 = 32'd3425
; 
32'd141745: dataIn1 = 32'd3451
; 
32'd141746: dataIn1 = 32'd271
; 
32'd141747: dataIn1 = 32'd409
; 
32'd141748: dataIn1 = 32'd784
; 
32'd141749: dataIn1 = 32'd2502
; 
32'd141750: dataIn1 = 32'd3424
; 
32'd141751: dataIn1 = 32'd3425
; 
32'd141752: dataIn1 = 32'd3426
; 
32'd141753: dataIn1 = 32'd3452
; 
32'd141754: dataIn1 = 32'd2
; 
32'd141755: dataIn1 = 32'd409
; 
32'd141756: dataIn1 = 32'd786
; 
32'd141757: dataIn1 = 32'd2510
; 
32'd141758: dataIn1 = 32'd3425
; 
32'd141759: dataIn1 = 32'd3426
; 
32'd141760: dataIn1 = 32'd3427
; 
32'd141761: dataIn1 = 32'd3452
; 
32'd141762: dataIn1 = 32'd2
; 
32'd141763: dataIn1 = 32'd411
; 
32'd141764: dataIn1 = 32'd786
; 
32'd141765: dataIn1 = 32'd2508
; 
32'd141766: dataIn1 = 32'd3426
; 
32'd141767: dataIn1 = 32'd3427
; 
32'd141768: dataIn1 = 32'd3428
; 
32'd141769: dataIn1 = 32'd3453
; 
32'd141770: dataIn1 = 32'd411
; 
32'd141771: dataIn1 = 32'd416
; 
32'd141772: dataIn1 = 32'd805
; 
32'd141773: dataIn1 = 32'd2518
; 
32'd141774: dataIn1 = 32'd3427
; 
32'd141775: dataIn1 = 32'd3428
; 
32'd141776: dataIn1 = 32'd3429
; 
32'd141777: dataIn1 = 32'd3453
; 
32'd141778: dataIn1 = 32'd413
; 
32'd141779: dataIn1 = 32'd416
; 
32'd141780: dataIn1 = 32'd805
; 
32'd141781: dataIn1 = 32'd981
; 
32'd141782: dataIn1 = 32'd2517
; 
32'd141783: dataIn1 = 32'd3428
; 
32'd141784: dataIn1 = 32'd3429
; 
32'd141785: dataIn1 = 32'd3454
; 
32'd141786: dataIn1 = 32'd10264
; 
32'd141787: dataIn1 = 32'd202
; 
32'd141788: dataIn1 = 32'd1038
; 
32'd141789: dataIn1 = 32'd1072
; 
32'd141790: dataIn1 = 32'd2553
; 
32'd141791: dataIn1 = 32'd2556
; 
32'd141792: dataIn1 = 32'd3430
; 
32'd141793: dataIn1 = 32'd3455
; 
32'd141794: dataIn1 = 32'd132
; 
32'd141795: dataIn1 = 32'd1043
; 
32'd141796: dataIn1 = 32'd1077
; 
32'd141797: dataIn1 = 32'd2565
; 
32'd141798: dataIn1 = 32'd2634
; 
32'd141799: dataIn1 = 32'd3431
; 
32'd141800: dataIn1 = 32'd3432
; 
32'd141801: dataIn1 = 32'd4887
; 
32'd141802: dataIn1 = 32'd132
; 
32'd141803: dataIn1 = 32'd1044
; 
32'd141804: dataIn1 = 32'd1078
; 
32'd141805: dataIn1 = 32'd2634
; 
32'd141806: dataIn1 = 32'd3431
; 
32'd141807: dataIn1 = 32'd3432
; 
32'd141808: dataIn1 = 32'd3456
; 
32'd141809: dataIn1 = 32'd4889
; 
32'd141810: dataIn1 = 32'd15
; 
32'd141811: dataIn1 = 32'd25
; 
32'd141812: dataIn1 = 32'd1135
; 
32'd141813: dataIn1 = 32'd2130
; 
32'd141814: dataIn1 = 32'd2737
; 
32'd141815: dataIn1 = 32'd3433
; 
32'd141816: dataIn1 = 32'd3434
; 
32'd141817: dataIn1 = 32'd3436
; 
32'd141818: dataIn1 = 32'd14
; 
32'd141819: dataIn1 = 32'd25
; 
32'd141820: dataIn1 = 32'd1135
; 
32'd141821: dataIn1 = 32'd2126
; 
32'd141822: dataIn1 = 32'd3433
; 
32'd141823: dataIn1 = 32'd3434
; 
32'd141824: dataIn1 = 32'd3457
; 
32'd141825: dataIn1 = 32'd5513
; 
32'd141826: dataIn1 = 32'd16
; 
32'd141827: dataIn1 = 32'd26
; 
32'd141828: dataIn1 = 32'd1136
; 
32'd141829: dataIn1 = 32'd2134
; 
32'd141830: dataIn1 = 32'd2742
; 
32'd141831: dataIn1 = 32'd3435
; 
32'd141832: dataIn1 = 32'd3436
; 
32'd141833: dataIn1 = 32'd3437
; 
32'd141834: dataIn1 = 32'd15
; 
32'd141835: dataIn1 = 32'd26
; 
32'd141836: dataIn1 = 32'd1136
; 
32'd141837: dataIn1 = 32'd2130
; 
32'd141838: dataIn1 = 32'd2741
; 
32'd141839: dataIn1 = 32'd3433
; 
32'd141840: dataIn1 = 32'd3435
; 
32'd141841: dataIn1 = 32'd3436
; 
32'd141842: dataIn1 = 32'd16
; 
32'd141843: dataIn1 = 32'd27
; 
32'd141844: dataIn1 = 32'd1137
; 
32'd141845: dataIn1 = 32'd2134
; 
32'd141846: dataIn1 = 32'd2746
; 
32'd141847: dataIn1 = 32'd3419
; 
32'd141848: dataIn1 = 32'd3435
; 
32'd141849: dataIn1 = 32'd3437
; 
32'd141850: dataIn1 = 32'd264
; 
32'd141851: dataIn1 = 32'd543
; 
32'd141852: dataIn1 = 32'd1243
; 
32'd141853: dataIn1 = 32'd1253
; 
32'd141854: dataIn1 = 32'd2754
; 
32'd141855: dataIn1 = 32'd3438
; 
32'd141856: dataIn1 = 32'd3458
; 
32'd141857: dataIn1 = 32'd783
; 
32'd141858: dataIn1 = 32'd1462
; 
32'd141859: dataIn1 = 32'd1489
; 
32'd141860: dataIn1 = 32'd2758
; 
32'd141861: dataIn1 = 32'd3439
; 
32'd141862: dataIn1 = 32'd3459
; 
32'd141863: dataIn1 = 32'd11668
; 
32'd141864: dataIn1 = 32'd11669
; 
32'd141865: dataIn1 = 32'd414
; 
32'd141866: dataIn1 = 32'd806
; 
32'd141867: dataIn1 = 32'd1514
; 
32'd141868: dataIn1 = 32'd2760
; 
32'd141869: dataIn1 = 32'd3040
; 
32'd141870: dataIn1 = 32'd3440
; 
32'd141871: dataIn1 = 32'd3445
; 
32'd141872: dataIn1 = 32'd1828
; 
32'd141873: dataIn1 = 32'd3023
; 
32'd141874: dataIn1 = 32'd3441
; 
32'd141875: dataIn1 = 32'd11197
; 
32'd141876: dataIn1 = 32'd389
; 
32'd141877: dataIn1 = 32'd1425
; 
32'd141878: dataIn1 = 32'd1429
; 
32'd141879: dataIn1 = 32'd1854
; 
32'd141880: dataIn1 = 32'd3027
; 
32'd141881: dataIn1 = 32'd3442
; 
32'd141882: dataIn1 = 32'd3460
; 
32'd141883: dataIn1 = 32'd412
; 
32'd141884: dataIn1 = 32'd1502
; 
32'd141885: dataIn1 = 32'd1868
; 
32'd141886: dataIn1 = 32'd1871
; 
32'd141887: dataIn1 = 32'd3036
; 
32'd141888: dataIn1 = 32'd3443
; 
32'd141889: dataIn1 = 32'd211
; 
32'd141890: dataIn1 = 32'd1501
; 
32'd141891: dataIn1 = 32'd1869
; 
32'd141892: dataIn1 = 32'd3035
; 
32'd141893: dataIn1 = 32'd3444
; 
32'd141894: dataIn1 = 32'd10260
; 
32'd141895: dataIn1 = 32'd10262
; 
32'd141896: dataIn1 = 32'd800
; 
32'd141897: dataIn1 = 32'd806
; 
32'd141898: dataIn1 = 32'd3040
; 
32'd141899: dataIn1 = 32'd3440
; 
32'd141900: dataIn1 = 32'd3445
; 
32'd141901: dataIn1 = 32'd10251
; 
32'd141902: dataIn1 = 32'd10252
; 
32'd141903: dataIn1 = 32'd740
; 
32'd141904: dataIn1 = 32'd1416
; 
32'd141905: dataIn1 = 32'd1847
; 
32'd141906: dataIn1 = 32'd1848
; 
32'd141907: dataIn1 = 32'd3409
; 
32'd141908: dataIn1 = 32'd3446
; 
32'd141909: dataIn1 = 32'd757
; 
32'd141910: dataIn1 = 32'd758
; 
32'd141911: dataIn1 = 32'd1445
; 
32'd141912: dataIn1 = 32'd1447
; 
32'd141913: dataIn1 = 32'd3412
; 
32'd141914: dataIn1 = 32'd3447
; 
32'd141915: dataIn1 = 32'd3461
; 
32'd141916: dataIn1 = 32'd745
; 
32'd141917: dataIn1 = 32'd746
; 
32'd141918: dataIn1 = 32'd1424
; 
32'd141919: dataIn1 = 32'd1430
; 
32'd141920: dataIn1 = 32'd3416
; 
32'd141921: dataIn1 = 32'd3448
; 
32'd141922: dataIn1 = 32'd3462
; 
32'd141923: dataIn1 = 32'd442
; 
32'd141924: dataIn1 = 32'd443
; 
32'd141925: dataIn1 = 32'd2295
; 
32'd141926: dataIn1 = 32'd3421
; 
32'd141927: dataIn1 = 32'd3449
; 
32'd141928: dataIn1 = 32'd3499
; 
32'd141929: dataIn1 = 32'd3502
; 
32'd141930: dataIn1 = 32'd151
; 
32'd141931: dataIn1 = 32'd270
; 
32'd141932: dataIn1 = 32'd960
; 
32'd141933: dataIn1 = 32'd976
; 
32'd141934: dataIn1 = 32'd3423
; 
32'd141935: dataIn1 = 32'd3450
; 
32'd141936: dataIn1 = 32'd3463
; 
32'd141937: dataIn1 = 32'd151
; 
32'd141938: dataIn1 = 32'd271
; 
32'd141939: dataIn1 = 32'd3422
; 
32'd141940: dataIn1 = 32'd3424
; 
32'd141941: dataIn1 = 32'd3451
; 
32'd141942: dataIn1 = 32'd3471
; 
32'd141943: dataIn1 = 32'd3475
; 
32'd141944: dataIn1 = 32'd2
; 
32'd141945: dataIn1 = 32'd271
; 
32'd141946: dataIn1 = 32'd3425
; 
32'd141947: dataIn1 = 32'd3426
; 
32'd141948: dataIn1 = 32'd3452
; 
32'd141949: dataIn1 = 32'd3479
; 
32'd141950: dataIn1 = 32'd3483
; 
32'd141951: dataIn1 = 32'd2
; 
32'd141952: dataIn1 = 32'd416
; 
32'd141953: dataIn1 = 32'd3427
; 
32'd141954: dataIn1 = 32'd3428
; 
32'd141955: dataIn1 = 32'd3453
; 
32'd141956: dataIn1 = 32'd3487
; 
32'd141957: dataIn1 = 32'd3491
; 
32'd141958: dataIn1 = 32'd156
; 
32'd141959: dataIn1 = 32'd416
; 
32'd141960: dataIn1 = 32'd981
; 
32'd141961: dataIn1 = 32'd3420
; 
32'd141962: dataIn1 = 32'd3429
; 
32'd141963: dataIn1 = 32'd3454
; 
32'd141964: dataIn1 = 32'd3464
; 
32'd141965: dataIn1 = 32'd10265
; 
32'd141966: dataIn1 = 32'd125
; 
32'd141967: dataIn1 = 32'd1038
; 
32'd141968: dataIn1 = 32'd1072
; 
32'd141969: dataIn1 = 32'd2613
; 
32'd141970: dataIn1 = 32'd3430
; 
32'd141971: dataIn1 = 32'd3455
; 
32'd141972: dataIn1 = 32'd3465
; 
32'd141973: dataIn1 = 32'd215
; 
32'd141974: dataIn1 = 32'd1044
; 
32'd141975: dataIn1 = 32'd1078
; 
32'd141976: dataIn1 = 32'd2571
; 
32'd141977: dataIn1 = 32'd3432
; 
32'd141978: dataIn1 = 32'd3456
; 
32'd141979: dataIn1 = 32'd3466
; 
32'd141980: dataIn1 = 32'd4690
; 
32'd141981: dataIn1 = 32'd14
; 
32'd141982: dataIn1 = 32'd24
; 
32'd141983: dataIn1 = 32'd2102
; 
32'd141984: dataIn1 = 32'd2126
; 
32'd141985: dataIn1 = 32'd3434
; 
32'd141986: dataIn1 = 32'd3457
; 
32'd141987: dataIn1 = 32'd3467
; 
32'd141988: dataIn1 = 32'd6730
; 
32'd141989: dataIn1 = 32'd9314
; 
32'd141990: dataIn1 = 32'd264
; 
32'd141991: dataIn1 = 32'd545
; 
32'd141992: dataIn1 = 32'd1253
; 
32'd141993: dataIn1 = 32'd1256
; 
32'd141994: dataIn1 = 32'd3438
; 
32'd141995: dataIn1 = 32'd3458
; 
32'd141996: dataIn1 = 32'd3468
; 
32'd141997: dataIn1 = 32'd782
; 
32'd141998: dataIn1 = 32'd783
; 
32'd141999: dataIn1 = 32'd976
; 
32'd142000: dataIn1 = 32'd1489
; 
32'd142001: dataIn1 = 32'd3439
; 
32'd142002: dataIn1 = 32'd3459
; 
32'd142003: dataIn1 = 32'd749
; 
32'd142004: dataIn1 = 32'd1429
; 
32'd142005: dataIn1 = 32'd1854
; 
32'd142006: dataIn1 = 32'd3442
; 
32'd142007: dataIn1 = 32'd3460
; 
32'd142008: dataIn1 = 32'd10256
; 
32'd142009: dataIn1 = 32'd10271
; 
32'd142010: dataIn1 = 32'd758
; 
32'd142011: dataIn1 = 32'd1447
; 
32'd142012: dataIn1 = 32'd1471
; 
32'd142013: dataIn1 = 32'd3447
; 
32'd142014: dataIn1 = 32'd3461
; 
32'd142015: dataIn1 = 32'd3469
; 
32'd142016: dataIn1 = 32'd10673
; 
32'd142017: dataIn1 = 32'd743
; 
32'd142018: dataIn1 = 32'd745
; 
32'd142019: dataIn1 = 32'd1421
; 
32'd142020: dataIn1 = 32'd1424
; 
32'd142021: dataIn1 = 32'd3448
; 
32'd142022: dataIn1 = 32'd3462
; 
32'd142023: dataIn1 = 32'd3470
; 
32'd142024: dataIn1 = 32'd151
; 
32'd142025: dataIn1 = 32'd268
; 
32'd142026: dataIn1 = 32'd552
; 
32'd142027: dataIn1 = 32'd960
; 
32'd142028: dataIn1 = 32'd3450
; 
32'd142029: dataIn1 = 32'd3463
; 
32'd142030: dataIn1 = 32'd3471
; 
32'd142031: dataIn1 = 32'd416
; 
32'd142032: dataIn1 = 32'd442
; 
32'd142033: dataIn1 = 32'd3420
; 
32'd142034: dataIn1 = 32'd3454
; 
32'd142035: dataIn1 = 32'd3464
; 
32'd142036: dataIn1 = 32'd3491
; 
32'd142037: dataIn1 = 32'd3495
; 
32'd142038: dataIn1 = 32'd125
; 
32'd142039: dataIn1 = 32'd1037
; 
32'd142040: dataIn1 = 32'd1071
; 
32'd142041: dataIn1 = 32'd2613
; 
32'd142042: dataIn1 = 32'd3455
; 
32'd142043: dataIn1 = 32'd3465
; 
32'd142044: dataIn1 = 32'd3472
; 
32'd142045: dataIn1 = 32'd215
; 
32'd142046: dataIn1 = 32'd1045
; 
32'd142047: dataIn1 = 32'd1079
; 
32'd142048: dataIn1 = 32'd2571
; 
32'd142049: dataIn1 = 32'd3456
; 
32'd142050: dataIn1 = 32'd3466
; 
32'd142051: dataIn1 = 32'd3473
; 
32'd142052: dataIn1 = 32'd4692
; 
32'd142053: dataIn1 = 32'd13
; 
32'd142054: dataIn1 = 32'd24
; 
32'd142055: dataIn1 = 32'd3457
; 
32'd142056: dataIn1 = 32'd3467
; 
32'd142057: dataIn1 = 32'd9314
; 
32'd142058: dataIn1 = 32'd545
; 
32'd142059: dataIn1 = 32'd546
; 
32'd142060: dataIn1 = 32'd1251
; 
32'd142061: dataIn1 = 32'd1256
; 
32'd142062: dataIn1 = 32'd3458
; 
32'd142063: dataIn1 = 32'd3468
; 
32'd142064: dataIn1 = 32'd3474
; 
32'd142065: dataIn1 = 32'd397
; 
32'd142066: dataIn1 = 32'd758
; 
32'd142067: dataIn1 = 32'd1471
; 
32'd142068: dataIn1 = 32'd3461
; 
32'd142069: dataIn1 = 32'd3469
; 
32'd142070: dataIn1 = 32'd10258
; 
32'd142071: dataIn1 = 32'd10259
; 
32'd142072: dataIn1 = 32'd390
; 
32'd142073: dataIn1 = 32'd745
; 
32'd142074: dataIn1 = 32'd1421
; 
32'd142075: dataIn1 = 32'd2041
; 
32'd142076: dataIn1 = 32'd3462
; 
32'd142077: dataIn1 = 32'd3470
; 
32'd142078: dataIn1 = 32'd151
; 
32'd142079: dataIn1 = 32'd269
; 
32'd142080: dataIn1 = 32'd552
; 
32'd142081: dataIn1 = 32'd3451
; 
32'd142082: dataIn1 = 32'd3463
; 
32'd142083: dataIn1 = 32'd3471
; 
32'd142084: dataIn1 = 32'd3475
; 
32'd142085: dataIn1 = 32'd199
; 
32'd142086: dataIn1 = 32'd1037
; 
32'd142087: dataIn1 = 32'd1071
; 
32'd142088: dataIn1 = 32'd2550
; 
32'd142089: dataIn1 = 32'd3465
; 
32'd142090: dataIn1 = 32'd3472
; 
32'd142091: dataIn1 = 32'd3476
; 
32'd142092: dataIn1 = 32'd134
; 
32'd142093: dataIn1 = 32'd1045
; 
32'd142094: dataIn1 = 32'd1079
; 
32'd142095: dataIn1 = 32'd2638
; 
32'd142096: dataIn1 = 32'd3466
; 
32'd142097: dataIn1 = 32'd3473
; 
32'd142098: dataIn1 = 32'd3477
; 
32'd142099: dataIn1 = 32'd4910
; 
32'd142100: dataIn1 = 32'd544
; 
32'd142101: dataIn1 = 32'd546
; 
32'd142102: dataIn1 = 32'd1251
; 
32'd142103: dataIn1 = 32'd1257
; 
32'd142104: dataIn1 = 32'd3468
; 
32'd142105: dataIn1 = 32'd3474
; 
32'd142106: dataIn1 = 32'd3478
; 
32'd142107: dataIn1 = 32'd269
; 
32'd142108: dataIn1 = 32'd271
; 
32'd142109: dataIn1 = 32'd559
; 
32'd142110: dataIn1 = 32'd3451
; 
32'd142111: dataIn1 = 32'd3471
; 
32'd142112: dataIn1 = 32'd3475
; 
32'd142113: dataIn1 = 32'd3479
; 
32'd142114: dataIn1 = 32'd199
; 
32'd142115: dataIn1 = 32'd1036
; 
32'd142116: dataIn1 = 32'd1070
; 
32'd142117: dataIn1 = 32'd2550
; 
32'd142118: dataIn1 = 32'd3472
; 
32'd142119: dataIn1 = 32'd3476
; 
32'd142120: dataIn1 = 32'd3480
; 
32'd142121: dataIn1 = 32'd134
; 
32'd142122: dataIn1 = 32'd1046
; 
32'd142123: dataIn1 = 32'd1080
; 
32'd142124: dataIn1 = 32'd2638
; 
32'd142125: dataIn1 = 32'd3473
; 
32'd142126: dataIn1 = 32'd3477
; 
32'd142127: dataIn1 = 32'd3481
; 
32'd142128: dataIn1 = 32'd4907
; 
32'd142129: dataIn1 = 32'd260
; 
32'd142130: dataIn1 = 32'd544
; 
32'd142131: dataIn1 = 32'd1252
; 
32'd142132: dataIn1 = 32'd1257
; 
32'd142133: dataIn1 = 32'd3474
; 
32'd142134: dataIn1 = 32'd3478
; 
32'd142135: dataIn1 = 32'd3482
; 
32'd142136: dataIn1 = 32'd271
; 
32'd142137: dataIn1 = 32'd272
; 
32'd142138: dataIn1 = 32'd559
; 
32'd142139: dataIn1 = 32'd3452
; 
32'd142140: dataIn1 = 32'd3475
; 
32'd142141: dataIn1 = 32'd3479
; 
32'd142142: dataIn1 = 32'd3483
; 
32'd142143: dataIn1 = 32'd122
; 
32'd142144: dataIn1 = 32'd1036
; 
32'd142145: dataIn1 = 32'd1070
; 
32'd142146: dataIn1 = 32'd2609
; 
32'd142147: dataIn1 = 32'd3476
; 
32'd142148: dataIn1 = 32'd3480
; 
32'd142149: dataIn1 = 32'd3484
; 
32'd142150: dataIn1 = 32'd218
; 
32'd142151: dataIn1 = 32'd1046
; 
32'd142152: dataIn1 = 32'd1080
; 
32'd142153: dataIn1 = 32'd2575
; 
32'd142154: dataIn1 = 32'd3477
; 
32'd142155: dataIn1 = 32'd3481
; 
32'd142156: dataIn1 = 32'd3485
; 
32'd142157: dataIn1 = 32'd4697
; 
32'd142158: dataIn1 = 32'd260
; 
32'd142159: dataIn1 = 32'd531
; 
32'd142160: dataIn1 = 32'd1211
; 
32'd142161: dataIn1 = 32'd1252
; 
32'd142162: dataIn1 = 32'd3478
; 
32'd142163: dataIn1 = 32'd3482
; 
32'd142164: dataIn1 = 32'd3486
; 
32'd142165: dataIn1 = 32'd2
; 
32'd142166: dataIn1 = 32'd272
; 
32'd142167: dataIn1 = 32'd569
; 
32'd142168: dataIn1 = 32'd3452
; 
32'd142169: dataIn1 = 32'd3479
; 
32'd142170: dataIn1 = 32'd3483
; 
32'd142171: dataIn1 = 32'd3487
; 
32'd142172: dataIn1 = 32'd122
; 
32'd142173: dataIn1 = 32'd1035
; 
32'd142174: dataIn1 = 32'd1069
; 
32'd142175: dataIn1 = 32'd2609
; 
32'd142176: dataIn1 = 32'd3480
; 
32'd142177: dataIn1 = 32'd3484
; 
32'd142178: dataIn1 = 32'd3488
; 
32'd142179: dataIn1 = 32'd218
; 
32'd142180: dataIn1 = 32'd1047
; 
32'd142181: dataIn1 = 32'd1081
; 
32'd142182: dataIn1 = 32'd2575
; 
32'd142183: dataIn1 = 32'd3481
; 
32'd142184: dataIn1 = 32'd3485
; 
32'd142185: dataIn1 = 32'd3489
; 
32'd142186: dataIn1 = 32'd4700
; 
32'd142187: dataIn1 = 32'd529
; 
32'd142188: dataIn1 = 32'd531
; 
32'd142189: dataIn1 = 32'd1211
; 
32'd142190: dataIn1 = 32'd1214
; 
32'd142191: dataIn1 = 32'd3482
; 
32'd142192: dataIn1 = 32'd3486
; 
32'd142193: dataIn1 = 32'd3490
; 
32'd142194: dataIn1 = 32'd2
; 
32'd142195: dataIn1 = 32'd277
; 
32'd142196: dataIn1 = 32'd569
; 
32'd142197: dataIn1 = 32'd3453
; 
32'd142198: dataIn1 = 32'd3483
; 
32'd142199: dataIn1 = 32'd3487
; 
32'd142200: dataIn1 = 32'd3491
; 
32'd142201: dataIn1 = 32'd195
; 
32'd142202: dataIn1 = 32'd1035
; 
32'd142203: dataIn1 = 32'd1069
; 
32'd142204: dataIn1 = 32'd2548
; 
32'd142205: dataIn1 = 32'd3484
; 
32'd142206: dataIn1 = 32'd3488
; 
32'd142207: dataIn1 = 32'd3492
; 
32'd142208: dataIn1 = 32'd135
; 
32'd142209: dataIn1 = 32'd1047
; 
32'd142210: dataIn1 = 32'd1081
; 
32'd142211: dataIn1 = 32'd2644
; 
32'd142212: dataIn1 = 32'd3485
; 
32'd142213: dataIn1 = 32'd3489
; 
32'd142214: dataIn1 = 32'd3493
; 
32'd142215: dataIn1 = 32'd4925
; 
32'd142216: dataIn1 = 32'd529
; 
32'd142217: dataIn1 = 32'd530
; 
32'd142218: dataIn1 = 32'd1213
; 
32'd142219: dataIn1 = 32'd1214
; 
32'd142220: dataIn1 = 32'd3486
; 
32'd142221: dataIn1 = 32'd3490
; 
32'd142222: dataIn1 = 32'd3494
; 
32'd142223: dataIn1 = 32'd277
; 
32'd142224: dataIn1 = 32'd416
; 
32'd142225: dataIn1 = 32'd3453
; 
32'd142226: dataIn1 = 32'd3464
; 
32'd142227: dataIn1 = 32'd3487
; 
32'd142228: dataIn1 = 32'd3491
; 
32'd142229: dataIn1 = 32'd3495
; 
32'd142230: dataIn1 = 32'd195
; 
32'd142231: dataIn1 = 32'd1034
; 
32'd142232: dataIn1 = 32'd1068
; 
32'd142233: dataIn1 = 32'd2548
; 
32'd142234: dataIn1 = 32'd3488
; 
32'd142235: dataIn1 = 32'd3492
; 
32'd142236: dataIn1 = 32'd3496
; 
32'd142237: dataIn1 = 32'd135
; 
32'd142238: dataIn1 = 32'd1048
; 
32'd142239: dataIn1 = 32'd1082
; 
32'd142240: dataIn1 = 32'd2644
; 
32'd142241: dataIn1 = 32'd3489
; 
32'd142242: dataIn1 = 32'd3493
; 
32'd142243: dataIn1 = 32'd3497
; 
32'd142244: dataIn1 = 32'd4927
; 
32'd142245: dataIn1 = 32'd261
; 
32'd142246: dataIn1 = 32'd530
; 
32'd142247: dataIn1 = 32'd1213
; 
32'd142248: dataIn1 = 32'd1227
; 
32'd142249: dataIn1 = 32'd3490
; 
32'd142250: dataIn1 = 32'd3494
; 
32'd142251: dataIn1 = 32'd3498
; 
32'd142252: dataIn1 = 32'd277
; 
32'd142253: dataIn1 = 32'd442
; 
32'd142254: dataIn1 = 32'd571
; 
32'd142255: dataIn1 = 32'd3464
; 
32'd142256: dataIn1 = 32'd3491
; 
32'd142257: dataIn1 = 32'd3495
; 
32'd142258: dataIn1 = 32'd3499
; 
32'd142259: dataIn1 = 32'd123
; 
32'd142260: dataIn1 = 32'd1034
; 
32'd142261: dataIn1 = 32'd1068
; 
32'd142262: dataIn1 = 32'd3492
; 
32'd142263: dataIn1 = 32'd3496
; 
32'd142264: dataIn1 = 32'd221
; 
32'd142265: dataIn1 = 32'd1048
; 
32'd142266: dataIn1 = 32'd1082
; 
32'd142267: dataIn1 = 32'd2577
; 
32'd142268: dataIn1 = 32'd3493
; 
32'd142269: dataIn1 = 32'd3497
; 
32'd142270: dataIn1 = 32'd3500
; 
32'd142271: dataIn1 = 32'd4708
; 
32'd142272: dataIn1 = 32'd261
; 
32'd142273: dataIn1 = 32'd535
; 
32'd142274: dataIn1 = 32'd1227
; 
32'd142275: dataIn1 = 32'd1231
; 
32'd142276: dataIn1 = 32'd3494
; 
32'd142277: dataIn1 = 32'd3498
; 
32'd142278: dataIn1 = 32'd3501
; 
32'd142279: dataIn1 = 32'd152
; 
32'd142280: dataIn1 = 32'd442
; 
32'd142281: dataIn1 = 32'd571
; 
32'd142282: dataIn1 = 32'd3449
; 
32'd142283: dataIn1 = 32'd3495
; 
32'd142284: dataIn1 = 32'd3499
; 
32'd142285: dataIn1 = 32'd3502
; 
32'd142286: dataIn1 = 32'd221
; 
32'd142287: dataIn1 = 32'd1049
; 
32'd142288: dataIn1 = 32'd1083
; 
32'd142289: dataIn1 = 32'd2577
; 
32'd142290: dataIn1 = 32'd3497
; 
32'd142291: dataIn1 = 32'd3500
; 
32'd142292: dataIn1 = 32'd3503
; 
32'd142293: dataIn1 = 32'd4710
; 
32'd142294: dataIn1 = 32'd535
; 
32'd142295: dataIn1 = 32'd536
; 
32'd142296: dataIn1 = 32'd1226
; 
32'd142297: dataIn1 = 32'd1231
; 
32'd142298: dataIn1 = 32'd3498
; 
32'd142299: dataIn1 = 32'd3501
; 
32'd142300: dataIn1 = 32'd3504
; 
32'd142301: dataIn1 = 32'd152
; 
32'd142302: dataIn1 = 32'd443
; 
32'd142303: dataIn1 = 32'd3449
; 
32'd142304: dataIn1 = 32'd3499
; 
32'd142305: dataIn1 = 32'd3502
; 
32'd142306: dataIn1 = 32'd5319
; 
32'd142307: dataIn1 = 32'd5457
; 
32'd142308: dataIn1 = 32'd137
; 
32'd142309: dataIn1 = 32'd1049
; 
32'd142310: dataIn1 = 32'd1083
; 
32'd142311: dataIn1 = 32'd2648
; 
32'd142312: dataIn1 = 32'd3500
; 
32'd142313: dataIn1 = 32'd3503
; 
32'd142314: dataIn1 = 32'd3505
; 
32'd142315: dataIn1 = 32'd4948
; 
32'd142316: dataIn1 = 32'd536
; 
32'd142317: dataIn1 = 32'd537
; 
32'd142318: dataIn1 = 32'd1226
; 
32'd142319: dataIn1 = 32'd1230
; 
32'd142320: dataIn1 = 32'd3501
; 
32'd142321: dataIn1 = 32'd3504
; 
32'd142322: dataIn1 = 32'd3506
; 
32'd142323: dataIn1 = 32'd137
; 
32'd142324: dataIn1 = 32'd1050
; 
32'd142325: dataIn1 = 32'd1084
; 
32'd142326: dataIn1 = 32'd2648
; 
32'd142327: dataIn1 = 32'd3503
; 
32'd142328: dataIn1 = 32'd3505
; 
32'd142329: dataIn1 = 32'd3507
; 
32'd142330: dataIn1 = 32'd4945
; 
32'd142331: dataIn1 = 32'd262
; 
32'd142332: dataIn1 = 32'd537
; 
32'd142333: dataIn1 = 32'd1230
; 
32'd142334: dataIn1 = 32'd1232
; 
32'd142335: dataIn1 = 32'd3504
; 
32'd142336: dataIn1 = 32'd3506
; 
32'd142337: dataIn1 = 32'd3508
; 
32'd142338: dataIn1 = 32'd224
; 
32'd142339: dataIn1 = 32'd1050
; 
32'd142340: dataIn1 = 32'd1084
; 
32'd142341: dataIn1 = 32'd2581
; 
32'd142342: dataIn1 = 32'd3505
; 
32'd142343: dataIn1 = 32'd3507
; 
32'd142344: dataIn1 = 32'd3509
; 
32'd142345: dataIn1 = 32'd4715
; 
32'd142346: dataIn1 = 32'd262
; 
32'd142347: dataIn1 = 32'd534
; 
32'd142348: dataIn1 = 32'd1219
; 
32'd142349: dataIn1 = 32'd1232
; 
32'd142350: dataIn1 = 32'd3506
; 
32'd142351: dataIn1 = 32'd3508
; 
32'd142352: dataIn1 = 32'd3510
; 
32'd142353: dataIn1 = 32'd224
; 
32'd142354: dataIn1 = 32'd1051
; 
32'd142355: dataIn1 = 32'd1085
; 
32'd142356: dataIn1 = 32'd2581
; 
32'd142357: dataIn1 = 32'd3507
; 
32'd142358: dataIn1 = 32'd3509
; 
32'd142359: dataIn1 = 32'd3511
; 
32'd142360: dataIn1 = 32'd4718
; 
32'd142361: dataIn1 = 32'd532
; 
32'd142362: dataIn1 = 32'd534
; 
32'd142363: dataIn1 = 32'd1219
; 
32'd142364: dataIn1 = 32'd1225
; 
32'd142365: dataIn1 = 32'd3508
; 
32'd142366: dataIn1 = 32'd3510
; 
32'd142367: dataIn1 = 32'd3512
; 
32'd142368: dataIn1 = 32'd138
; 
32'd142369: dataIn1 = 32'd1051
; 
32'd142370: dataIn1 = 32'd1085
; 
32'd142371: dataIn1 = 32'd2654
; 
32'd142372: dataIn1 = 32'd3509
; 
32'd142373: dataIn1 = 32'd3511
; 
32'd142374: dataIn1 = 32'd3513
; 
32'd142375: dataIn1 = 32'd4963
; 
32'd142376: dataIn1 = 32'd532
; 
32'd142377: dataIn1 = 32'd533
; 
32'd142378: dataIn1 = 32'd1221
; 
32'd142379: dataIn1 = 32'd1225
; 
32'd142380: dataIn1 = 32'd3510
; 
32'd142381: dataIn1 = 32'd3512
; 
32'd142382: dataIn1 = 32'd3514
; 
32'd142383: dataIn1 = 32'd138
; 
32'd142384: dataIn1 = 32'd1052
; 
32'd142385: dataIn1 = 32'd1086
; 
32'd142386: dataIn1 = 32'd2654
; 
32'd142387: dataIn1 = 32'd3511
; 
32'd142388: dataIn1 = 32'd3513
; 
32'd142389: dataIn1 = 32'd3515
; 
32'd142390: dataIn1 = 32'd4965
; 
32'd142391: dataIn1 = 32'd263
; 
32'd142392: dataIn1 = 32'd533
; 
32'd142393: dataIn1 = 32'd1221
; 
32'd142394: dataIn1 = 32'd1239
; 
32'd142395: dataIn1 = 32'd3512
; 
32'd142396: dataIn1 = 32'd3514
; 
32'd142397: dataIn1 = 32'd3516
; 
32'd142398: dataIn1 = 32'd227
; 
32'd142399: dataIn1 = 32'd1052
; 
32'd142400: dataIn1 = 32'd1086
; 
32'd142401: dataIn1 = 32'd2583
; 
32'd142402: dataIn1 = 32'd3513
; 
32'd142403: dataIn1 = 32'd3515
; 
32'd142404: dataIn1 = 32'd3517
; 
32'd142405: dataIn1 = 32'd4726
; 
32'd142406: dataIn1 = 32'd263
; 
32'd142407: dataIn1 = 32'd540
; 
32'd142408: dataIn1 = 32'd1236
; 
32'd142409: dataIn1 = 32'd1239
; 
32'd142410: dataIn1 = 32'd3514
; 
32'd142411: dataIn1 = 32'd3516
; 
32'd142412: dataIn1 = 32'd3518
; 
32'd142413: dataIn1 = 32'd227
; 
32'd142414: dataIn1 = 32'd1053
; 
32'd142415: dataIn1 = 32'd1087
; 
32'd142416: dataIn1 = 32'd2583
; 
32'd142417: dataIn1 = 32'd3515
; 
32'd142418: dataIn1 = 32'd3517
; 
32'd142419: dataIn1 = 32'd3519
; 
32'd142420: dataIn1 = 32'd4728
; 
32'd142421: dataIn1 = 32'd538
; 
32'd142422: dataIn1 = 32'd540
; 
32'd142423: dataIn1 = 32'd1233
; 
32'd142424: dataIn1 = 32'd1236
; 
32'd142425: dataIn1 = 32'd3516
; 
32'd142426: dataIn1 = 32'd3518
; 
32'd142427: dataIn1 = 32'd3520
; 
32'd142428: dataIn1 = 32'd140
; 
32'd142429: dataIn1 = 32'd1053
; 
32'd142430: dataIn1 = 32'd1087
; 
32'd142431: dataIn1 = 32'd2658
; 
32'd142432: dataIn1 = 32'd3517
; 
32'd142433: dataIn1 = 32'd3519
; 
32'd142434: dataIn1 = 32'd3521
; 
32'd142435: dataIn1 = 32'd4986
; 
32'd142436: dataIn1 = 32'd538
; 
32'd142437: dataIn1 = 32'd539
; 
32'd142438: dataIn1 = 32'd1233
; 
32'd142439: dataIn1 = 32'd1237
; 
32'd142440: dataIn1 = 32'd3518
; 
32'd142441: dataIn1 = 32'd3520
; 
32'd142442: dataIn1 = 32'd3522
; 
32'd142443: dataIn1 = 32'd140
; 
32'd142444: dataIn1 = 32'd1054
; 
32'd142445: dataIn1 = 32'd1088
; 
32'd142446: dataIn1 = 32'd2658
; 
32'd142447: dataIn1 = 32'd3519
; 
32'd142448: dataIn1 = 32'd3521
; 
32'd142449: dataIn1 = 32'd3523
; 
32'd142450: dataIn1 = 32'd4983
; 
32'd142451: dataIn1 = 32'd259
; 
32'd142452: dataIn1 = 32'd539
; 
32'd142453: dataIn1 = 32'd1237
; 
32'd142454: dataIn1 = 32'd1238
; 
32'd142455: dataIn1 = 32'd3520
; 
32'd142456: dataIn1 = 32'd3522
; 
32'd142457: dataIn1 = 32'd3524
; 
32'd142458: dataIn1 = 32'd230
; 
32'd142459: dataIn1 = 32'd1054
; 
32'd142460: dataIn1 = 32'd1088
; 
32'd142461: dataIn1 = 32'd2587
; 
32'd142462: dataIn1 = 32'd3521
; 
32'd142463: dataIn1 = 32'd3523
; 
32'd142464: dataIn1 = 32'd3525
; 
32'd142465: dataIn1 = 32'd4733
; 
32'd142466: dataIn1 = 32'd259
; 
32'd142467: dataIn1 = 32'd528
; 
32'd142468: dataIn1 = 32'd1203
; 
32'd142469: dataIn1 = 32'd1238
; 
32'd142470: dataIn1 = 32'd3522
; 
32'd142471: dataIn1 = 32'd3524
; 
32'd142472: dataIn1 = 32'd3526
; 
32'd142473: dataIn1 = 32'd230
; 
32'd142474: dataIn1 = 32'd1055
; 
32'd142475: dataIn1 = 32'd1089
; 
32'd142476: dataIn1 = 32'd2587
; 
32'd142477: dataIn1 = 32'd3523
; 
32'd142478: dataIn1 = 32'd3525
; 
32'd142479: dataIn1 = 32'd3527
; 
32'd142480: dataIn1 = 32'd4736
; 
32'd142481: dataIn1 = 32'd527
; 
32'd142482: dataIn1 = 32'd528
; 
32'd142483: dataIn1 = 32'd1203
; 
32'd142484: dataIn1 = 32'd1206
; 
32'd142485: dataIn1 = 32'd3524
; 
32'd142486: dataIn1 = 32'd3526
; 
32'd142487: dataIn1 = 32'd3528
; 
32'd142488: dataIn1 = 32'd141
; 
32'd142489: dataIn1 = 32'd1055
; 
32'd142490: dataIn1 = 32'd1089
; 
32'd142491: dataIn1 = 32'd2664
; 
32'd142492: dataIn1 = 32'd3525
; 
32'd142493: dataIn1 = 32'd3527
; 
32'd142494: dataIn1 = 32'd3529
; 
32'd142495: dataIn1 = 32'd5001
; 
32'd142496: dataIn1 = 32'd526
; 
32'd142497: dataIn1 = 32'd527
; 
32'd142498: dataIn1 = 32'd1204
; 
32'd142499: dataIn1 = 32'd1206
; 
32'd142500: dataIn1 = 32'd3526
; 
32'd142501: dataIn1 = 32'd3528
; 
32'd142502: dataIn1 = 32'd3530
; 
32'd142503: dataIn1 = 32'd141
; 
32'd142504: dataIn1 = 32'd1056
; 
32'd142505: dataIn1 = 32'd1090
; 
32'd142506: dataIn1 = 32'd2664
; 
32'd142507: dataIn1 = 32'd3527
; 
32'd142508: dataIn1 = 32'd3529
; 
32'd142509: dataIn1 = 32'd3531
; 
32'd142510: dataIn1 = 32'd5003
; 
32'd142511: dataIn1 = 32'd258
; 
32'd142512: dataIn1 = 32'd526
; 
32'd142513: dataIn1 = 32'd1199
; 
32'd142514: dataIn1 = 32'd1204
; 
32'd142515: dataIn1 = 32'd3528
; 
32'd142516: dataIn1 = 32'd3530
; 
32'd142517: dataIn1 = 32'd3532
; 
32'd142518: dataIn1 = 32'd233
; 
32'd142519: dataIn1 = 32'd1056
; 
32'd142520: dataIn1 = 32'd1090
; 
32'd142521: dataIn1 = 32'd2589
; 
32'd142522: dataIn1 = 32'd3529
; 
32'd142523: dataIn1 = 32'd3531
; 
32'd142524: dataIn1 = 32'd3533
; 
32'd142525: dataIn1 = 32'd4744
; 
32'd142526: dataIn1 = 32'd258
; 
32'd142527: dataIn1 = 32'd525
; 
32'd142528: dataIn1 = 32'd1196
; 
32'd142529: dataIn1 = 32'd1199
; 
32'd142530: dataIn1 = 32'd3530
; 
32'd142531: dataIn1 = 32'd3532
; 
32'd142532: dataIn1 = 32'd3534
; 
32'd142533: dataIn1 = 32'd233
; 
32'd142534: dataIn1 = 32'd1057
; 
32'd142535: dataIn1 = 32'd1091
; 
32'd142536: dataIn1 = 32'd2589
; 
32'd142537: dataIn1 = 32'd3531
; 
32'd142538: dataIn1 = 32'd3533
; 
32'd142539: dataIn1 = 32'd3535
; 
32'd142540: dataIn1 = 32'd4746
; 
32'd142541: dataIn1 = 32'd523
; 
32'd142542: dataIn1 = 32'd525
; 
32'd142543: dataIn1 = 32'd1192
; 
32'd142544: dataIn1 = 32'd1196
; 
32'd142545: dataIn1 = 32'd3532
; 
32'd142546: dataIn1 = 32'd3534
; 
32'd142547: dataIn1 = 32'd3536
; 
32'd142548: dataIn1 = 32'd143
; 
32'd142549: dataIn1 = 32'd1057
; 
32'd142550: dataIn1 = 32'd1091
; 
32'd142551: dataIn1 = 32'd2668
; 
32'd142552: dataIn1 = 32'd3533
; 
32'd142553: dataIn1 = 32'd3535
; 
32'd142554: dataIn1 = 32'd3537
; 
32'd142555: dataIn1 = 32'd5024
; 
32'd142556: dataIn1 = 32'd523
; 
32'd142557: dataIn1 = 32'd524
; 
32'd142558: dataIn1 = 32'd1192
; 
32'd142559: dataIn1 = 32'd1197
; 
32'd142560: dataIn1 = 32'd3534
; 
32'd142561: dataIn1 = 32'd3536
; 
32'd142562: dataIn1 = 32'd3538
; 
32'd142563: dataIn1 = 32'd143
; 
32'd142564: dataIn1 = 32'd1058
; 
32'd142565: dataIn1 = 32'd1092
; 
32'd142566: dataIn1 = 32'd2668
; 
32'd142567: dataIn1 = 32'd3535
; 
32'd142568: dataIn1 = 32'd3537
; 
32'd142569: dataIn1 = 32'd3539
; 
32'd142570: dataIn1 = 32'd5021
; 
32'd142571: dataIn1 = 32'd257
; 
32'd142572: dataIn1 = 32'd524
; 
32'd142573: dataIn1 = 32'd1197
; 
32'd142574: dataIn1 = 32'd1198
; 
32'd142575: dataIn1 = 32'd3536
; 
32'd142576: dataIn1 = 32'd3538
; 
32'd142577: dataIn1 = 32'd3540
; 
32'd142578: dataIn1 = 32'd236
; 
32'd142579: dataIn1 = 32'd1058
; 
32'd142580: dataIn1 = 32'd1092
; 
32'd142581: dataIn1 = 32'd2593
; 
32'd142582: dataIn1 = 32'd3537
; 
32'd142583: dataIn1 = 32'd3539
; 
32'd142584: dataIn1 = 32'd3541
; 
32'd142585: dataIn1 = 32'd4751
; 
32'd142586: dataIn1 = 32'd257
; 
32'd142587: dataIn1 = 32'd518
; 
32'd142588: dataIn1 = 32'd1180
; 
32'd142589: dataIn1 = 32'd1198
; 
32'd142590: dataIn1 = 32'd3538
; 
32'd142591: dataIn1 = 32'd3540
; 
32'd142592: dataIn1 = 32'd3542
; 
32'd142593: dataIn1 = 32'd236
; 
32'd142594: dataIn1 = 32'd1059
; 
32'd142595: dataIn1 = 32'd1093
; 
32'd142596: dataIn1 = 32'd2593
; 
32'd142597: dataIn1 = 32'd3539
; 
32'd142598: dataIn1 = 32'd3541
; 
32'd142599: dataIn1 = 32'd3543
; 
32'd142600: dataIn1 = 32'd4754
; 
32'd142601: dataIn1 = 32'd517
; 
32'd142602: dataIn1 = 32'd518
; 
32'd142603: dataIn1 = 32'd1180
; 
32'd142604: dataIn1 = 32'd1183
; 
32'd142605: dataIn1 = 32'd3540
; 
32'd142606: dataIn1 = 32'd3542
; 
32'd142607: dataIn1 = 32'd3544
; 
32'd142608: dataIn1 = 32'd144
; 
32'd142609: dataIn1 = 32'd1059
; 
32'd142610: dataIn1 = 32'd1093
; 
32'd142611: dataIn1 = 32'd2674
; 
32'd142612: dataIn1 = 32'd3541
; 
32'd142613: dataIn1 = 32'd3543
; 
32'd142614: dataIn1 = 32'd3545
; 
32'd142615: dataIn1 = 32'd5039
; 
32'd142616: dataIn1 = 32'd517
; 
32'd142617: dataIn1 = 32'd519
; 
32'd142618: dataIn1 = 32'd1179
; 
32'd142619: dataIn1 = 32'd1183
; 
32'd142620: dataIn1 = 32'd3542
; 
32'd142621: dataIn1 = 32'd3544
; 
32'd142622: dataIn1 = 32'd3546
; 
32'd142623: dataIn1 = 32'd144
; 
32'd142624: dataIn1 = 32'd1060
; 
32'd142625: dataIn1 = 32'd1094
; 
32'd142626: dataIn1 = 32'd2674
; 
32'd142627: dataIn1 = 32'd3543
; 
32'd142628: dataIn1 = 32'd3545
; 
32'd142629: dataIn1 = 32'd3547
; 
32'd142630: dataIn1 = 32'd5041
; 
32'd142631: dataIn1 = 32'd256
; 
32'd142632: dataIn1 = 32'd519
; 
32'd142633: dataIn1 = 32'd1179
; 
32'd142634: dataIn1 = 32'd1187
; 
32'd142635: dataIn1 = 32'd3544
; 
32'd142636: dataIn1 = 32'd3546
; 
32'd142637: dataIn1 = 32'd3548
; 
32'd142638: dataIn1 = 32'd239
; 
32'd142639: dataIn1 = 32'd1060
; 
32'd142640: dataIn1 = 32'd1094
; 
32'd142641: dataIn1 = 32'd2595
; 
32'd142642: dataIn1 = 32'd3545
; 
32'd142643: dataIn1 = 32'd3547
; 
32'd142644: dataIn1 = 32'd3549
; 
32'd142645: dataIn1 = 32'd4762
; 
32'd142646: dataIn1 = 32'd256
; 
32'd142647: dataIn1 = 32'd521
; 
32'd142648: dataIn1 = 32'd1187
; 
32'd142649: dataIn1 = 32'd1190
; 
32'd142650: dataIn1 = 32'd3546
; 
32'd142651: dataIn1 = 32'd3548
; 
32'd142652: dataIn1 = 32'd3550
; 
32'd142653: dataIn1 = 32'd239
; 
32'd142654: dataIn1 = 32'd1061
; 
32'd142655: dataIn1 = 32'd1095
; 
32'd142656: dataIn1 = 32'd2595
; 
32'd142657: dataIn1 = 32'd3547
; 
32'd142658: dataIn1 = 32'd3549
; 
32'd142659: dataIn1 = 32'd3551
; 
32'd142660: dataIn1 = 32'd4764
; 
32'd142661: dataIn1 = 32'd521
; 
32'd142662: dataIn1 = 32'd522
; 
32'd142663: dataIn1 = 32'd1185
; 
32'd142664: dataIn1 = 32'd1190
; 
32'd142665: dataIn1 = 32'd3548
; 
32'd142666: dataIn1 = 32'd3550
; 
32'd142667: dataIn1 = 32'd3552
; 
32'd142668: dataIn1 = 32'd146
; 
32'd142669: dataIn1 = 32'd1061
; 
32'd142670: dataIn1 = 32'd1095
; 
32'd142671: dataIn1 = 32'd2678
; 
32'd142672: dataIn1 = 32'd3549
; 
32'd142673: dataIn1 = 32'd3551
; 
32'd142674: dataIn1 = 32'd3553
; 
32'd142675: dataIn1 = 32'd5062
; 
32'd142676: dataIn1 = 32'd520
; 
32'd142677: dataIn1 = 32'd522
; 
32'd142678: dataIn1 = 32'd1185
; 
32'd142679: dataIn1 = 32'd1191
; 
32'd142680: dataIn1 = 32'd3550
; 
32'd142681: dataIn1 = 32'd3552
; 
32'd142682: dataIn1 = 32'd3554
; 
32'd142683: dataIn1 = 32'd146
; 
32'd142684: dataIn1 = 32'd1062
; 
32'd142685: dataIn1 = 32'd1096
; 
32'd142686: dataIn1 = 32'd2678
; 
32'd142687: dataIn1 = 32'd3551
; 
32'd142688: dataIn1 = 32'd3553
; 
32'd142689: dataIn1 = 32'd3555
; 
32'd142690: dataIn1 = 32'd5059
; 
32'd142691: dataIn1 = 32'd251
; 
32'd142692: dataIn1 = 32'd520
; 
32'd142693: dataIn1 = 32'd1186
; 
32'd142694: dataIn1 = 32'd1191
; 
32'd142695: dataIn1 = 32'd3552
; 
32'd142696: dataIn1 = 32'd3554
; 
32'd142697: dataIn1 = 32'd3556
; 
32'd142698: dataIn1 = 32'd242
; 
32'd142699: dataIn1 = 32'd1062
; 
32'd142700: dataIn1 = 32'd1096
; 
32'd142701: dataIn1 = 32'd2599
; 
32'd142702: dataIn1 = 32'd3553
; 
32'd142703: dataIn1 = 32'd3555
; 
32'd142704: dataIn1 = 32'd3557
; 
32'd142705: dataIn1 = 32'd4769
; 
32'd142706: dataIn1 = 32'd251
; 
32'd142707: dataIn1 = 32'd506
; 
32'd142708: dataIn1 = 32'd1146
; 
32'd142709: dataIn1 = 32'd1186
; 
32'd142710: dataIn1 = 32'd3554
; 
32'd142711: dataIn1 = 32'd3556
; 
32'd142712: dataIn1 = 32'd3558
; 
32'd142713: dataIn1 = 32'd242
; 
32'd142714: dataIn1 = 32'd1063
; 
32'd142715: dataIn1 = 32'd1097
; 
32'd142716: dataIn1 = 32'd2599
; 
32'd142717: dataIn1 = 32'd3555
; 
32'd142718: dataIn1 = 32'd3557
; 
32'd142719: dataIn1 = 32'd3559
; 
32'd142720: dataIn1 = 32'd4772
; 
32'd142721: dataIn1 = 32'd504
; 
32'd142722: dataIn1 = 32'd506
; 
32'd142723: dataIn1 = 32'd1146
; 
32'd142724: dataIn1 = 32'd1149
; 
32'd142725: dataIn1 = 32'd3556
; 
32'd142726: dataIn1 = 32'd3558
; 
32'd142727: dataIn1 = 32'd3560
; 
32'd142728: dataIn1 = 32'd147
; 
32'd142729: dataIn1 = 32'd1063
; 
32'd142730: dataIn1 = 32'd1097
; 
32'd142731: dataIn1 = 32'd2684
; 
32'd142732: dataIn1 = 32'd3557
; 
32'd142733: dataIn1 = 32'd3559
; 
32'd142734: dataIn1 = 32'd3561
; 
32'd142735: dataIn1 = 32'd5077
; 
32'd142736: dataIn1 = 32'd504
; 
32'd142737: dataIn1 = 32'd505
; 
32'd142738: dataIn1 = 32'd1148
; 
32'd142739: dataIn1 = 32'd1149
; 
32'd142740: dataIn1 = 32'd3558
; 
32'd142741: dataIn1 = 32'd3560
; 
32'd142742: dataIn1 = 32'd3562
; 
32'd142743: dataIn1 = 32'd147
; 
32'd142744: dataIn1 = 32'd1064
; 
32'd142745: dataIn1 = 32'd1098
; 
32'd142746: dataIn1 = 32'd2684
; 
32'd142747: dataIn1 = 32'd3559
; 
32'd142748: dataIn1 = 32'd3561
; 
32'd142749: dataIn1 = 32'd3563
; 
32'd142750: dataIn1 = 32'd5079
; 
32'd142751: dataIn1 = 32'd252
; 
32'd142752: dataIn1 = 32'd505
; 
32'd142753: dataIn1 = 32'd1148
; 
32'd142754: dataIn1 = 32'd1162
; 
32'd142755: dataIn1 = 32'd3560
; 
32'd142756: dataIn1 = 32'd3562
; 
32'd142757: dataIn1 = 32'd3564
; 
32'd142758: dataIn1 = 32'd245
; 
32'd142759: dataIn1 = 32'd1064
; 
32'd142760: dataIn1 = 32'd1098
; 
32'd142761: dataIn1 = 32'd2601
; 
32'd142762: dataIn1 = 32'd3561
; 
32'd142763: dataIn1 = 32'd3563
; 
32'd142764: dataIn1 = 32'd3565
; 
32'd142765: dataIn1 = 32'd4780
; 
32'd142766: dataIn1 = 32'd252
; 
32'd142767: dataIn1 = 32'd510
; 
32'd142768: dataIn1 = 32'd1162
; 
32'd142769: dataIn1 = 32'd1166
; 
32'd142770: dataIn1 = 32'd3562
; 
32'd142771: dataIn1 = 32'd3564
; 
32'd142772: dataIn1 = 32'd3566
; 
32'd142773: dataIn1 = 32'd245
; 
32'd142774: dataIn1 = 32'd1065
; 
32'd142775: dataIn1 = 32'd1099
; 
32'd142776: dataIn1 = 32'd2601
; 
32'd142777: dataIn1 = 32'd3563
; 
32'd142778: dataIn1 = 32'd3565
; 
32'd142779: dataIn1 = 32'd3567
; 
32'd142780: dataIn1 = 32'd4782
; 
32'd142781: dataIn1 = 32'd510
; 
32'd142782: dataIn1 = 32'd511
; 
32'd142783: dataIn1 = 32'd1161
; 
32'd142784: dataIn1 = 32'd1166
; 
32'd142785: dataIn1 = 32'd3564
; 
32'd142786: dataIn1 = 32'd3566
; 
32'd142787: dataIn1 = 32'd3568
; 
32'd142788: dataIn1 = 32'd149
; 
32'd142789: dataIn1 = 32'd1065
; 
32'd142790: dataIn1 = 32'd1099
; 
32'd142791: dataIn1 = 32'd2688
; 
32'd142792: dataIn1 = 32'd3565
; 
32'd142793: dataIn1 = 32'd3567
; 
32'd142794: dataIn1 = 32'd3569
; 
32'd142795: dataIn1 = 32'd5100
; 
32'd142796: dataIn1 = 32'd511
; 
32'd142797: dataIn1 = 32'd512
; 
32'd142798: dataIn1 = 32'd1161
; 
32'd142799: dataIn1 = 32'd1165
; 
32'd142800: dataIn1 = 32'd3566
; 
32'd142801: dataIn1 = 32'd3568
; 
32'd142802: dataIn1 = 32'd3570
; 
32'd142803: dataIn1 = 32'd149
; 
32'd142804: dataIn1 = 32'd1066
; 
32'd142805: dataIn1 = 32'd1100
; 
32'd142806: dataIn1 = 32'd2688
; 
32'd142807: dataIn1 = 32'd3567
; 
32'd142808: dataIn1 = 32'd3569
; 
32'd142809: dataIn1 = 32'd3571
; 
32'd142810: dataIn1 = 32'd5097
; 
32'd142811: dataIn1 = 32'd253
; 
32'd142812: dataIn1 = 32'd512
; 
32'd142813: dataIn1 = 32'd1165
; 
32'd142814: dataIn1 = 32'd1167
; 
32'd142815: dataIn1 = 32'd3568
; 
32'd142816: dataIn1 = 32'd3570
; 
32'd142817: dataIn1 = 32'd3572
; 
32'd142818: dataIn1 = 32'd248
; 
32'd142819: dataIn1 = 32'd1066
; 
32'd142820: dataIn1 = 32'd1100
; 
32'd142821: dataIn1 = 32'd3569
; 
32'd142822: dataIn1 = 32'd3571
; 
32'd142823: dataIn1 = 32'd3573
; 
32'd142824: dataIn1 = 32'd4787
; 
32'd142825: dataIn1 = 32'd253
; 
32'd142826: dataIn1 = 32'd509
; 
32'd142827: dataIn1 = 32'd1154
; 
32'd142828: dataIn1 = 32'd1167
; 
32'd142829: dataIn1 = 32'd3570
; 
32'd142830: dataIn1 = 32'd3572
; 
32'd142831: dataIn1 = 32'd3574
; 
32'd142832: dataIn1 = 32'd248
; 
32'd142833: dataIn1 = 32'd1067
; 
32'd142834: dataIn1 = 32'd2605
; 
32'd142835: dataIn1 = 32'd3571
; 
32'd142836: dataIn1 = 32'd3573
; 
32'd142837: dataIn1 = 32'd3575
; 
32'd142838: dataIn1 = 32'd4787
; 
32'd142839: dataIn1 = 32'd4790
; 
32'd142840: dataIn1 = 32'd507
; 
32'd142841: dataIn1 = 32'd509
; 
32'd142842: dataIn1 = 32'd1154
; 
32'd142843: dataIn1 = 32'd1160
; 
32'd142844: dataIn1 = 32'd3572
; 
32'd142845: dataIn1 = 32'd3574
; 
32'd142846: dataIn1 = 32'd3576
; 
32'd142847: dataIn1 = 32'd150
; 
32'd142848: dataIn1 = 32'd1067
; 
32'd142849: dataIn1 = 32'd1101
; 
32'd142850: dataIn1 = 32'd3573
; 
32'd142851: dataIn1 = 32'd3575
; 
32'd142852: dataIn1 = 32'd4790
; 
32'd142853: dataIn1 = 32'd507
; 
32'd142854: dataIn1 = 32'd508
; 
32'd142855: dataIn1 = 32'd1156
; 
32'd142856: dataIn1 = 32'd1160
; 
32'd142857: dataIn1 = 32'd3574
; 
32'd142858: dataIn1 = 32'd3576
; 
32'd142859: dataIn1 = 32'd3577
; 
32'd142860: dataIn1 = 32'd254
; 
32'd142861: dataIn1 = 32'd508
; 
32'd142862: dataIn1 = 32'd1156
; 
32'd142863: dataIn1 = 32'd1175
; 
32'd142864: dataIn1 = 32'd3576
; 
32'd142865: dataIn1 = 32'd3577
; 
32'd142866: dataIn1 = 32'd3578
; 
32'd142867: dataIn1 = 32'd254
; 
32'd142868: dataIn1 = 32'd515
; 
32'd142869: dataIn1 = 32'd1171
; 
32'd142870: dataIn1 = 32'd1175
; 
32'd142871: dataIn1 = 32'd3577
; 
32'd142872: dataIn1 = 32'd3578
; 
32'd142873: dataIn1 = 32'd3579
; 
32'd142874: dataIn1 = 32'd513
; 
32'd142875: dataIn1 = 32'd515
; 
32'd142876: dataIn1 = 32'd1168
; 
32'd142877: dataIn1 = 32'd1171
; 
32'd142878: dataIn1 = 32'd3578
; 
32'd142879: dataIn1 = 32'd3579
; 
32'd142880: dataIn1 = 32'd3580
; 
32'd142881: dataIn1 = 32'd513
; 
32'd142882: dataIn1 = 32'd514
; 
32'd142883: dataIn1 = 32'd1168
; 
32'd142884: dataIn1 = 32'd1173
; 
32'd142885: dataIn1 = 32'd3579
; 
32'd142886: dataIn1 = 32'd3580
; 
32'd142887: dataIn1 = 32'd3581
; 
32'd142888: dataIn1 = 32'd255
; 
32'd142889: dataIn1 = 32'd514
; 
32'd142890: dataIn1 = 32'd1173
; 
32'd142891: dataIn1 = 32'd1174
; 
32'd142892: dataIn1 = 32'd3580
; 
32'd142893: dataIn1 = 32'd3581
; 
32'd142894: dataIn1 = 32'd3582
; 
32'd142895: dataIn1 = 32'd255
; 
32'd142896: dataIn1 = 32'd516
; 
32'd142897: dataIn1 = 32'd1174
; 
32'd142898: dataIn1 = 32'd3581
; 
32'd142899: dataIn1 = 32'd3582
; 
32'd142900: dataIn1 = 32'd3583
; 
32'd142901: dataIn1 = 32'd6805
; 
32'd142902: dataIn1 = 32'd6806
; 
32'd142903: dataIn1 = 32'd6819
; 
32'd142904: dataIn1 = 32'd6824
; 
32'd142905: dataIn1 = 32'd9265
; 
32'd142906: dataIn1 = 32'd3584
; 
32'd142907: dataIn1 = 32'd9353
; 
32'd142908: dataIn1 = 32'd9354
; 
32'd142909: dataIn1 = 32'd9375
; 
32'd142910: dataIn1 = 32'd9389
; 
32'd142911: dataIn1 = 32'd3585
; 
32'd142912: dataIn1 = 32'd6831
; 
32'd142913: dataIn1 = 32'd6832
; 
32'd142914: dataIn1 = 32'd6845
; 
32'd142915: dataIn1 = 32'd6850
; 
32'd142916: dataIn1 = 32'd9267
; 
32'd142917: dataIn1 = 32'd3586
; 
32'd142918: dataIn1 = 32'd9412
; 
32'd142919: dataIn1 = 32'd9413
; 
32'd142920: dataIn1 = 32'd9434
; 
32'd142921: dataIn1 = 32'd9441
; 
32'd142922: dataIn1 = 32'd3587
; 
32'd142923: dataIn1 = 32'd3591
; 
32'd142924: dataIn1 = 32'd9469
; 
32'd142925: dataIn1 = 32'd9470
; 
32'd142926: dataIn1 = 32'd9474
; 
32'd142927: dataIn1 = 32'd9476
; 
32'd142928: dataIn1 = 32'd9850
; 
32'd142929: dataIn1 = 32'd9859
; 
32'd142930: dataIn1 = 32'd10159
; 
32'd142931: dataIn1 = 32'd3588
; 
32'd142932: dataIn1 = 32'd9853
; 
32'd142933: dataIn1 = 32'd9854
; 
32'd142934: dataIn1 = 32'd9857
; 
32'd142935: dataIn1 = 32'd9909
; 
32'd142936: dataIn1 = 32'd10158
; 
32'd142937: dataIn1 = 32'd10172
; 
32'd142938: dataIn1 = 32'd3589
; 
32'd142939: dataIn1 = 32'd9471
; 
32'd142940: dataIn1 = 32'd9771
; 
32'd142941: dataIn1 = 32'd9855
; 
32'd142942: dataIn1 = 32'd9856
; 
32'd142943: dataIn1 = 32'd9864
; 
32'd142944: dataIn1 = 32'd10160
; 
32'd142945: dataIn1 = 32'd2178
; 
32'd142946: dataIn1 = 32'd3590
; 
32'd142947: dataIn1 = 32'd3591
; 
32'd142948: dataIn1 = 32'd9466
; 
32'd142949: dataIn1 = 32'd9475
; 
32'd142950: dataIn1 = 32'd9476
; 
32'd142951: dataIn1 = 32'd9844
; 
32'd142952: dataIn1 = 32'd52
; 
32'd142953: dataIn1 = 32'd2178
; 
32'd142954: dataIn1 = 32'd3587
; 
32'd142955: dataIn1 = 32'd3590
; 
32'd142956: dataIn1 = 32'd3591
; 
32'd142957: dataIn1 = 32'd3593
; 
32'd142958: dataIn1 = 32'd3597
; 
32'd142959: dataIn1 = 32'd9476
; 
32'd142960: dataIn1 = 32'd10159
; 
32'd142961: dataIn1 = 32'd2178
; 
32'd142962: dataIn1 = 32'd2180
; 
32'd142963: dataIn1 = 32'd3592
; 
32'd142964: dataIn1 = 32'd3593
; 
32'd142965: dataIn1 = 32'd3594
; 
32'd142966: dataIn1 = 32'd3595
; 
32'd142967: dataIn1 = 32'd3596
; 
32'd142968: dataIn1 = 32'd2178
; 
32'd142969: dataIn1 = 32'd2179
; 
32'd142970: dataIn1 = 32'd3591
; 
32'd142971: dataIn1 = 32'd3592
; 
32'd142972: dataIn1 = 32'd3593
; 
32'd142973: dataIn1 = 32'd3594
; 
32'd142974: dataIn1 = 32'd3597
; 
32'd142975: dataIn1 = 32'd2179
; 
32'd142976: dataIn1 = 32'd2180
; 
32'd142977: dataIn1 = 32'd3592
; 
32'd142978: dataIn1 = 32'd3593
; 
32'd142979: dataIn1 = 32'd3594
; 
32'd142980: dataIn1 = 32'd3598
; 
32'd142981: dataIn1 = 32'd3599
; 
32'd142982: dataIn1 = 32'd42
; 
32'd142983: dataIn1 = 32'd2178
; 
32'd142984: dataIn1 = 32'd3592
; 
32'd142985: dataIn1 = 32'd3595
; 
32'd142986: dataIn1 = 32'd3596
; 
32'd142987: dataIn1 = 32'd9466
; 
32'd142988: dataIn1 = 32'd9477
; 
32'd142989: dataIn1 = 32'd42
; 
32'd142990: dataIn1 = 32'd2180
; 
32'd142991: dataIn1 = 32'd3592
; 
32'd142992: dataIn1 = 32'd3595
; 
32'd142993: dataIn1 = 32'd3596
; 
32'd142994: dataIn1 = 32'd3600
; 
32'd142995: dataIn1 = 32'd3603
; 
32'd142996: dataIn1 = 32'd52
; 
32'd142997: dataIn1 = 32'd2179
; 
32'd142998: dataIn1 = 32'd3591
; 
32'd142999: dataIn1 = 32'd3593
; 
32'd143000: dataIn1 = 32'd3597
; 
32'd143001: dataIn1 = 32'd3637
; 
32'd143002: dataIn1 = 32'd3641
; 
32'd143003: dataIn1 = 32'd53
; 
32'd143004: dataIn1 = 32'd2180
; 
32'd143005: dataIn1 = 32'd3594
; 
32'd143006: dataIn1 = 32'd3598
; 
32'd143007: dataIn1 = 32'd3599
; 
32'd143008: dataIn1 = 32'd3601
; 
32'd143009: dataIn1 = 32'd3604
; 
32'd143010: dataIn1 = 32'd53
; 
32'd143011: dataIn1 = 32'd2179
; 
32'd143012: dataIn1 = 32'd3594
; 
32'd143013: dataIn1 = 32'd3598
; 
32'd143014: dataIn1 = 32'd3599
; 
32'd143015: dataIn1 = 32'd3643
; 
32'd143016: dataIn1 = 32'd3645
; 
32'd143017: dataIn1 = 32'd2151
; 
32'd143018: dataIn1 = 32'd2180
; 
32'd143019: dataIn1 = 32'd3596
; 
32'd143020: dataIn1 = 32'd3600
; 
32'd143021: dataIn1 = 32'd3601
; 
32'd143022: dataIn1 = 32'd3602
; 
32'd143023: dataIn1 = 32'd3603
; 
32'd143024: dataIn1 = 32'd2180
; 
32'd143025: dataIn1 = 32'd2181
; 
32'd143026: dataIn1 = 32'd3598
; 
32'd143027: dataIn1 = 32'd3600
; 
32'd143028: dataIn1 = 32'd3601
; 
32'd143029: dataIn1 = 32'd3602
; 
32'd143030: dataIn1 = 32'd3604
; 
32'd143031: dataIn1 = 32'd2151
; 
32'd143032: dataIn1 = 32'd2181
; 
32'd143033: dataIn1 = 32'd3600
; 
32'd143034: dataIn1 = 32'd3601
; 
32'd143035: dataIn1 = 32'd3602
; 
32'd143036: dataIn1 = 32'd3605
; 
32'd143037: dataIn1 = 32'd3606
; 
32'd143038: dataIn1 = 32'd42
; 
32'd143039: dataIn1 = 32'd2150
; 
32'd143040: dataIn1 = 32'd2151
; 
32'd143041: dataIn1 = 32'd3596
; 
32'd143042: dataIn1 = 32'd3600
; 
32'd143043: dataIn1 = 32'd3603
; 
32'd143044: dataIn1 = 32'd53
; 
32'd143045: dataIn1 = 32'd2181
; 
32'd143046: dataIn1 = 32'd3598
; 
32'd143047: dataIn1 = 32'd3601
; 
32'd143048: dataIn1 = 32'd3604
; 
32'd143049: dataIn1 = 32'd3608
; 
32'd143050: dataIn1 = 32'd3610
; 
32'd143051: dataIn1 = 32'd43
; 
32'd143052: dataIn1 = 32'd2151
; 
32'd143053: dataIn1 = 32'd2152
; 
32'd143054: dataIn1 = 32'd3602
; 
32'd143055: dataIn1 = 32'd3605
; 
32'd143056: dataIn1 = 32'd3606
; 
32'd143057: dataIn1 = 32'd43
; 
32'd143058: dataIn1 = 32'd2181
; 
32'd143059: dataIn1 = 32'd3602
; 
32'd143060: dataIn1 = 32'd3605
; 
32'd143061: dataIn1 = 32'd3606
; 
32'd143062: dataIn1 = 32'd3607
; 
32'd143063: dataIn1 = 32'd5308
; 
32'd143064: dataIn1 = 32'd2181
; 
32'd143065: dataIn1 = 32'd2183
; 
32'd143066: dataIn1 = 32'd3606
; 
32'd143067: dataIn1 = 32'd3607
; 
32'd143068: dataIn1 = 32'd3608
; 
32'd143069: dataIn1 = 32'd3609
; 
32'd143070: dataIn1 = 32'd5308
; 
32'd143071: dataIn1 = 32'd2181
; 
32'd143072: dataIn1 = 32'd2182
; 
32'd143073: dataIn1 = 32'd3604
; 
32'd143074: dataIn1 = 32'd3607
; 
32'd143075: dataIn1 = 32'd3608
; 
32'd143076: dataIn1 = 32'd3609
; 
32'd143077: dataIn1 = 32'd3610
; 
32'd143078: dataIn1 = 32'd54
; 
32'd143079: dataIn1 = 32'd2182
; 
32'd143080: dataIn1 = 32'd2183
; 
32'd143081: dataIn1 = 32'd3607
; 
32'd143082: dataIn1 = 32'd3608
; 
32'd143083: dataIn1 = 32'd3609
; 
32'd143084: dataIn1 = 32'd53
; 
32'd143085: dataIn1 = 32'd2182
; 
32'd143086: dataIn1 = 32'd3604
; 
32'd143087: dataIn1 = 32'd3608
; 
32'd143088: dataIn1 = 32'd3610
; 
32'd143089: dataIn1 = 32'd3649
; 
32'd143090: dataIn1 = 32'd3653
; 
32'd143091: dataIn1 = 32'd50
; 
32'd143092: dataIn1 = 32'd2200
; 
32'd143093: dataIn1 = 32'd2202
; 
32'd143094: dataIn1 = 32'd3611
; 
32'd143095: dataIn1 = 32'd3612
; 
32'd143096: dataIn1 = 32'd3613
; 
32'd143097: dataIn1 = 32'd2200
; 
32'd143098: dataIn1 = 32'd2201
; 
32'd143099: dataIn1 = 32'd3611
; 
32'd143100: dataIn1 = 32'd3612
; 
32'd143101: dataIn1 = 32'd3613
; 
32'd143102: dataIn1 = 32'd3614
; 
32'd143103: dataIn1 = 32'd3615
; 
32'd143104: dataIn1 = 32'd2201
; 
32'd143105: dataIn1 = 32'd2202
; 
32'd143106: dataIn1 = 32'd3611
; 
32'd143107: dataIn1 = 32'd3612
; 
32'd143108: dataIn1 = 32'd3613
; 
32'd143109: dataIn1 = 32'd3616
; 
32'd143110: dataIn1 = 32'd3617
; 
32'd143111: dataIn1 = 32'd60
; 
32'd143112: dataIn1 = 32'd2199
; 
32'd143113: dataIn1 = 32'd2200
; 
32'd143114: dataIn1 = 32'd3612
; 
32'd143115: dataIn1 = 32'd3614
; 
32'd143116: dataIn1 = 32'd3615
; 
32'd143117: dataIn1 = 32'd60
; 
32'd143118: dataIn1 = 32'd2201
; 
32'd143119: dataIn1 = 32'd3612
; 
32'd143120: dataIn1 = 32'd3614
; 
32'd143121: dataIn1 = 32'd3615
; 
32'd143122: dataIn1 = 32'd3690
; 
32'd143123: dataIn1 = 32'd3694
; 
32'd143124: dataIn1 = 32'd10192
; 
32'd143125: dataIn1 = 32'd61
; 
32'd143126: dataIn1 = 32'd2202
; 
32'd143127: dataIn1 = 32'd3613
; 
32'd143128: dataIn1 = 32'd3616
; 
32'd143129: dataIn1 = 32'd3617
; 
32'd143130: dataIn1 = 32'd3618
; 
32'd143131: dataIn1 = 32'd3619
; 
32'd143132: dataIn1 = 32'd9550
; 
32'd143133: dataIn1 = 32'd10196
; 
32'd143134: dataIn1 = 32'd2201
; 
32'd143135: dataIn1 = 32'd3613
; 
32'd143136: dataIn1 = 32'd3616
; 
32'd143137: dataIn1 = 32'd3617
; 
32'd143138: dataIn1 = 32'd9546
; 
32'd143139: dataIn1 = 32'd9547
; 
32'd143140: dataIn1 = 32'd9550
; 
32'd143141: dataIn1 = 32'd2173
; 
32'd143142: dataIn1 = 32'd2202
; 
32'd143143: dataIn1 = 32'd2203
; 
32'd143144: dataIn1 = 32'd3616
; 
32'd143145: dataIn1 = 32'd3618
; 
32'd143146: dataIn1 = 32'd3619
; 
32'd143147: dataIn1 = 32'd2203
; 
32'd143148: dataIn1 = 32'd3616
; 
32'd143149: dataIn1 = 32'd3618
; 
32'd143150: dataIn1 = 32'd3619
; 
32'd143151: dataIn1 = 32'd10164
; 
32'd143152: dataIn1 = 32'd10165
; 
32'd143153: dataIn1 = 32'd10196
; 
32'd143154: dataIn1 = 32'd2203
; 
32'd143155: dataIn1 = 32'd3620
; 
32'd143156: dataIn1 = 32'd3623
; 
32'd143157: dataIn1 = 32'd9479
; 
32'd143158: dataIn1 = 32'd9480
; 
32'd143159: dataIn1 = 32'd9484
; 
32'd143160: dataIn1 = 32'd10229
; 
32'd143161: dataIn1 = 32'd2203
; 
32'd143162: dataIn1 = 32'd3621
; 
32'd143163: dataIn1 = 32'd9480
; 
32'd143164: dataIn1 = 32'd9873
; 
32'd143165: dataIn1 = 32'd9874
; 
32'd143166: dataIn1 = 32'd9881
; 
32'd143167: dataIn1 = 32'd10165
; 
32'd143168: dataIn1 = 32'd3622
; 
32'd143169: dataIn1 = 32'd9867
; 
32'd143170: dataIn1 = 32'd9868
; 
32'd143171: dataIn1 = 32'd9875
; 
32'd143172: dataIn1 = 32'd9876
; 
32'd143173: dataIn1 = 32'd9889
; 
32'd143174: dataIn1 = 32'd10162
; 
32'd143175: dataIn1 = 32'd51
; 
32'd143176: dataIn1 = 32'd2173
; 
32'd143177: dataIn1 = 32'd2203
; 
32'd143178: dataIn1 = 32'd3620
; 
32'd143179: dataIn1 = 32'd3623
; 
32'd143180: dataIn1 = 32'd3624
; 
32'd143181: dataIn1 = 32'd10229
; 
32'd143182: dataIn1 = 32'd51
; 
32'd143183: dataIn1 = 32'd3623
; 
32'd143184: dataIn1 = 32'd3624
; 
32'd143185: dataIn1 = 32'd3631
; 
32'd143186: dataIn1 = 32'd10169
; 
32'd143187: dataIn1 = 32'd10170
; 
32'd143188: dataIn1 = 32'd10229
; 
32'd143189: dataIn1 = 32'd3625
; 
32'd143190: dataIn1 = 32'd9882
; 
32'd143191: dataIn1 = 32'd9883
; 
32'd143192: dataIn1 = 32'd10018
; 
32'd143193: dataIn1 = 32'd10019
; 
32'd143194: dataIn1 = 32'd10025
; 
32'd143195: dataIn1 = 32'd10164
; 
32'd143196: dataIn1 = 32'd62
; 
32'd143197: dataIn1 = 32'd3626
; 
32'd143198: dataIn1 = 32'd3632
; 
32'd143199: dataIn1 = 32'd9487
; 
32'd143200: dataIn1 = 32'd9488
; 
32'd143201: dataIn1 = 32'd9496
; 
32'd143202: dataIn1 = 32'd9884
; 
32'd143203: dataIn1 = 32'd10166
; 
32'd143204: dataIn1 = 32'd62
; 
32'd143205: dataIn1 = 32'd3627
; 
32'd143206: dataIn1 = 32'd3708
; 
32'd143207: dataIn1 = 32'd3710
; 
32'd143208: dataIn1 = 32'd10162
; 
32'd143209: dataIn1 = 32'd10163
; 
32'd143210: dataIn1 = 32'd10166
; 
32'd143211: dataIn1 = 32'd3628
; 
32'd143212: dataIn1 = 32'd3631
; 
32'd143213: dataIn1 = 32'd9493
; 
32'd143214: dataIn1 = 32'd9893
; 
32'd143215: dataIn1 = 32'd9894
; 
32'd143216: dataIn1 = 32'd9902
; 
32'd143217: dataIn1 = 32'd10170
; 
32'd143218: dataIn1 = 32'd3629
; 
32'd143219: dataIn1 = 32'd3632
; 
32'd143220: dataIn1 = 32'd9489
; 
32'd143221: dataIn1 = 32'd9491
; 
32'd143222: dataIn1 = 32'd9494
; 
32'd143223: dataIn1 = 32'd9496
; 
32'd143224: dataIn1 = 32'd9891
; 
32'd143225: dataIn1 = 32'd9900
; 
32'd143226: dataIn1 = 32'd10168
; 
32'd143227: dataIn1 = 32'd3630
; 
32'd143228: dataIn1 = 32'd9895
; 
32'd143229: dataIn1 = 32'd9896
; 
32'd143230: dataIn1 = 32'd9897
; 
32'd143231: dataIn1 = 32'd9910
; 
32'd143232: dataIn1 = 32'd10167
; 
32'd143233: dataIn1 = 32'd10171
; 
32'd143234: dataIn1 = 32'd51
; 
32'd143235: dataIn1 = 32'd2176
; 
32'd143236: dataIn1 = 32'd3624
; 
32'd143237: dataIn1 = 32'd3628
; 
32'd143238: dataIn1 = 32'd3631
; 
32'd143239: dataIn1 = 32'd9493
; 
32'd143240: dataIn1 = 32'd9771
; 
32'd143241: dataIn1 = 32'd9780
; 
32'd143242: dataIn1 = 32'd10170
; 
32'd143243: dataIn1 = 32'd62
; 
32'd143244: dataIn1 = 32'd2206
; 
32'd143245: dataIn1 = 32'd3626
; 
32'd143246: dataIn1 = 32'd3629
; 
32'd143247: dataIn1 = 32'd3632
; 
32'd143248: dataIn1 = 32'd3635
; 
32'd143249: dataIn1 = 32'd3638
; 
32'd143250: dataIn1 = 32'd9496
; 
32'd143251: dataIn1 = 32'd10168
; 
32'd143252: dataIn1 = 32'd3633
; 
32'd143253: dataIn1 = 32'd3634
; 
32'd143254: dataIn1 = 32'd3637
; 
32'd143255: dataIn1 = 32'd10171
; 
32'd143256: dataIn1 = 32'd10172
; 
32'd143257: dataIn1 = 32'd10226
; 
32'd143258: dataIn1 = 32'd10228
; 
32'd143259: dataIn1 = 32'd2206
; 
32'd143260: dataIn1 = 32'd2208
; 
32'd143261: dataIn1 = 32'd3633
; 
32'd143262: dataIn1 = 32'd3634
; 
32'd143263: dataIn1 = 32'd3635
; 
32'd143264: dataIn1 = 32'd3636
; 
32'd143265: dataIn1 = 32'd3637
; 
32'd143266: dataIn1 = 32'd10228
; 
32'd143267: dataIn1 = 32'd2206
; 
32'd143268: dataIn1 = 32'd2207
; 
32'd143269: dataIn1 = 32'd3632
; 
32'd143270: dataIn1 = 32'd3634
; 
32'd143271: dataIn1 = 32'd3635
; 
32'd143272: dataIn1 = 32'd3636
; 
32'd143273: dataIn1 = 32'd3638
; 
32'd143274: dataIn1 = 32'd2207
; 
32'd143275: dataIn1 = 32'd2208
; 
32'd143276: dataIn1 = 32'd3634
; 
32'd143277: dataIn1 = 32'd3635
; 
32'd143278: dataIn1 = 32'd3636
; 
32'd143279: dataIn1 = 32'd3639
; 
32'd143280: dataIn1 = 32'd3640
; 
32'd143281: dataIn1 = 32'd52
; 
32'd143282: dataIn1 = 32'd2208
; 
32'd143283: dataIn1 = 32'd3597
; 
32'd143284: dataIn1 = 32'd3633
; 
32'd143285: dataIn1 = 32'd3634
; 
32'd143286: dataIn1 = 32'd3637
; 
32'd143287: dataIn1 = 32'd3641
; 
32'd143288: dataIn1 = 32'd10226
; 
32'd143289: dataIn1 = 32'd62
; 
32'd143290: dataIn1 = 32'd2207
; 
32'd143291: dataIn1 = 32'd3632
; 
32'd143292: dataIn1 = 32'd3635
; 
32'd143293: dataIn1 = 32'd3638
; 
32'd143294: dataIn1 = 32'd3714
; 
32'd143295: dataIn1 = 32'd3718
; 
32'd143296: dataIn1 = 32'd63
; 
32'd143297: dataIn1 = 32'd2208
; 
32'd143298: dataIn1 = 32'd3636
; 
32'd143299: dataIn1 = 32'd3639
; 
32'd143300: dataIn1 = 32'd3640
; 
32'd143301: dataIn1 = 32'd3642
; 
32'd143302: dataIn1 = 32'd3644
; 
32'd143303: dataIn1 = 32'd63
; 
32'd143304: dataIn1 = 32'd2207
; 
32'd143305: dataIn1 = 32'd3636
; 
32'd143306: dataIn1 = 32'd3639
; 
32'd143307: dataIn1 = 32'd3640
; 
32'd143308: dataIn1 = 32'd3720
; 
32'd143309: dataIn1 = 32'd3722
; 
32'd143310: dataIn1 = 32'd2179
; 
32'd143311: dataIn1 = 32'd2208
; 
32'd143312: dataIn1 = 32'd3597
; 
32'd143313: dataIn1 = 32'd3637
; 
32'd143314: dataIn1 = 32'd3641
; 
32'd143315: dataIn1 = 32'd3642
; 
32'd143316: dataIn1 = 32'd3643
; 
32'd143317: dataIn1 = 32'd2208
; 
32'd143318: dataIn1 = 32'd2209
; 
32'd143319: dataIn1 = 32'd3639
; 
32'd143320: dataIn1 = 32'd3641
; 
32'd143321: dataIn1 = 32'd3642
; 
32'd143322: dataIn1 = 32'd3643
; 
32'd143323: dataIn1 = 32'd3644
; 
32'd143324: dataIn1 = 32'd2179
; 
32'd143325: dataIn1 = 32'd2209
; 
32'd143326: dataIn1 = 32'd3599
; 
32'd143327: dataIn1 = 32'd3641
; 
32'd143328: dataIn1 = 32'd3642
; 
32'd143329: dataIn1 = 32'd3643
; 
32'd143330: dataIn1 = 32'd3645
; 
32'd143331: dataIn1 = 32'd63
; 
32'd143332: dataIn1 = 32'd2209
; 
32'd143333: dataIn1 = 32'd3639
; 
32'd143334: dataIn1 = 32'd3642
; 
32'd143335: dataIn1 = 32'd3644
; 
32'd143336: dataIn1 = 32'd3647
; 
32'd143337: dataIn1 = 32'd3650
; 
32'd143338: dataIn1 = 32'd53
; 
32'd143339: dataIn1 = 32'd2209
; 
32'd143340: dataIn1 = 32'd3599
; 
32'd143341: dataIn1 = 32'd3643
; 
32'd143342: dataIn1 = 32'd3645
; 
32'd143343: dataIn1 = 32'd3646
; 
32'd143344: dataIn1 = 32'd3649
; 
32'd143345: dataIn1 = 32'd2209
; 
32'd143346: dataIn1 = 32'd2211
; 
32'd143347: dataIn1 = 32'd3645
; 
32'd143348: dataIn1 = 32'd3646
; 
32'd143349: dataIn1 = 32'd3647
; 
32'd143350: dataIn1 = 32'd3648
; 
32'd143351: dataIn1 = 32'd3649
; 
32'd143352: dataIn1 = 32'd2209
; 
32'd143353: dataIn1 = 32'd2210
; 
32'd143354: dataIn1 = 32'd3644
; 
32'd143355: dataIn1 = 32'd3646
; 
32'd143356: dataIn1 = 32'd3647
; 
32'd143357: dataIn1 = 32'd3648
; 
32'd143358: dataIn1 = 32'd3650
; 
32'd143359: dataIn1 = 32'd2210
; 
32'd143360: dataIn1 = 32'd2211
; 
32'd143361: dataIn1 = 32'd3646
; 
32'd143362: dataIn1 = 32'd3647
; 
32'd143363: dataIn1 = 32'd3648
; 
32'd143364: dataIn1 = 32'd3651
; 
32'd143365: dataIn1 = 32'd3652
; 
32'd143366: dataIn1 = 32'd53
; 
32'd143367: dataIn1 = 32'd2211
; 
32'd143368: dataIn1 = 32'd3610
; 
32'd143369: dataIn1 = 32'd3645
; 
32'd143370: dataIn1 = 32'd3646
; 
32'd143371: dataIn1 = 32'd3649
; 
32'd143372: dataIn1 = 32'd3653
; 
32'd143373: dataIn1 = 32'd63
; 
32'd143374: dataIn1 = 32'd2210
; 
32'd143375: dataIn1 = 32'd3644
; 
32'd143376: dataIn1 = 32'd3647
; 
32'd143377: dataIn1 = 32'd3650
; 
32'd143378: dataIn1 = 32'd3726
; 
32'd143379: dataIn1 = 32'd3728
; 
32'd143380: dataIn1 = 32'd64
; 
32'd143381: dataIn1 = 32'd2211
; 
32'd143382: dataIn1 = 32'd3648
; 
32'd143383: dataIn1 = 32'd3651
; 
32'd143384: dataIn1 = 32'd3652
; 
32'd143385: dataIn1 = 32'd3654
; 
32'd143386: dataIn1 = 32'd3655
; 
32'd143387: dataIn1 = 32'd64
; 
32'd143388: dataIn1 = 32'd2210
; 
32'd143389: dataIn1 = 32'd3648
; 
32'd143390: dataIn1 = 32'd3651
; 
32'd143391: dataIn1 = 32'd3652
; 
32'd143392: dataIn1 = 32'd3730
; 
32'd143393: dataIn1 = 32'd3731
; 
32'd143394: dataIn1 = 32'd2182
; 
32'd143395: dataIn1 = 32'd2211
; 
32'd143396: dataIn1 = 32'd3610
; 
32'd143397: dataIn1 = 32'd3649
; 
32'd143398: dataIn1 = 32'd3653
; 
32'd143399: dataIn1 = 32'd3654
; 
32'd143400: dataIn1 = 32'd5309
; 
32'd143401: dataIn1 = 32'd2211
; 
32'd143402: dataIn1 = 32'd2212
; 
32'd143403: dataIn1 = 32'd3651
; 
32'd143404: dataIn1 = 32'd3653
; 
32'd143405: dataIn1 = 32'd3654
; 
32'd143406: dataIn1 = 32'd3655
; 
32'd143407: dataIn1 = 32'd5309
; 
32'd143408: dataIn1 = 32'd64
; 
32'd143409: dataIn1 = 32'd2212
; 
32'd143410: dataIn1 = 32'd2213
; 
32'd143411: dataIn1 = 32'd3651
; 
32'd143412: dataIn1 = 32'd3654
; 
32'd143413: dataIn1 = 32'd3655
; 
32'd143414: dataIn1 = 32'd66
; 
32'd143415: dataIn1 = 32'd2216
; 
32'd143416: dataIn1 = 32'd3656
; 
32'd143417: dataIn1 = 32'd3657
; 
32'd143418: dataIn1 = 32'd3658
; 
32'd143419: dataIn1 = 32'd55
; 
32'd143420: dataIn1 = 32'd2185
; 
32'd143421: dataIn1 = 32'd2215
; 
32'd143422: dataIn1 = 32'd2216
; 
32'd143423: dataIn1 = 32'd3656
; 
32'd143424: dataIn1 = 32'd3657
; 
32'd143425: dataIn1 = 32'd3658
; 
32'd143426: dataIn1 = 32'd66
; 
32'd143427: dataIn1 = 32'd2215
; 
32'd143428: dataIn1 = 32'd3656
; 
32'd143429: dataIn1 = 32'd3657
; 
32'd143430: dataIn1 = 32'd3658
; 
32'd143431: dataIn1 = 32'd3744
; 
32'd143432: dataIn1 = 32'd5310
; 
32'd143433: dataIn1 = 32'd9567
; 
32'd143434: dataIn1 = 32'd2221
; 
32'd143435: dataIn1 = 32'd3659
; 
32'd143436: dataIn1 = 32'd3662
; 
32'd143437: dataIn1 = 32'd10213
; 
32'd143438: dataIn1 = 32'd10214
; 
32'd143439: dataIn1 = 32'd10242
; 
32'd143440: dataIn1 = 32'd10243
; 
32'd143441: dataIn1 = 32'd3660
; 
32'd143442: dataIn1 = 32'd10083
; 
32'd143443: dataIn1 = 32'd10084
; 
32'd143444: dataIn1 = 32'd10088
; 
32'd143445: dataIn1 = 32'd10093
; 
32'd143446: dataIn1 = 32'd10211
; 
32'd143447: dataIn1 = 32'd10214
; 
32'd143448: dataIn1 = 32'd2221
; 
32'd143449: dataIn1 = 32'd3661
; 
32'd143450: dataIn1 = 32'd9784
; 
32'd143451: dataIn1 = 32'd10211
; 
32'd143452: dataIn1 = 32'd10212
; 
32'd143453: dataIn1 = 32'd10241
; 
32'd143454: dataIn1 = 32'd10242
; 
32'd143455: dataIn1 = 32'd2192
; 
32'd143456: dataIn1 = 32'd2221
; 
32'd143457: dataIn1 = 32'd2222
; 
32'd143458: dataIn1 = 32'd3659
; 
32'd143459: dataIn1 = 32'd3662
; 
32'd143460: dataIn1 = 32'd3663
; 
32'd143461: dataIn1 = 32'd10243
; 
32'd143462: dataIn1 = 32'd2222
; 
32'd143463: dataIn1 = 32'd3662
; 
32'd143464: dataIn1 = 32'd3663
; 
32'd143465: dataIn1 = 32'd10215
; 
32'd143466: dataIn1 = 32'd10216
; 
32'd143467: dataIn1 = 32'd10243
; 
32'd143468: dataIn1 = 32'd10244
; 
32'd143469: dataIn1 = 32'd58
; 
32'd143470: dataIn1 = 32'd2222
; 
32'd143471: dataIn1 = 32'd2224
; 
32'd143472: dataIn1 = 32'd3664
; 
32'd143473: dataIn1 = 32'd3665
; 
32'd143474: dataIn1 = 32'd3666
; 
32'd143475: dataIn1 = 32'd10245
; 
32'd143476: dataIn1 = 32'd2222
; 
32'd143477: dataIn1 = 32'd3664
; 
32'd143478: dataIn1 = 32'd3665
; 
32'd143479: dataIn1 = 32'd10217
; 
32'd143480: dataIn1 = 32'd10218
; 
32'd143481: dataIn1 = 32'd10244
; 
32'd143482: dataIn1 = 32'd10245
; 
32'd143483: dataIn1 = 32'd2224
; 
32'd143484: dataIn1 = 32'd3664
; 
32'd143485: dataIn1 = 32'd3666
; 
32'd143486: dataIn1 = 32'd9498
; 
32'd143487: dataIn1 = 32'd9499
; 
32'd143488: dataIn1 = 32'd9501
; 
32'd143489: dataIn1 = 32'd10245
; 
32'd143490: dataIn1 = 32'd3667
; 
32'd143491: dataIn1 = 32'd10101
; 
32'd143492: dataIn1 = 32'd10102
; 
32'd143493: dataIn1 = 32'd10108
; 
32'd143494: dataIn1 = 32'd10113
; 
32'd143495: dataIn1 = 32'd10215
; 
32'd143496: dataIn1 = 32'd10217
; 
32'd143497: dataIn1 = 32'd2224
; 
32'd143498: dataIn1 = 32'd3668
; 
32'd143499: dataIn1 = 32'd3670
; 
32'd143500: dataIn1 = 32'd9499
; 
32'd143501: dataIn1 = 32'd9500
; 
32'd143502: dataIn1 = 32'd9504
; 
32'd143503: dataIn1 = 32'd9506
; 
32'd143504: dataIn1 = 32'd9916
; 
32'd143505: dataIn1 = 32'd3669
; 
32'd143506: dataIn1 = 32'd9911
; 
32'd143507: dataIn1 = 32'd9913
; 
32'd143508: dataIn1 = 32'd9914
; 
32'd143509: dataIn1 = 32'd9919
; 
32'd143510: dataIn1 = 32'd10117
; 
32'd143511: dataIn1 = 32'd10174
; 
32'd143512: dataIn1 = 32'd2195
; 
32'd143513: dataIn1 = 32'd2224
; 
32'd143514: dataIn1 = 32'd2225
; 
32'd143515: dataIn1 = 32'd3668
; 
32'd143516: dataIn1 = 32'd3670
; 
32'd143517: dataIn1 = 32'd3671
; 
32'd143518: dataIn1 = 32'd9506
; 
32'd143519: dataIn1 = 32'd2225
; 
32'd143520: dataIn1 = 32'd3670
; 
32'd143521: dataIn1 = 32'd3671
; 
32'd143522: dataIn1 = 32'd9505
; 
32'd143523: dataIn1 = 32'd9506
; 
32'd143524: dataIn1 = 32'd9511
; 
32'd143525: dataIn1 = 32'd9512
; 
32'd143526: dataIn1 = 32'd9939
; 
32'd143527: dataIn1 = 32'd2225
; 
32'd143528: dataIn1 = 32'd3672
; 
32'd143529: dataIn1 = 32'd3675
; 
32'd143530: dataIn1 = 32'd3676
; 
32'd143531: dataIn1 = 32'd10175
; 
32'd143532: dataIn1 = 32'd10176
; 
32'd143533: dataIn1 = 32'd10231
; 
32'd143534: dataIn1 = 32'd2225
; 
32'd143535: dataIn1 = 32'd3673
; 
32'd143536: dataIn1 = 32'd9507
; 
32'd143537: dataIn1 = 32'd9509
; 
32'd143538: dataIn1 = 32'd9510
; 
32'd143539: dataIn1 = 32'd9512
; 
32'd143540: dataIn1 = 32'd9925
; 
32'd143541: dataIn1 = 32'd9935
; 
32'd143542: dataIn1 = 32'd10176
; 
32'd143543: dataIn1 = 32'd3674
; 
32'd143544: dataIn1 = 32'd9929
; 
32'd143545: dataIn1 = 32'd9930
; 
32'd143546: dataIn1 = 32'd9949
; 
32'd143547: dataIn1 = 32'd9950
; 
32'd143548: dataIn1 = 32'd10175
; 
32'd143549: dataIn1 = 32'd10181
; 
32'd143550: dataIn1 = 32'd59
; 
32'd143551: dataIn1 = 32'd2195
; 
32'd143552: dataIn1 = 32'd2225
; 
32'd143553: dataIn1 = 32'd3672
; 
32'd143554: dataIn1 = 32'd3675
; 
32'd143555: dataIn1 = 32'd3676
; 
32'd143556: dataIn1 = 32'd59
; 
32'd143557: dataIn1 = 32'd2227
; 
32'd143558: dataIn1 = 32'd3672
; 
32'd143559: dataIn1 = 32'd3675
; 
32'd143560: dataIn1 = 32'd3676
; 
32'd143561: dataIn1 = 32'd3680
; 
32'd143562: dataIn1 = 32'd3683
; 
32'd143563: dataIn1 = 32'd10231
; 
32'd143564: dataIn1 = 32'd3677
; 
32'd143565: dataIn1 = 32'd9931
; 
32'd143566: dataIn1 = 32'd9932
; 
32'd143567: dataIn1 = 32'd9938
; 
32'd143568: dataIn1 = 32'd9943
; 
32'd143569: dataIn1 = 32'd10177
; 
32'd143570: dataIn1 = 32'd10179
; 
32'd143571: dataIn1 = 32'd3678
; 
32'd143572: dataIn1 = 32'd9523
; 
32'd143573: dataIn1 = 32'd9947
; 
32'd143574: dataIn1 = 32'd9948
; 
32'd143575: dataIn1 = 32'd9953
; 
32'd143576: dataIn1 = 32'd9962
; 
32'd143577: dataIn1 = 32'd10182
; 
32'd143578: dataIn1 = 32'd3679
; 
32'd143579: dataIn1 = 32'd3782
; 
32'd143580: dataIn1 = 32'd3784
; 
32'd143581: dataIn1 = 32'd9515
; 
32'd143582: dataIn1 = 32'd9517
; 
32'd143583: dataIn1 = 32'd9518
; 
32'd143584: dataIn1 = 32'd9519
; 
32'd143585: dataIn1 = 32'd9945
; 
32'd143586: dataIn1 = 32'd2198
; 
32'd143587: dataIn1 = 32'd2227
; 
32'd143588: dataIn1 = 32'd3676
; 
32'd143589: dataIn1 = 32'd3680
; 
32'd143590: dataIn1 = 32'd3681
; 
32'd143591: dataIn1 = 32'd3682
; 
32'd143592: dataIn1 = 32'd3683
; 
32'd143593: dataIn1 = 32'd10233
; 
32'd143594: dataIn1 = 32'd3680
; 
32'd143595: dataIn1 = 32'd3681
; 
32'd143596: dataIn1 = 32'd3682
; 
32'd143597: dataIn1 = 32'd9521
; 
32'd143598: dataIn1 = 32'd9523
; 
32'd143599: dataIn1 = 32'd9525
; 
32'd143600: dataIn1 = 32'd10233
; 
32'd143601: dataIn1 = 32'd2198
; 
32'd143602: dataIn1 = 32'd2228
; 
32'd143603: dataIn1 = 32'd3680
; 
32'd143604: dataIn1 = 32'd3681
; 
32'd143605: dataIn1 = 32'd3682
; 
32'd143606: dataIn1 = 32'd3685
; 
32'd143607: dataIn1 = 32'd3686
; 
32'd143608: dataIn1 = 32'd9525
; 
32'd143609: dataIn1 = 32'd59
; 
32'd143610: dataIn1 = 32'd2197
; 
32'd143611: dataIn1 = 32'd2198
; 
32'd143612: dataIn1 = 32'd3676
; 
32'd143613: dataIn1 = 32'd3680
; 
32'd143614: dataIn1 = 32'd3683
; 
32'd143615: dataIn1 = 32'd3684
; 
32'd143616: dataIn1 = 32'd9954
; 
32'd143617: dataIn1 = 32'd9955
; 
32'd143618: dataIn1 = 32'd9957
; 
32'd143619: dataIn1 = 32'd9963
; 
32'd143620: dataIn1 = 32'd9982
; 
32'd143621: dataIn1 = 32'd10184
; 
32'd143622: dataIn1 = 32'd60
; 
32'd143623: dataIn1 = 32'd2198
; 
32'd143624: dataIn1 = 32'd2199
; 
32'd143625: dataIn1 = 32'd3682
; 
32'd143626: dataIn1 = 32'd3685
; 
32'd143627: dataIn1 = 32'd3686
; 
32'd143628: dataIn1 = 32'd60
; 
32'd143629: dataIn1 = 32'd2228
; 
32'd143630: dataIn1 = 32'd3682
; 
32'd143631: dataIn1 = 32'd3685
; 
32'd143632: dataIn1 = 32'd3686
; 
32'd143633: dataIn1 = 32'd3687
; 
32'd143634: dataIn1 = 32'd3690
; 
32'd143635: dataIn1 = 32'd9533
; 
32'd143636: dataIn1 = 32'd10188
; 
32'd143637: dataIn1 = 32'd3686
; 
32'd143638: dataIn1 = 32'd3687
; 
32'd143639: dataIn1 = 32'd9533
; 
32'd143640: dataIn1 = 32'd9967
; 
32'd143641: dataIn1 = 32'd9968
; 
32'd143642: dataIn1 = 32'd9974
; 
32'd143643: dataIn1 = 32'd10188
; 
32'd143644: dataIn1 = 32'd3688
; 
32'd143645: dataIn1 = 32'd9969
; 
32'd143646: dataIn1 = 32'd9970
; 
32'd143647: dataIn1 = 32'd9978
; 
32'd143648: dataIn1 = 32'd9983
; 
32'd143649: dataIn1 = 32'd10186
; 
32'd143650: dataIn1 = 32'd10189
; 
32'd143651: dataIn1 = 32'd3689
; 
32'd143652: dataIn1 = 32'd3693
; 
32'd143653: dataIn1 = 32'd9527
; 
32'd143654: dataIn1 = 32'd9528
; 
32'd143655: dataIn1 = 32'd9530
; 
32'd143656: dataIn1 = 32'd9535
; 
32'd143657: dataIn1 = 32'd9966
; 
32'd143658: dataIn1 = 32'd9973
; 
32'd143659: dataIn1 = 32'd10185
; 
32'd143660: dataIn1 = 32'd60
; 
32'd143661: dataIn1 = 32'd3615
; 
32'd143662: dataIn1 = 32'd3686
; 
32'd143663: dataIn1 = 32'd3690
; 
32'd143664: dataIn1 = 32'd10187
; 
32'd143665: dataIn1 = 32'd10188
; 
32'd143666: dataIn1 = 32'd10192
; 
32'd143667: dataIn1 = 32'd3691
; 
32'd143668: dataIn1 = 32'd3788
; 
32'd143669: dataIn1 = 32'd3792
; 
32'd143670: dataIn1 = 32'd10183
; 
32'd143671: dataIn1 = 32'd10184
; 
32'd143672: dataIn1 = 32'd10189
; 
32'd143673: dataIn1 = 32'd10234
; 
32'd143674: dataIn1 = 32'd71
; 
32'd143675: dataIn1 = 32'd3692
; 
32'd143676: dataIn1 = 32'd3693
; 
32'd143677: dataIn1 = 32'd9535
; 
32'd143678: dataIn1 = 32'd9536
; 
32'd143679: dataIn1 = 32'd9544
; 
32'd143680: dataIn1 = 32'd10235
; 
32'd143681: dataIn1 = 32'd71
; 
32'd143682: dataIn1 = 32'd2229
; 
32'd143683: dataIn1 = 32'd3689
; 
32'd143684: dataIn1 = 32'd3692
; 
32'd143685: dataIn1 = 32'd3693
; 
32'd143686: dataIn1 = 32'd3794
; 
32'd143687: dataIn1 = 32'd3796
; 
32'd143688: dataIn1 = 32'd9535
; 
32'd143689: dataIn1 = 32'd10185
; 
32'd143690: dataIn1 = 32'd2201
; 
32'd143691: dataIn1 = 32'd3615
; 
32'd143692: dataIn1 = 32'd3694
; 
32'd143693: dataIn1 = 32'd9538
; 
32'd143694: dataIn1 = 32'd9539
; 
32'd143695: dataIn1 = 32'd9543
; 
32'd143696: dataIn1 = 32'd9995
; 
32'd143697: dataIn1 = 32'd10192
; 
32'd143698: dataIn1 = 32'd3695
; 
32'd143699: dataIn1 = 32'd9544
; 
32'd143700: dataIn1 = 32'd9986
; 
32'd143701: dataIn1 = 32'd9988
; 
32'd143702: dataIn1 = 32'd9992
; 
32'd143703: dataIn1 = 32'd9998
; 
32'd143704: dataIn1 = 32'd10190
; 
32'd143705: dataIn1 = 32'd2201
; 
32'd143706: dataIn1 = 32'd3696
; 
32'd143707: dataIn1 = 32'd9538
; 
32'd143708: dataIn1 = 32'd9546
; 
32'd143709: dataIn1 = 32'd9993
; 
32'd143710: dataIn1 = 32'd9994
; 
32'd143711: dataIn1 = 32'd10009
; 
32'd143712: dataIn1 = 32'd71
; 
32'd143713: dataIn1 = 32'd3697
; 
32'd143714: dataIn1 = 32'd3700
; 
32'd143715: dataIn1 = 32'd3703
; 
32'd143716: dataIn1 = 32'd10190
; 
32'd143717: dataIn1 = 32'd10191
; 
32'd143718: dataIn1 = 32'd10235
; 
32'd143719: dataIn1 = 32'd3698
; 
32'd143720: dataIn1 = 32'd10002
; 
32'd143721: dataIn1 = 32'd10004
; 
32'd143722: dataIn1 = 32'd10008
; 
32'd143723: dataIn1 = 32'd10011
; 
32'd143724: dataIn1 = 32'd10015
; 
32'd143725: dataIn1 = 32'd10194
; 
32'd143726: dataIn1 = 32'd2233
; 
32'd143727: dataIn1 = 32'd3699
; 
32'd143728: dataIn1 = 32'd3700
; 
32'd143729: dataIn1 = 32'd3701
; 
32'd143730: dataIn1 = 32'd10193
; 
32'd143731: dataIn1 = 32'd10194
; 
32'd143732: dataIn1 = 32'd10195
; 
32'd143733: dataIn1 = 32'd2231
; 
32'd143734: dataIn1 = 32'd2232
; 
32'd143735: dataIn1 = 32'd3697
; 
32'd143736: dataIn1 = 32'd3699
; 
32'd143737: dataIn1 = 32'd3700
; 
32'd143738: dataIn1 = 32'd3701
; 
32'd143739: dataIn1 = 32'd3703
; 
32'd143740: dataIn1 = 32'd10191
; 
32'd143741: dataIn1 = 32'd10193
; 
32'd143742: dataIn1 = 32'd2232
; 
32'd143743: dataIn1 = 32'd2233
; 
32'd143744: dataIn1 = 32'd3699
; 
32'd143745: dataIn1 = 32'd3700
; 
32'd143746: dataIn1 = 32'd3701
; 
32'd143747: dataIn1 = 32'd3704
; 
32'd143748: dataIn1 = 32'd3705
; 
32'd143749: dataIn1 = 32'd2233
; 
32'd143750: dataIn1 = 32'd3702
; 
32'd143751: dataIn1 = 32'd9555
; 
32'd143752: dataIn1 = 32'd10016
; 
32'd143753: dataIn1 = 32'd10017
; 
32'd143754: dataIn1 = 32'd10024
; 
32'd143755: dataIn1 = 32'd10195
; 
32'd143756: dataIn1 = 32'd71
; 
32'd143757: dataIn1 = 32'd2232
; 
32'd143758: dataIn1 = 32'd3697
; 
32'd143759: dataIn1 = 32'd3700
; 
32'd143760: dataIn1 = 32'd3703
; 
32'd143761: dataIn1 = 32'd3800
; 
32'd143762: dataIn1 = 32'd3804
; 
32'd143763: dataIn1 = 32'd72
; 
32'd143764: dataIn1 = 32'd2233
; 
32'd143765: dataIn1 = 32'd3701
; 
32'd143766: dataIn1 = 32'd3704
; 
32'd143767: dataIn1 = 32'd3705
; 
32'd143768: dataIn1 = 32'd3707
; 
32'd143769: dataIn1 = 32'd3709
; 
32'd143770: dataIn1 = 32'd72
; 
32'd143771: dataIn1 = 32'd2232
; 
32'd143772: dataIn1 = 32'd3701
; 
32'd143773: dataIn1 = 32'd3704
; 
32'd143774: dataIn1 = 32'd3705
; 
32'd143775: dataIn1 = 32'd3806
; 
32'd143776: dataIn1 = 32'd3808
; 
32'd143777: dataIn1 = 32'd2233
; 
32'd143778: dataIn1 = 32'd3706
; 
32'd143779: dataIn1 = 32'd3707
; 
32'd143780: dataIn1 = 32'd3708
; 
32'd143781: dataIn1 = 32'd9554
; 
32'd143782: dataIn1 = 32'd9555
; 
32'd143783: dataIn1 = 32'd9557
; 
32'd143784: dataIn1 = 32'd2233
; 
32'd143785: dataIn1 = 32'd2234
; 
32'd143786: dataIn1 = 32'd3704
; 
32'd143787: dataIn1 = 32'd3706
; 
32'd143788: dataIn1 = 32'd3707
; 
32'd143789: dataIn1 = 32'd3708
; 
32'd143790: dataIn1 = 32'd3709
; 
32'd143791: dataIn1 = 32'd2204
; 
32'd143792: dataIn1 = 32'd2234
; 
32'd143793: dataIn1 = 32'd3627
; 
32'd143794: dataIn1 = 32'd3706
; 
32'd143795: dataIn1 = 32'd3707
; 
32'd143796: dataIn1 = 32'd3708
; 
32'd143797: dataIn1 = 32'd3710
; 
32'd143798: dataIn1 = 32'd9557
; 
32'd143799: dataIn1 = 32'd10163
; 
32'd143800: dataIn1 = 32'd72
; 
32'd143801: dataIn1 = 32'd2234
; 
32'd143802: dataIn1 = 32'd3704
; 
32'd143803: dataIn1 = 32'd3707
; 
32'd143804: dataIn1 = 32'd3709
; 
32'd143805: dataIn1 = 32'd3712
; 
32'd143806: dataIn1 = 32'd3715
; 
32'd143807: dataIn1 = 32'd62
; 
32'd143808: dataIn1 = 32'd2234
; 
32'd143809: dataIn1 = 32'd3627
; 
32'd143810: dataIn1 = 32'd3708
; 
32'd143811: dataIn1 = 32'd3710
; 
32'd143812: dataIn1 = 32'd3711
; 
32'd143813: dataIn1 = 32'd3714
; 
32'd143814: dataIn1 = 32'd2234
; 
32'd143815: dataIn1 = 32'd2236
; 
32'd143816: dataIn1 = 32'd3710
; 
32'd143817: dataIn1 = 32'd3711
; 
32'd143818: dataIn1 = 32'd3712
; 
32'd143819: dataIn1 = 32'd3713
; 
32'd143820: dataIn1 = 32'd3714
; 
32'd143821: dataIn1 = 32'd2234
; 
32'd143822: dataIn1 = 32'd2235
; 
32'd143823: dataIn1 = 32'd3709
; 
32'd143824: dataIn1 = 32'd3711
; 
32'd143825: dataIn1 = 32'd3712
; 
32'd143826: dataIn1 = 32'd3713
; 
32'd143827: dataIn1 = 32'd3715
; 
32'd143828: dataIn1 = 32'd2235
; 
32'd143829: dataIn1 = 32'd2236
; 
32'd143830: dataIn1 = 32'd3711
; 
32'd143831: dataIn1 = 32'd3712
; 
32'd143832: dataIn1 = 32'd3713
; 
32'd143833: dataIn1 = 32'd3716
; 
32'd143834: dataIn1 = 32'd3717
; 
32'd143835: dataIn1 = 32'd62
; 
32'd143836: dataIn1 = 32'd2236
; 
32'd143837: dataIn1 = 32'd3638
; 
32'd143838: dataIn1 = 32'd3710
; 
32'd143839: dataIn1 = 32'd3711
; 
32'd143840: dataIn1 = 32'd3714
; 
32'd143841: dataIn1 = 32'd3718
; 
32'd143842: dataIn1 = 32'd72
; 
32'd143843: dataIn1 = 32'd2235
; 
32'd143844: dataIn1 = 32'd3709
; 
32'd143845: dataIn1 = 32'd3712
; 
32'd143846: dataIn1 = 32'd3715
; 
32'd143847: dataIn1 = 32'd3812
; 
32'd143848: dataIn1 = 32'd3816
; 
32'd143849: dataIn1 = 32'd73
; 
32'd143850: dataIn1 = 32'd2236
; 
32'd143851: dataIn1 = 32'd3713
; 
32'd143852: dataIn1 = 32'd3716
; 
32'd143853: dataIn1 = 32'd3717
; 
32'd143854: dataIn1 = 32'd3719
; 
32'd143855: dataIn1 = 32'd3721
; 
32'd143856: dataIn1 = 32'd73
; 
32'd143857: dataIn1 = 32'd2235
; 
32'd143858: dataIn1 = 32'd3713
; 
32'd143859: dataIn1 = 32'd3716
; 
32'd143860: dataIn1 = 32'd3717
; 
32'd143861: dataIn1 = 32'd3818
; 
32'd143862: dataIn1 = 32'd3820
; 
32'd143863: dataIn1 = 32'd2207
; 
32'd143864: dataIn1 = 32'd2236
; 
32'd143865: dataIn1 = 32'd3638
; 
32'd143866: dataIn1 = 32'd3714
; 
32'd143867: dataIn1 = 32'd3718
; 
32'd143868: dataIn1 = 32'd3719
; 
32'd143869: dataIn1 = 32'd3720
; 
32'd143870: dataIn1 = 32'd2236
; 
32'd143871: dataIn1 = 32'd2237
; 
32'd143872: dataIn1 = 32'd3716
; 
32'd143873: dataIn1 = 32'd3718
; 
32'd143874: dataIn1 = 32'd3719
; 
32'd143875: dataIn1 = 32'd3720
; 
32'd143876: dataIn1 = 32'd3721
; 
32'd143877: dataIn1 = 32'd2207
; 
32'd143878: dataIn1 = 32'd2237
; 
32'd143879: dataIn1 = 32'd3640
; 
32'd143880: dataIn1 = 32'd3718
; 
32'd143881: dataIn1 = 32'd3719
; 
32'd143882: dataIn1 = 32'd3720
; 
32'd143883: dataIn1 = 32'd3722
; 
32'd143884: dataIn1 = 32'd73
; 
32'd143885: dataIn1 = 32'd2237
; 
32'd143886: dataIn1 = 32'd3716
; 
32'd143887: dataIn1 = 32'd3719
; 
32'd143888: dataIn1 = 32'd3721
; 
32'd143889: dataIn1 = 32'd3724
; 
32'd143890: dataIn1 = 32'd3727
; 
32'd143891: dataIn1 = 32'd63
; 
32'd143892: dataIn1 = 32'd2237
; 
32'd143893: dataIn1 = 32'd3640
; 
32'd143894: dataIn1 = 32'd3720
; 
32'd143895: dataIn1 = 32'd3722
; 
32'd143896: dataIn1 = 32'd3723
; 
32'd143897: dataIn1 = 32'd3726
; 
32'd143898: dataIn1 = 32'd2237
; 
32'd143899: dataIn1 = 32'd2239
; 
32'd143900: dataIn1 = 32'd3722
; 
32'd143901: dataIn1 = 32'd3723
; 
32'd143902: dataIn1 = 32'd3724
; 
32'd143903: dataIn1 = 32'd3725
; 
32'd143904: dataIn1 = 32'd3726
; 
32'd143905: dataIn1 = 32'd2237
; 
32'd143906: dataIn1 = 32'd2238
; 
32'd143907: dataIn1 = 32'd3721
; 
32'd143908: dataIn1 = 32'd3723
; 
32'd143909: dataIn1 = 32'd3724
; 
32'd143910: dataIn1 = 32'd3725
; 
32'd143911: dataIn1 = 32'd3727
; 
32'd143912: dataIn1 = 32'd74
; 
32'd143913: dataIn1 = 32'd2238
; 
32'd143914: dataIn1 = 32'd2239
; 
32'd143915: dataIn1 = 32'd3723
; 
32'd143916: dataIn1 = 32'd3724
; 
32'd143917: dataIn1 = 32'd3725
; 
32'd143918: dataIn1 = 32'd63
; 
32'd143919: dataIn1 = 32'd2239
; 
32'd143920: dataIn1 = 32'd3650
; 
32'd143921: dataIn1 = 32'd3722
; 
32'd143922: dataIn1 = 32'd3723
; 
32'd143923: dataIn1 = 32'd3726
; 
32'd143924: dataIn1 = 32'd3728
; 
32'd143925: dataIn1 = 32'd73
; 
32'd143926: dataIn1 = 32'd2238
; 
32'd143927: dataIn1 = 32'd2264
; 
32'd143928: dataIn1 = 32'd3721
; 
32'd143929: dataIn1 = 32'd3724
; 
32'd143930: dataIn1 = 32'd3727
; 
32'd143931: dataIn1 = 32'd2210
; 
32'd143932: dataIn1 = 32'd2239
; 
32'd143933: dataIn1 = 32'd3650
; 
32'd143934: dataIn1 = 32'd3726
; 
32'd143935: dataIn1 = 32'd3728
; 
32'd143936: dataIn1 = 32'd3729
; 
32'd143937: dataIn1 = 32'd3730
; 
32'd143938: dataIn1 = 32'd74
; 
32'd143939: dataIn1 = 32'd2239
; 
32'd143940: dataIn1 = 32'd2240
; 
32'd143941: dataIn1 = 32'd3728
; 
32'd143942: dataIn1 = 32'd3729
; 
32'd143943: dataIn1 = 32'd3730
; 
32'd143944: dataIn1 = 32'd2210
; 
32'd143945: dataIn1 = 32'd2240
; 
32'd143946: dataIn1 = 32'd3652
; 
32'd143947: dataIn1 = 32'd3728
; 
32'd143948: dataIn1 = 32'd3729
; 
32'd143949: dataIn1 = 32'd3730
; 
32'd143950: dataIn1 = 32'd3731
; 
32'd143951: dataIn1 = 32'd64
; 
32'd143952: dataIn1 = 32'd2240
; 
32'd143953: dataIn1 = 32'd3652
; 
32'd143954: dataIn1 = 32'd3730
; 
32'd143955: dataIn1 = 32'd3731
; 
32'd143956: dataIn1 = 32'd5312
; 
32'd143957: dataIn1 = 32'd2243
; 
32'd143958: dataIn1 = 32'd3732
; 
32'd143959: dataIn1 = 32'd3733
; 
32'd143960: dataIn1 = 32'd10197
; 
32'd143961: dataIn1 = 32'd10198
; 
32'd143962: dataIn1 = 32'd10236
; 
32'd143963: dataIn1 = 32'd2241
; 
32'd143964: dataIn1 = 32'd2243
; 
32'd143965: dataIn1 = 32'd3732
; 
32'd143966: dataIn1 = 32'd3733
; 
32'd143967: dataIn1 = 32'd3734
; 
32'd143968: dataIn1 = 32'd3737
; 
32'd143969: dataIn1 = 32'd3738
; 
32'd143970: dataIn1 = 32'd10236
; 
32'd143971: dataIn1 = 32'd2241
; 
32'd143972: dataIn1 = 32'd2242
; 
32'd143973: dataIn1 = 32'd3733
; 
32'd143974: dataIn1 = 32'd3734
; 
32'd143975: dataIn1 = 32'd3739
; 
32'd143976: dataIn1 = 32'd3740
; 
32'd143977: dataIn1 = 32'd10236
; 
32'd143978: dataIn1 = 32'd3735
; 
32'd143979: dataIn1 = 32'd10030
; 
32'd143980: dataIn1 = 32'd10031
; 
32'd143981: dataIn1 = 32'd10287
; 
32'd143982: dataIn1 = 32'd3736
; 
32'd143983: dataIn1 = 32'd10032
; 
32'd143984: dataIn1 = 32'd10033
; 
32'd143985: dataIn1 = 32'd10046
; 
32'd143986: dataIn1 = 32'd10047
; 
32'd143987: dataIn1 = 32'd10197
; 
32'd143988: dataIn1 = 32'd10201
; 
32'd143989: dataIn1 = 32'd76
; 
32'd143990: dataIn1 = 32'd2243
; 
32'd143991: dataIn1 = 32'd3733
; 
32'd143992: dataIn1 = 32'd3737
; 
32'd143993: dataIn1 = 32'd3738
; 
32'd143994: dataIn1 = 32'd76
; 
32'd143995: dataIn1 = 32'd2241
; 
32'd143996: dataIn1 = 32'd3733
; 
32'd143997: dataIn1 = 32'd3737
; 
32'd143998: dataIn1 = 32'd3738
; 
32'd143999: dataIn1 = 32'd3821
; 
32'd144000: dataIn1 = 32'd3824
; 
32'd144001: dataIn1 = 32'd77
; 
32'd144002: dataIn1 = 32'd2242
; 
32'd144003: dataIn1 = 32'd3734
; 
32'd144004: dataIn1 = 32'd3739
; 
32'd144005: dataIn1 = 32'd3740
; 
32'd144006: dataIn1 = 32'd3742
; 
32'd144007: dataIn1 = 32'd3745
; 
32'd144008: dataIn1 = 32'd10237
; 
32'd144009: dataIn1 = 32'd77
; 
32'd144010: dataIn1 = 32'd2241
; 
32'd144011: dataIn1 = 32'd3734
; 
32'd144012: dataIn1 = 32'd3739
; 
32'd144013: dataIn1 = 32'd3740
; 
32'd144014: dataIn1 = 32'd3823
; 
32'd144015: dataIn1 = 32'd3825
; 
32'd144016: dataIn1 = 32'd3741
; 
32'd144017: dataIn1 = 32'd10037
; 
32'd144018: dataIn1 = 32'd10038
; 
32'd144019: dataIn1 = 32'd10044
; 
32'd144020: dataIn1 = 32'd10045
; 
32'd144021: dataIn1 = 32'd10200
; 
32'd144022: dataIn1 = 32'd10202
; 
32'd144023: dataIn1 = 32'd2244
; 
32'd144024: dataIn1 = 32'd3739
; 
32'd144025: dataIn1 = 32'd3742
; 
32'd144026: dataIn1 = 32'd3745
; 
32'd144027: dataIn1 = 32'd10199
; 
32'd144028: dataIn1 = 32'd10200
; 
32'd144029: dataIn1 = 32'd10237
; 
32'd144030: dataIn1 = 32'd2244
; 
32'd144031: dataIn1 = 32'd3743
; 
32'd144032: dataIn1 = 32'd9561
; 
32'd144033: dataIn1 = 32'd9562
; 
32'd144034: dataIn1 = 32'd9569
; 
32'd144035: dataIn1 = 32'd9570
; 
32'd144036: dataIn1 = 32'd10036
; 
32'd144037: dataIn1 = 32'd10055
; 
32'd144038: dataIn1 = 32'd10199
; 
32'd144039: dataIn1 = 32'd3658
; 
32'd144040: dataIn1 = 32'd3744
; 
32'd144041: dataIn1 = 32'd5310
; 
32'd144042: dataIn1 = 32'd9564
; 
32'd144043: dataIn1 = 32'd9565
; 
32'd144044: dataIn1 = 32'd9567
; 
32'd144045: dataIn1 = 32'd9568
; 
32'd144046: dataIn1 = 32'd10043
; 
32'd144047: dataIn1 = 32'd77
; 
32'd144048: dataIn1 = 32'd2244
; 
32'd144049: dataIn1 = 32'd3739
; 
32'd144050: dataIn1 = 32'd3742
; 
32'd144051: dataIn1 = 32'd3745
; 
32'd144052: dataIn1 = 32'd3749
; 
32'd144053: dataIn1 = 32'd3752
; 
32'd144054: dataIn1 = 32'd3746
; 
32'd144055: dataIn1 = 32'd10051
; 
32'd144056: dataIn1 = 32'd10052
; 
32'd144057: dataIn1 = 32'd10056
; 
32'd144058: dataIn1 = 32'd10061
; 
32'd144059: dataIn1 = 32'd10203
; 
32'd144060: dataIn1 = 32'd10206
; 
32'd144061: dataIn1 = 32'd2244
; 
32'd144062: dataIn1 = 32'd3747
; 
32'd144063: dataIn1 = 32'd3748
; 
32'd144064: dataIn1 = 32'd9569
; 
32'd144065: dataIn1 = 32'd9571
; 
32'd144066: dataIn1 = 32'd9573
; 
32'd144067: dataIn1 = 32'd9575
; 
32'd144068: dataIn1 = 32'd10059
; 
32'd144069: dataIn1 = 32'd2244
; 
32'd144070: dataIn1 = 32'd2246
; 
32'd144071: dataIn1 = 32'd3747
; 
32'd144072: dataIn1 = 32'd3748
; 
32'd144073: dataIn1 = 32'd3749
; 
32'd144074: dataIn1 = 32'd3750
; 
32'd144075: dataIn1 = 32'd3751
; 
32'd144076: dataIn1 = 32'd9575
; 
32'd144077: dataIn1 = 32'd2244
; 
32'd144078: dataIn1 = 32'd2245
; 
32'd144079: dataIn1 = 32'd3745
; 
32'd144080: dataIn1 = 32'd3748
; 
32'd144081: dataIn1 = 32'd3749
; 
32'd144082: dataIn1 = 32'd3750
; 
32'd144083: dataIn1 = 32'd3752
; 
32'd144084: dataIn1 = 32'd2245
; 
32'd144085: dataIn1 = 32'd2246
; 
32'd144086: dataIn1 = 32'd3748
; 
32'd144087: dataIn1 = 32'd3749
; 
32'd144088: dataIn1 = 32'd3750
; 
32'd144089: dataIn1 = 32'd3753
; 
32'd144090: dataIn1 = 32'd3754
; 
32'd144091: dataIn1 = 32'd2246
; 
32'd144092: dataIn1 = 32'd3748
; 
32'd144093: dataIn1 = 32'd3751
; 
32'd144094: dataIn1 = 32'd9575
; 
32'd144095: dataIn1 = 32'd9576
; 
32'd144096: dataIn1 = 32'd9580
; 
32'd144097: dataIn1 = 32'd9582
; 
32'd144098: dataIn1 = 32'd10073
; 
32'd144099: dataIn1 = 32'd77
; 
32'd144100: dataIn1 = 32'd2245
; 
32'd144101: dataIn1 = 32'd3745
; 
32'd144102: dataIn1 = 32'd3749
; 
32'd144103: dataIn1 = 32'd3752
; 
32'd144104: dataIn1 = 32'd3827
; 
32'd144105: dataIn1 = 32'd3831
; 
32'd144106: dataIn1 = 32'd78
; 
32'd144107: dataIn1 = 32'd2246
; 
32'd144108: dataIn1 = 32'd3750
; 
32'd144109: dataIn1 = 32'd3753
; 
32'd144110: dataIn1 = 32'd3754
; 
32'd144111: dataIn1 = 32'd3756
; 
32'd144112: dataIn1 = 32'd3759
; 
32'd144113: dataIn1 = 32'd78
; 
32'd144114: dataIn1 = 32'd2245
; 
32'd144115: dataIn1 = 32'd3750
; 
32'd144116: dataIn1 = 32'd3753
; 
32'd144117: dataIn1 = 32'd3754
; 
32'd144118: dataIn1 = 32'd3833
; 
32'd144119: dataIn1 = 32'd3835
; 
32'd144120: dataIn1 = 32'd2246
; 
32'd144121: dataIn1 = 32'd3755
; 
32'd144122: dataIn1 = 32'd3756
; 
32'd144123: dataIn1 = 32'd9578
; 
32'd144124: dataIn1 = 32'd9579
; 
32'd144125: dataIn1 = 32'd9581
; 
32'd144126: dataIn1 = 32'd9582
; 
32'd144127: dataIn1 = 32'd10077
; 
32'd144128: dataIn1 = 32'd2246
; 
32'd144129: dataIn1 = 32'd2247
; 
32'd144130: dataIn1 = 32'd3753
; 
32'd144131: dataIn1 = 32'd3755
; 
32'd144132: dataIn1 = 32'd3756
; 
32'd144133: dataIn1 = 32'd3757
; 
32'd144134: dataIn1 = 32'd3759
; 
32'd144135: dataIn1 = 32'd9578
; 
32'd144136: dataIn1 = 32'd2247
; 
32'd144137: dataIn1 = 32'd3756
; 
32'd144138: dataIn1 = 32'd3757
; 
32'd144139: dataIn1 = 32'd9577
; 
32'd144140: dataIn1 = 32'd9578
; 
32'd144141: dataIn1 = 32'd9585
; 
32'd144142: dataIn1 = 32'd9586
; 
32'd144143: dataIn1 = 32'd10087
; 
32'd144144: dataIn1 = 32'd3758
; 
32'd144145: dataIn1 = 32'd10069
; 
32'd144146: dataIn1 = 32'd10070
; 
32'd144147: dataIn1 = 32'd10076
; 
32'd144148: dataIn1 = 32'd10081
; 
32'd144149: dataIn1 = 32'd10207
; 
32'd144150: dataIn1 = 32'd10209
; 
32'd144151: dataIn1 = 32'd78
; 
32'd144152: dataIn1 = 32'd2247
; 
32'd144153: dataIn1 = 32'd3753
; 
32'd144154: dataIn1 = 32'd3756
; 
32'd144155: dataIn1 = 32'd3759
; 
32'd144156: dataIn1 = 32'd3762
; 
32'd144157: dataIn1 = 32'd3765
; 
32'd144158: dataIn1 = 32'd2247
; 
32'd144159: dataIn1 = 32'd3760
; 
32'd144160: dataIn1 = 32'd3761
; 
32'd144161: dataIn1 = 32'd9585
; 
32'd144162: dataIn1 = 32'd9587
; 
32'd144163: dataIn1 = 32'd9589
; 
32'd144164: dataIn1 = 32'd9591
; 
32'd144165: dataIn1 = 32'd10091
; 
32'd144166: dataIn1 = 32'd2247
; 
32'd144167: dataIn1 = 32'd2249
; 
32'd144168: dataIn1 = 32'd3760
; 
32'd144169: dataIn1 = 32'd3761
; 
32'd144170: dataIn1 = 32'd3762
; 
32'd144171: dataIn1 = 32'd3763
; 
32'd144172: dataIn1 = 32'd3764
; 
32'd144173: dataIn1 = 32'd9591
; 
32'd144174: dataIn1 = 32'd2247
; 
32'd144175: dataIn1 = 32'd2248
; 
32'd144176: dataIn1 = 32'd3759
; 
32'd144177: dataIn1 = 32'd3761
; 
32'd144178: dataIn1 = 32'd3762
; 
32'd144179: dataIn1 = 32'd3763
; 
32'd144180: dataIn1 = 32'd3765
; 
32'd144181: dataIn1 = 32'd2248
; 
32'd144182: dataIn1 = 32'd2249
; 
32'd144183: dataIn1 = 32'd3761
; 
32'd144184: dataIn1 = 32'd3762
; 
32'd144185: dataIn1 = 32'd3763
; 
32'd144186: dataIn1 = 32'd3766
; 
32'd144187: dataIn1 = 32'd3767
; 
32'd144188: dataIn1 = 32'd2249
; 
32'd144189: dataIn1 = 32'd3761
; 
32'd144190: dataIn1 = 32'd3764
; 
32'd144191: dataIn1 = 32'd9591
; 
32'd144192: dataIn1 = 32'd9592
; 
32'd144193: dataIn1 = 32'd9596
; 
32'd144194: dataIn1 = 32'd9598
; 
32'd144195: dataIn1 = 32'd10105
; 
32'd144196: dataIn1 = 32'd78
; 
32'd144197: dataIn1 = 32'd2248
; 
32'd144198: dataIn1 = 32'd3759
; 
32'd144199: dataIn1 = 32'd3762
; 
32'd144200: dataIn1 = 32'd3765
; 
32'd144201: dataIn1 = 32'd3837
; 
32'd144202: dataIn1 = 32'd3843
; 
32'd144203: dataIn1 = 32'd79
; 
32'd144204: dataIn1 = 32'd2249
; 
32'd144205: dataIn1 = 32'd3763
; 
32'd144206: dataIn1 = 32'd3766
; 
32'd144207: dataIn1 = 32'd3767
; 
32'd144208: dataIn1 = 32'd3769
; 
32'd144209: dataIn1 = 32'd3771
; 
32'd144210: dataIn1 = 32'd79
; 
32'd144211: dataIn1 = 32'd2248
; 
32'd144212: dataIn1 = 32'd3763
; 
32'd144213: dataIn1 = 32'd3766
; 
32'd144214: dataIn1 = 32'd3767
; 
32'd144215: dataIn1 = 32'd3845
; 
32'd144216: dataIn1 = 32'd3847
; 
32'd144217: dataIn1 = 32'd2249
; 
32'd144218: dataIn1 = 32'd3768
; 
32'd144219: dataIn1 = 32'd3769
; 
32'd144220: dataIn1 = 32'd9594
; 
32'd144221: dataIn1 = 32'd9595
; 
32'd144222: dataIn1 = 32'd9597
; 
32'd144223: dataIn1 = 32'd9598
; 
32'd144224: dataIn1 = 32'd10109
; 
32'd144225: dataIn1 = 32'd2249
; 
32'd144226: dataIn1 = 32'd2250
; 
32'd144227: dataIn1 = 32'd3766
; 
32'd144228: dataIn1 = 32'd3768
; 
32'd144229: dataIn1 = 32'd3769
; 
32'd144230: dataIn1 = 32'd3770
; 
32'd144231: dataIn1 = 32'd3771
; 
32'd144232: dataIn1 = 32'd9594
; 
32'd144233: dataIn1 = 32'd2250
; 
32'd144234: dataIn1 = 32'd3769
; 
32'd144235: dataIn1 = 32'd3770
; 
32'd144236: dataIn1 = 32'd9593
; 
32'd144237: dataIn1 = 32'd9594
; 
32'd144238: dataIn1 = 32'd9601
; 
32'd144239: dataIn1 = 32'd10116
; 
32'd144240: dataIn1 = 32'd10219
; 
32'd144241: dataIn1 = 32'd79
; 
32'd144242: dataIn1 = 32'd2250
; 
32'd144243: dataIn1 = 32'd3766
; 
32'd144244: dataIn1 = 32'd3769
; 
32'd144245: dataIn1 = 32'd3771
; 
32'd144246: dataIn1 = 32'd3774
; 
32'd144247: dataIn1 = 32'd3777
; 
32'd144248: dataIn1 = 32'd2250
; 
32'd144249: dataIn1 = 32'd3772
; 
32'd144250: dataIn1 = 32'd3773
; 
32'd144251: dataIn1 = 32'd10173
; 
32'd144252: dataIn1 = 32'd10174
; 
32'd144253: dataIn1 = 32'd10219
; 
32'd144254: dataIn1 = 32'd10230
; 
32'd144255: dataIn1 = 32'd2250
; 
32'd144256: dataIn1 = 32'd2252
; 
32'd144257: dataIn1 = 32'd3772
; 
32'd144258: dataIn1 = 32'd3773
; 
32'd144259: dataIn1 = 32'd3774
; 
32'd144260: dataIn1 = 32'd3775
; 
32'd144261: dataIn1 = 32'd3776
; 
32'd144262: dataIn1 = 32'd10230
; 
32'd144263: dataIn1 = 32'd2250
; 
32'd144264: dataIn1 = 32'd2251
; 
32'd144265: dataIn1 = 32'd3771
; 
32'd144266: dataIn1 = 32'd3773
; 
32'd144267: dataIn1 = 32'd3774
; 
32'd144268: dataIn1 = 32'd3775
; 
32'd144269: dataIn1 = 32'd3777
; 
32'd144270: dataIn1 = 32'd2251
; 
32'd144271: dataIn1 = 32'd2252
; 
32'd144272: dataIn1 = 32'd3773
; 
32'd144273: dataIn1 = 32'd3774
; 
32'd144274: dataIn1 = 32'd3775
; 
32'd144275: dataIn1 = 32'd3778
; 
32'd144276: dataIn1 = 32'd3779
; 
32'd144277: dataIn1 = 32'd2252
; 
32'd144278: dataIn1 = 32'd3773
; 
32'd144279: dataIn1 = 32'd3776
; 
32'd144280: dataIn1 = 32'd10179
; 
32'd144281: dataIn1 = 32'd10180
; 
32'd144282: dataIn1 = 32'd10230
; 
32'd144283: dataIn1 = 32'd10232
; 
32'd144284: dataIn1 = 32'd79
; 
32'd144285: dataIn1 = 32'd2251
; 
32'd144286: dataIn1 = 32'd3771
; 
32'd144287: dataIn1 = 32'd3774
; 
32'd144288: dataIn1 = 32'd3777
; 
32'd144289: dataIn1 = 32'd3849
; 
32'd144290: dataIn1 = 32'd3850
; 
32'd144291: dataIn1 = 32'd80
; 
32'd144292: dataIn1 = 32'd2252
; 
32'd144293: dataIn1 = 32'd3775
; 
32'd144294: dataIn1 = 32'd3778
; 
32'd144295: dataIn1 = 32'd3779
; 
32'd144296: dataIn1 = 32'd3781
; 
32'd144297: dataIn1 = 32'd3783
; 
32'd144298: dataIn1 = 32'd80
; 
32'd144299: dataIn1 = 32'd2251
; 
32'd144300: dataIn1 = 32'd3775
; 
32'd144301: dataIn1 = 32'd3778
; 
32'd144302: dataIn1 = 32'd3779
; 
32'd144303: dataIn1 = 32'd3852
; 
32'd144304: dataIn1 = 32'd3853
; 
32'd144305: dataIn1 = 32'd2252
; 
32'd144306: dataIn1 = 32'd3780
; 
32'd144307: dataIn1 = 32'd3781
; 
32'd144308: dataIn1 = 32'd3782
; 
32'd144309: dataIn1 = 32'd10177
; 
32'd144310: dataIn1 = 32'd10178
; 
32'd144311: dataIn1 = 32'd10232
; 
32'd144312: dataIn1 = 32'd2252
; 
32'd144313: dataIn1 = 32'd2253
; 
32'd144314: dataIn1 = 32'd3778
; 
32'd144315: dataIn1 = 32'd3780
; 
32'd144316: dataIn1 = 32'd3781
; 
32'd144317: dataIn1 = 32'd3782
; 
32'd144318: dataIn1 = 32'd3783
; 
32'd144319: dataIn1 = 32'd2226
; 
32'd144320: dataIn1 = 32'd2253
; 
32'd144321: dataIn1 = 32'd3679
; 
32'd144322: dataIn1 = 32'd3780
; 
32'd144323: dataIn1 = 32'd3781
; 
32'd144324: dataIn1 = 32'd3782
; 
32'd144325: dataIn1 = 32'd3784
; 
32'd144326: dataIn1 = 32'd9518
; 
32'd144327: dataIn1 = 32'd10178
; 
32'd144328: dataIn1 = 32'd80
; 
32'd144329: dataIn1 = 32'd2253
; 
32'd144330: dataIn1 = 32'd3778
; 
32'd144331: dataIn1 = 32'd3781
; 
32'd144332: dataIn1 = 32'd3783
; 
32'd144333: dataIn1 = 32'd3786
; 
32'd144334: dataIn1 = 32'd3789
; 
32'd144335: dataIn1 = 32'd70
; 
32'd144336: dataIn1 = 32'd2253
; 
32'd144337: dataIn1 = 32'd3679
; 
32'd144338: dataIn1 = 32'd3782
; 
32'd144339: dataIn1 = 32'd3784
; 
32'd144340: dataIn1 = 32'd3785
; 
32'd144341: dataIn1 = 32'd3788
; 
32'd144342: dataIn1 = 32'd9519
; 
32'd144343: dataIn1 = 32'd2253
; 
32'd144344: dataIn1 = 32'd2255
; 
32'd144345: dataIn1 = 32'd3784
; 
32'd144346: dataIn1 = 32'd3785
; 
32'd144347: dataIn1 = 32'd3786
; 
32'd144348: dataIn1 = 32'd3787
; 
32'd144349: dataIn1 = 32'd3788
; 
32'd144350: dataIn1 = 32'd2253
; 
32'd144351: dataIn1 = 32'd2254
; 
32'd144352: dataIn1 = 32'd3783
; 
32'd144353: dataIn1 = 32'd3785
; 
32'd144354: dataIn1 = 32'd3786
; 
32'd144355: dataIn1 = 32'd3787
; 
32'd144356: dataIn1 = 32'd3789
; 
32'd144357: dataIn1 = 32'd2254
; 
32'd144358: dataIn1 = 32'd2255
; 
32'd144359: dataIn1 = 32'd3785
; 
32'd144360: dataIn1 = 32'd3786
; 
32'd144361: dataIn1 = 32'd3787
; 
32'd144362: dataIn1 = 32'd3790
; 
32'd144363: dataIn1 = 32'd3791
; 
32'd144364: dataIn1 = 32'd70
; 
32'd144365: dataIn1 = 32'd2255
; 
32'd144366: dataIn1 = 32'd3691
; 
32'd144367: dataIn1 = 32'd3784
; 
32'd144368: dataIn1 = 32'd3785
; 
32'd144369: dataIn1 = 32'd3788
; 
32'd144370: dataIn1 = 32'd3792
; 
32'd144371: dataIn1 = 32'd10183
; 
32'd144372: dataIn1 = 32'd80
; 
32'd144373: dataIn1 = 32'd2254
; 
32'd144374: dataIn1 = 32'd3783
; 
32'd144375: dataIn1 = 32'd3786
; 
32'd144376: dataIn1 = 32'd3789
; 
32'd144377: dataIn1 = 32'd3855
; 
32'd144378: dataIn1 = 32'd3856
; 
32'd144379: dataIn1 = 32'd81
; 
32'd144380: dataIn1 = 32'd2255
; 
32'd144381: dataIn1 = 32'd3787
; 
32'd144382: dataIn1 = 32'd3790
; 
32'd144383: dataIn1 = 32'd3791
; 
32'd144384: dataIn1 = 32'd3793
; 
32'd144385: dataIn1 = 32'd3795
; 
32'd144386: dataIn1 = 32'd81
; 
32'd144387: dataIn1 = 32'd2254
; 
32'd144388: dataIn1 = 32'd3787
; 
32'd144389: dataIn1 = 32'd3790
; 
32'd144390: dataIn1 = 32'd3791
; 
32'd144391: dataIn1 = 32'd3858
; 
32'd144392: dataIn1 = 32'd3859
; 
32'd144393: dataIn1 = 32'd2229
; 
32'd144394: dataIn1 = 32'd2255
; 
32'd144395: dataIn1 = 32'd3691
; 
32'd144396: dataIn1 = 32'd3788
; 
32'd144397: dataIn1 = 32'd3792
; 
32'd144398: dataIn1 = 32'd3793
; 
32'd144399: dataIn1 = 32'd3794
; 
32'd144400: dataIn1 = 32'd10234
; 
32'd144401: dataIn1 = 32'd2255
; 
32'd144402: dataIn1 = 32'd2256
; 
32'd144403: dataIn1 = 32'd3790
; 
32'd144404: dataIn1 = 32'd3792
; 
32'd144405: dataIn1 = 32'd3793
; 
32'd144406: dataIn1 = 32'd3794
; 
32'd144407: dataIn1 = 32'd3795
; 
32'd144408: dataIn1 = 32'd2229
; 
32'd144409: dataIn1 = 32'd2256
; 
32'd144410: dataIn1 = 32'd3693
; 
32'd144411: dataIn1 = 32'd3792
; 
32'd144412: dataIn1 = 32'd3793
; 
32'd144413: dataIn1 = 32'd3794
; 
32'd144414: dataIn1 = 32'd3796
; 
32'd144415: dataIn1 = 32'd81
; 
32'd144416: dataIn1 = 32'd2256
; 
32'd144417: dataIn1 = 32'd3790
; 
32'd144418: dataIn1 = 32'd3793
; 
32'd144419: dataIn1 = 32'd3795
; 
32'd144420: dataIn1 = 32'd3798
; 
32'd144421: dataIn1 = 32'd3801
; 
32'd144422: dataIn1 = 32'd71
; 
32'd144423: dataIn1 = 32'd2256
; 
32'd144424: dataIn1 = 32'd3693
; 
32'd144425: dataIn1 = 32'd3794
; 
32'd144426: dataIn1 = 32'd3796
; 
32'd144427: dataIn1 = 32'd3797
; 
32'd144428: dataIn1 = 32'd3800
; 
32'd144429: dataIn1 = 32'd2256
; 
32'd144430: dataIn1 = 32'd2258
; 
32'd144431: dataIn1 = 32'd3796
; 
32'd144432: dataIn1 = 32'd3797
; 
32'd144433: dataIn1 = 32'd3798
; 
32'd144434: dataIn1 = 32'd3799
; 
32'd144435: dataIn1 = 32'd3800
; 
32'd144436: dataIn1 = 32'd2256
; 
32'd144437: dataIn1 = 32'd2257
; 
32'd144438: dataIn1 = 32'd3795
; 
32'd144439: dataIn1 = 32'd3797
; 
32'd144440: dataIn1 = 32'd3798
; 
32'd144441: dataIn1 = 32'd3799
; 
32'd144442: dataIn1 = 32'd3801
; 
32'd144443: dataIn1 = 32'd2257
; 
32'd144444: dataIn1 = 32'd2258
; 
32'd144445: dataIn1 = 32'd3797
; 
32'd144446: dataIn1 = 32'd3798
; 
32'd144447: dataIn1 = 32'd3799
; 
32'd144448: dataIn1 = 32'd3802
; 
32'd144449: dataIn1 = 32'd3803
; 
32'd144450: dataIn1 = 32'd71
; 
32'd144451: dataIn1 = 32'd2258
; 
32'd144452: dataIn1 = 32'd3703
; 
32'd144453: dataIn1 = 32'd3796
; 
32'd144454: dataIn1 = 32'd3797
; 
32'd144455: dataIn1 = 32'd3800
; 
32'd144456: dataIn1 = 32'd3804
; 
32'd144457: dataIn1 = 32'd81
; 
32'd144458: dataIn1 = 32'd2257
; 
32'd144459: dataIn1 = 32'd3795
; 
32'd144460: dataIn1 = 32'd3798
; 
32'd144461: dataIn1 = 32'd3801
; 
32'd144462: dataIn1 = 32'd3861
; 
32'd144463: dataIn1 = 32'd3862
; 
32'd144464: dataIn1 = 32'd82
; 
32'd144465: dataIn1 = 32'd2258
; 
32'd144466: dataIn1 = 32'd3799
; 
32'd144467: dataIn1 = 32'd3802
; 
32'd144468: dataIn1 = 32'd3803
; 
32'd144469: dataIn1 = 32'd3805
; 
32'd144470: dataIn1 = 32'd3807
; 
32'd144471: dataIn1 = 32'd82
; 
32'd144472: dataIn1 = 32'd2257
; 
32'd144473: dataIn1 = 32'd2282
; 
32'd144474: dataIn1 = 32'd3799
; 
32'd144475: dataIn1 = 32'd3802
; 
32'd144476: dataIn1 = 32'd3803
; 
32'd144477: dataIn1 = 32'd2232
; 
32'd144478: dataIn1 = 32'd2258
; 
32'd144479: dataIn1 = 32'd3703
; 
32'd144480: dataIn1 = 32'd3800
; 
32'd144481: dataIn1 = 32'd3804
; 
32'd144482: dataIn1 = 32'd3805
; 
32'd144483: dataIn1 = 32'd3806
; 
32'd144484: dataIn1 = 32'd2258
; 
32'd144485: dataIn1 = 32'd2259
; 
32'd144486: dataIn1 = 32'd3802
; 
32'd144487: dataIn1 = 32'd3804
; 
32'd144488: dataIn1 = 32'd3805
; 
32'd144489: dataIn1 = 32'd3806
; 
32'd144490: dataIn1 = 32'd3807
; 
32'd144491: dataIn1 = 32'd2232
; 
32'd144492: dataIn1 = 32'd2259
; 
32'd144493: dataIn1 = 32'd3705
; 
32'd144494: dataIn1 = 32'd3804
; 
32'd144495: dataIn1 = 32'd3805
; 
32'd144496: dataIn1 = 32'd3806
; 
32'd144497: dataIn1 = 32'd3808
; 
32'd144498: dataIn1 = 32'd82
; 
32'd144499: dataIn1 = 32'd2259
; 
32'd144500: dataIn1 = 32'd3802
; 
32'd144501: dataIn1 = 32'd3805
; 
32'd144502: dataIn1 = 32'd3807
; 
32'd144503: dataIn1 = 32'd3810
; 
32'd144504: dataIn1 = 32'd3813
; 
32'd144505: dataIn1 = 32'd72
; 
32'd144506: dataIn1 = 32'd2259
; 
32'd144507: dataIn1 = 32'd3705
; 
32'd144508: dataIn1 = 32'd3806
; 
32'd144509: dataIn1 = 32'd3808
; 
32'd144510: dataIn1 = 32'd3809
; 
32'd144511: dataIn1 = 32'd3812
; 
32'd144512: dataIn1 = 32'd2259
; 
32'd144513: dataIn1 = 32'd2261
; 
32'd144514: dataIn1 = 32'd3808
; 
32'd144515: dataIn1 = 32'd3809
; 
32'd144516: dataIn1 = 32'd3810
; 
32'd144517: dataIn1 = 32'd3811
; 
32'd144518: dataIn1 = 32'd3812
; 
32'd144519: dataIn1 = 32'd2259
; 
32'd144520: dataIn1 = 32'd2260
; 
32'd144521: dataIn1 = 32'd3807
; 
32'd144522: dataIn1 = 32'd3809
; 
32'd144523: dataIn1 = 32'd3810
; 
32'd144524: dataIn1 = 32'd3811
; 
32'd144525: dataIn1 = 32'd3813
; 
32'd144526: dataIn1 = 32'd2260
; 
32'd144527: dataIn1 = 32'd2261
; 
32'd144528: dataIn1 = 32'd3809
; 
32'd144529: dataIn1 = 32'd3810
; 
32'd144530: dataIn1 = 32'd3811
; 
32'd144531: dataIn1 = 32'd3814
; 
32'd144532: dataIn1 = 32'd3815
; 
32'd144533: dataIn1 = 32'd72
; 
32'd144534: dataIn1 = 32'd2261
; 
32'd144535: dataIn1 = 32'd3715
; 
32'd144536: dataIn1 = 32'd3808
; 
32'd144537: dataIn1 = 32'd3809
; 
32'd144538: dataIn1 = 32'd3812
; 
32'd144539: dataIn1 = 32'd3816
; 
32'd144540: dataIn1 = 32'd82
; 
32'd144541: dataIn1 = 32'd2260
; 
32'd144542: dataIn1 = 32'd2284
; 
32'd144543: dataIn1 = 32'd3807
; 
32'd144544: dataIn1 = 32'd3810
; 
32'd144545: dataIn1 = 32'd3813
; 
32'd144546: dataIn1 = 32'd83
; 
32'd144547: dataIn1 = 32'd2261
; 
32'd144548: dataIn1 = 32'd3811
; 
32'd144549: dataIn1 = 32'd3814
; 
32'd144550: dataIn1 = 32'd3815
; 
32'd144551: dataIn1 = 32'd3817
; 
32'd144552: dataIn1 = 32'd3819
; 
32'd144553: dataIn1 = 32'd83
; 
32'd144554: dataIn1 = 32'd2260
; 
32'd144555: dataIn1 = 32'd2285
; 
32'd144556: dataIn1 = 32'd3811
; 
32'd144557: dataIn1 = 32'd3814
; 
32'd144558: dataIn1 = 32'd3815
; 
32'd144559: dataIn1 = 32'd2235
; 
32'd144560: dataIn1 = 32'd2261
; 
32'd144561: dataIn1 = 32'd3715
; 
32'd144562: dataIn1 = 32'd3812
; 
32'd144563: dataIn1 = 32'd3816
; 
32'd144564: dataIn1 = 32'd3817
; 
32'd144565: dataIn1 = 32'd3818
; 
32'd144566: dataIn1 = 32'd2261
; 
32'd144567: dataIn1 = 32'd2262
; 
32'd144568: dataIn1 = 32'd3814
; 
32'd144569: dataIn1 = 32'd3816
; 
32'd144570: dataIn1 = 32'd3817
; 
32'd144571: dataIn1 = 32'd3818
; 
32'd144572: dataIn1 = 32'd3819
; 
32'd144573: dataIn1 = 32'd2235
; 
32'd144574: dataIn1 = 32'd2262
; 
32'd144575: dataIn1 = 32'd3717
; 
32'd144576: dataIn1 = 32'd3816
; 
32'd144577: dataIn1 = 32'd3817
; 
32'd144578: dataIn1 = 32'd3818
; 
32'd144579: dataIn1 = 32'd3820
; 
32'd144580: dataIn1 = 32'd83
; 
32'd144581: dataIn1 = 32'd2262
; 
32'd144582: dataIn1 = 32'd2263
; 
32'd144583: dataIn1 = 32'd3814
; 
32'd144584: dataIn1 = 32'd3817
; 
32'd144585: dataIn1 = 32'd3819
; 
32'd144586: dataIn1 = 32'd73
; 
32'd144587: dataIn1 = 32'd2262
; 
32'd144588: dataIn1 = 32'd2264
; 
32'd144589: dataIn1 = 32'd3717
; 
32'd144590: dataIn1 = 32'd3818
; 
32'd144591: dataIn1 = 32'd3820
; 
32'd144592: dataIn1 = 32'd2241
; 
32'd144593: dataIn1 = 32'd2267
; 
32'd144594: dataIn1 = 32'd3738
; 
32'd144595: dataIn1 = 32'd3821
; 
32'd144596: dataIn1 = 32'd3822
; 
32'd144597: dataIn1 = 32'd3823
; 
32'd144598: dataIn1 = 32'd3824
; 
32'd144599: dataIn1 = 32'd87
; 
32'd144600: dataIn1 = 32'd2266
; 
32'd144601: dataIn1 = 32'd2267
; 
32'd144602: dataIn1 = 32'd3821
; 
32'd144603: dataIn1 = 32'd3822
; 
32'd144604: dataIn1 = 32'd3823
; 
32'd144605: dataIn1 = 32'd2241
; 
32'd144606: dataIn1 = 32'd2266
; 
32'd144607: dataIn1 = 32'd3740
; 
32'd144608: dataIn1 = 32'd3821
; 
32'd144609: dataIn1 = 32'd3822
; 
32'd144610: dataIn1 = 32'd3823
; 
32'd144611: dataIn1 = 32'd3825
; 
32'd144612: dataIn1 = 32'd76
; 
32'd144613: dataIn1 = 32'd2267
; 
32'd144614: dataIn1 = 32'd3738
; 
32'd144615: dataIn1 = 32'd3821
; 
32'd144616: dataIn1 = 32'd3824
; 
32'd144617: dataIn1 = 32'd77
; 
32'd144618: dataIn1 = 32'd2266
; 
32'd144619: dataIn1 = 32'd3740
; 
32'd144620: dataIn1 = 32'd3823
; 
32'd144621: dataIn1 = 32'd3825
; 
32'd144622: dataIn1 = 32'd3826
; 
32'd144623: dataIn1 = 32'd3827
; 
32'd144624: dataIn1 = 32'd2266
; 
32'd144625: dataIn1 = 32'd2269
; 
32'd144626: dataIn1 = 32'd3825
; 
32'd144627: dataIn1 = 32'd3826
; 
32'd144628: dataIn1 = 32'd3827
; 
32'd144629: dataIn1 = 32'd3830
; 
32'd144630: dataIn1 = 32'd5313
; 
32'd144631: dataIn1 = 32'd77
; 
32'd144632: dataIn1 = 32'd2269
; 
32'd144633: dataIn1 = 32'd3752
; 
32'd144634: dataIn1 = 32'd3825
; 
32'd144635: dataIn1 = 32'd3826
; 
32'd144636: dataIn1 = 32'd3827
; 
32'd144637: dataIn1 = 32'd3831
; 
32'd144638: dataIn1 = 32'd88
; 
32'd144639: dataIn1 = 32'd2269
; 
32'd144640: dataIn1 = 32'd3828
; 
32'd144641: dataIn1 = 32'd3829
; 
32'd144642: dataIn1 = 32'd3830
; 
32'd144643: dataIn1 = 32'd3832
; 
32'd144644: dataIn1 = 32'd3834
; 
32'd144645: dataIn1 = 32'd88
; 
32'd144646: dataIn1 = 32'd2268
; 
32'd144647: dataIn1 = 32'd3828
; 
32'd144648: dataIn1 = 32'd3829
; 
32'd144649: dataIn1 = 32'd3830
; 
32'd144650: dataIn1 = 32'd5314
; 
32'd144651: dataIn1 = 32'd2268
; 
32'd144652: dataIn1 = 32'd2269
; 
32'd144653: dataIn1 = 32'd3826
; 
32'd144654: dataIn1 = 32'd3828
; 
32'd144655: dataIn1 = 32'd3829
; 
32'd144656: dataIn1 = 32'd3830
; 
32'd144657: dataIn1 = 32'd5313
; 
32'd144658: dataIn1 = 32'd2245
; 
32'd144659: dataIn1 = 32'd2269
; 
32'd144660: dataIn1 = 32'd3752
; 
32'd144661: dataIn1 = 32'd3827
; 
32'd144662: dataIn1 = 32'd3831
; 
32'd144663: dataIn1 = 32'd3832
; 
32'd144664: dataIn1 = 32'd3833
; 
32'd144665: dataIn1 = 32'd2269
; 
32'd144666: dataIn1 = 32'd2270
; 
32'd144667: dataIn1 = 32'd3828
; 
32'd144668: dataIn1 = 32'd3831
; 
32'd144669: dataIn1 = 32'd3832
; 
32'd144670: dataIn1 = 32'd3833
; 
32'd144671: dataIn1 = 32'd3834
; 
32'd144672: dataIn1 = 32'd2245
; 
32'd144673: dataIn1 = 32'd2270
; 
32'd144674: dataIn1 = 32'd3754
; 
32'd144675: dataIn1 = 32'd3831
; 
32'd144676: dataIn1 = 32'd3832
; 
32'd144677: dataIn1 = 32'd3833
; 
32'd144678: dataIn1 = 32'd3835
; 
32'd144679: dataIn1 = 32'd88
; 
32'd144680: dataIn1 = 32'd2270
; 
32'd144681: dataIn1 = 32'd3828
; 
32'd144682: dataIn1 = 32'd3832
; 
32'd144683: dataIn1 = 32'd3834
; 
32'd144684: dataIn1 = 32'd3838
; 
32'd144685: dataIn1 = 32'd3839
; 
32'd144686: dataIn1 = 32'd78
; 
32'd144687: dataIn1 = 32'd2270
; 
32'd144688: dataIn1 = 32'd3754
; 
32'd144689: dataIn1 = 32'd3833
; 
32'd144690: dataIn1 = 32'd3835
; 
32'd144691: dataIn1 = 32'd3836
; 
32'd144692: dataIn1 = 32'd3837
; 
32'd144693: dataIn1 = 32'd2270
; 
32'd144694: dataIn1 = 32'd2272
; 
32'd144695: dataIn1 = 32'd3835
; 
32'd144696: dataIn1 = 32'd3836
; 
32'd144697: dataIn1 = 32'd3837
; 
32'd144698: dataIn1 = 32'd3838
; 
32'd144699: dataIn1 = 32'd3842
; 
32'd144700: dataIn1 = 32'd78
; 
32'd144701: dataIn1 = 32'd2272
; 
32'd144702: dataIn1 = 32'd3765
; 
32'd144703: dataIn1 = 32'd3835
; 
32'd144704: dataIn1 = 32'd3836
; 
32'd144705: dataIn1 = 32'd3837
; 
32'd144706: dataIn1 = 32'd3843
; 
32'd144707: dataIn1 = 32'd2270
; 
32'd144708: dataIn1 = 32'd2271
; 
32'd144709: dataIn1 = 32'd3834
; 
32'd144710: dataIn1 = 32'd3836
; 
32'd144711: dataIn1 = 32'd3838
; 
32'd144712: dataIn1 = 32'd3839
; 
32'd144713: dataIn1 = 32'd3842
; 
32'd144714: dataIn1 = 32'd88
; 
32'd144715: dataIn1 = 32'd2271
; 
32'd144716: dataIn1 = 32'd3834
; 
32'd144717: dataIn1 = 32'd3838
; 
32'd144718: dataIn1 = 32'd3839
; 
32'd144719: dataIn1 = 32'd5317
; 
32'd144720: dataIn1 = 32'd89
; 
32'd144721: dataIn1 = 32'd2272
; 
32'd144722: dataIn1 = 32'd3840
; 
32'd144723: dataIn1 = 32'd3841
; 
32'd144724: dataIn1 = 32'd3842
; 
32'd144725: dataIn1 = 32'd3844
; 
32'd144726: dataIn1 = 32'd3846
; 
32'd144727: dataIn1 = 32'd89
; 
32'd144728: dataIn1 = 32'd2271
; 
32'd144729: dataIn1 = 32'd3840
; 
32'd144730: dataIn1 = 32'd3841
; 
32'd144731: dataIn1 = 32'd3842
; 
32'd144732: dataIn1 = 32'd5316
; 
32'd144733: dataIn1 = 32'd2271
; 
32'd144734: dataIn1 = 32'd2272
; 
32'd144735: dataIn1 = 32'd3836
; 
32'd144736: dataIn1 = 32'd3838
; 
32'd144737: dataIn1 = 32'd3840
; 
32'd144738: dataIn1 = 32'd3841
; 
32'd144739: dataIn1 = 32'd3842
; 
32'd144740: dataIn1 = 32'd2248
; 
32'd144741: dataIn1 = 32'd2272
; 
32'd144742: dataIn1 = 32'd3765
; 
32'd144743: dataIn1 = 32'd3837
; 
32'd144744: dataIn1 = 32'd3843
; 
32'd144745: dataIn1 = 32'd3844
; 
32'd144746: dataIn1 = 32'd3845
; 
32'd144747: dataIn1 = 32'd2272
; 
32'd144748: dataIn1 = 32'd2273
; 
32'd144749: dataIn1 = 32'd3840
; 
32'd144750: dataIn1 = 32'd3843
; 
32'd144751: dataIn1 = 32'd3844
; 
32'd144752: dataIn1 = 32'd3845
; 
32'd144753: dataIn1 = 32'd3846
; 
32'd144754: dataIn1 = 32'd2248
; 
32'd144755: dataIn1 = 32'd2273
; 
32'd144756: dataIn1 = 32'd3767
; 
32'd144757: dataIn1 = 32'd3843
; 
32'd144758: dataIn1 = 32'd3844
; 
32'd144759: dataIn1 = 32'd3845
; 
32'd144760: dataIn1 = 32'd3847
; 
32'd144761: dataIn1 = 32'd89
; 
32'd144762: dataIn1 = 32'd2273
; 
32'd144763: dataIn1 = 32'd2274
; 
32'd144764: dataIn1 = 32'd3840
; 
32'd144765: dataIn1 = 32'd3844
; 
32'd144766: dataIn1 = 32'd3846
; 
32'd144767: dataIn1 = 32'd79
; 
32'd144768: dataIn1 = 32'd2273
; 
32'd144769: dataIn1 = 32'd3767
; 
32'd144770: dataIn1 = 32'd3845
; 
32'd144771: dataIn1 = 32'd3847
; 
32'd144772: dataIn1 = 32'd3848
; 
32'd144773: dataIn1 = 32'd3849
; 
32'd144774: dataIn1 = 32'd2273
; 
32'd144775: dataIn1 = 32'd2274
; 
32'd144776: dataIn1 = 32'd2275
; 
32'd144777: dataIn1 = 32'd3847
; 
32'd144778: dataIn1 = 32'd3848
; 
32'd144779: dataIn1 = 32'd3849
; 
32'd144780: dataIn1 = 32'd79
; 
32'd144781: dataIn1 = 32'd2275
; 
32'd144782: dataIn1 = 32'd3777
; 
32'd144783: dataIn1 = 32'd3847
; 
32'd144784: dataIn1 = 32'd3848
; 
32'd144785: dataIn1 = 32'd3849
; 
32'd144786: dataIn1 = 32'd3850
; 
32'd144787: dataIn1 = 32'd2251
; 
32'd144788: dataIn1 = 32'd2275
; 
32'd144789: dataIn1 = 32'd3777
; 
32'd144790: dataIn1 = 32'd3849
; 
32'd144791: dataIn1 = 32'd3850
; 
32'd144792: dataIn1 = 32'd3851
; 
32'd144793: dataIn1 = 32'd3852
; 
32'd144794: dataIn1 = 32'd90
; 
32'd144795: dataIn1 = 32'd2275
; 
32'd144796: dataIn1 = 32'd2276
; 
32'd144797: dataIn1 = 32'd3850
; 
32'd144798: dataIn1 = 32'd3851
; 
32'd144799: dataIn1 = 32'd3852
; 
32'd144800: dataIn1 = 32'd2251
; 
32'd144801: dataIn1 = 32'd2276
; 
32'd144802: dataIn1 = 32'd3779
; 
32'd144803: dataIn1 = 32'd3850
; 
32'd144804: dataIn1 = 32'd3851
; 
32'd144805: dataIn1 = 32'd3852
; 
32'd144806: dataIn1 = 32'd3853
; 
32'd144807: dataIn1 = 32'd80
; 
32'd144808: dataIn1 = 32'd2276
; 
32'd144809: dataIn1 = 32'd3779
; 
32'd144810: dataIn1 = 32'd3852
; 
32'd144811: dataIn1 = 32'd3853
; 
32'd144812: dataIn1 = 32'd3854
; 
32'd144813: dataIn1 = 32'd3855
; 
32'd144814: dataIn1 = 32'd2276
; 
32'd144815: dataIn1 = 32'd2277
; 
32'd144816: dataIn1 = 32'd2278
; 
32'd144817: dataIn1 = 32'd3853
; 
32'd144818: dataIn1 = 32'd3854
; 
32'd144819: dataIn1 = 32'd3855
; 
32'd144820: dataIn1 = 32'd80
; 
32'd144821: dataIn1 = 32'd2278
; 
32'd144822: dataIn1 = 32'd3789
; 
32'd144823: dataIn1 = 32'd3853
; 
32'd144824: dataIn1 = 32'd3854
; 
32'd144825: dataIn1 = 32'd3855
; 
32'd144826: dataIn1 = 32'd3856
; 
32'd144827: dataIn1 = 32'd2254
; 
32'd144828: dataIn1 = 32'd2278
; 
32'd144829: dataIn1 = 32'd3789
; 
32'd144830: dataIn1 = 32'd3855
; 
32'd144831: dataIn1 = 32'd3856
; 
32'd144832: dataIn1 = 32'd3857
; 
32'd144833: dataIn1 = 32'd3858
; 
32'd144834: dataIn1 = 32'd91
; 
32'd144835: dataIn1 = 32'd2278
; 
32'd144836: dataIn1 = 32'd2279
; 
32'd144837: dataIn1 = 32'd3856
; 
32'd144838: dataIn1 = 32'd3857
; 
32'd144839: dataIn1 = 32'd3858
; 
32'd144840: dataIn1 = 32'd2254
; 
32'd144841: dataIn1 = 32'd2279
; 
32'd144842: dataIn1 = 32'd3791
; 
32'd144843: dataIn1 = 32'd3856
; 
32'd144844: dataIn1 = 32'd3857
; 
32'd144845: dataIn1 = 32'd3858
; 
32'd144846: dataIn1 = 32'd3859
; 
32'd144847: dataIn1 = 32'd81
; 
32'd144848: dataIn1 = 32'd2279
; 
32'd144849: dataIn1 = 32'd3791
; 
32'd144850: dataIn1 = 32'd3858
; 
32'd144851: dataIn1 = 32'd3859
; 
32'd144852: dataIn1 = 32'd3860
; 
32'd144853: dataIn1 = 32'd3861
; 
32'd144854: dataIn1 = 32'd2279
; 
32'd144855: dataIn1 = 32'd2280
; 
32'd144856: dataIn1 = 32'd2281
; 
32'd144857: dataIn1 = 32'd3859
; 
32'd144858: dataIn1 = 32'd3860
; 
32'd144859: dataIn1 = 32'd3861
; 
32'd144860: dataIn1 = 32'd81
; 
32'd144861: dataIn1 = 32'd2281
; 
32'd144862: dataIn1 = 32'd3801
; 
32'd144863: dataIn1 = 32'd3859
; 
32'd144864: dataIn1 = 32'd3860
; 
32'd144865: dataIn1 = 32'd3861
; 
32'd144866: dataIn1 = 32'd3862
; 
32'd144867: dataIn1 = 32'd2257
; 
32'd144868: dataIn1 = 32'd2281
; 
32'd144869: dataIn1 = 32'd2282
; 
32'd144870: dataIn1 = 32'd3801
; 
32'd144871: dataIn1 = 32'd3861
; 
32'd144872: dataIn1 = 32'd3862
; 
32'd144873: dataIn1 = 32'd2286
; 
32'd144874: dataIn1 = 32'd2287
; 
32'd144875: dataIn1 = 32'd3863
; 
32'd144876: dataIn1 = 32'd3864
; 
32'd144877: dataIn1 = 32'd3865
; 
32'd144878: dataIn1 = 32'd10263
; 
32'd144879: dataIn1 = 32'd10272
; 
32'd144880: dataIn1 = 32'd126
; 
32'd144881: dataIn1 = 32'd2287
; 
32'd144882: dataIn1 = 32'd3863
; 
32'd144883: dataIn1 = 32'd3864
; 
32'd144884: dataIn1 = 32'd3865
; 
32'd144885: dataIn1 = 32'd4607
; 
32'd144886: dataIn1 = 32'd4610
; 
32'd144887: dataIn1 = 32'd126
; 
32'd144888: dataIn1 = 32'd2286
; 
32'd144889: dataIn1 = 32'd3863
; 
32'd144890: dataIn1 = 32'd3864
; 
32'd144891: dataIn1 = 32'd3865
; 
32'd144892: dataIn1 = 32'd3866
; 
32'd144893: dataIn1 = 32'd3867
; 
32'd144894: dataIn1 = 32'd126
; 
32'd144895: dataIn1 = 32'd2288
; 
32'd144896: dataIn1 = 32'd3865
; 
32'd144897: dataIn1 = 32'd3866
; 
32'd144898: dataIn1 = 32'd3867
; 
32'd144899: dataIn1 = 32'd5690
; 
32'd144900: dataIn1 = 32'd5951
; 
32'd144901: dataIn1 = 32'd2286
; 
32'd144902: dataIn1 = 32'd2288
; 
32'd144903: dataIn1 = 32'd2289
; 
32'd144904: dataIn1 = 32'd3865
; 
32'd144905: dataIn1 = 32'd3866
; 
32'd144906: dataIn1 = 32'd3867
; 
32'd144907: dataIn1 = 32'd1726
; 
32'd144908: dataIn1 = 32'd2295
; 
32'd144909: dataIn1 = 32'd2769
; 
32'd144910: dataIn1 = 32'd3868
; 
32'd144911: dataIn1 = 32'd3869
; 
32'd144912: dataIn1 = 32'd3870
; 
32'd144913: dataIn1 = 32'd5304
; 
32'd144914: dataIn1 = 32'd1726
; 
32'd144915: dataIn1 = 32'd2294
; 
32'd144916: dataIn1 = 32'd2770
; 
32'd144917: dataIn1 = 32'd3868
; 
32'd144918: dataIn1 = 32'd3869
; 
32'd144919: dataIn1 = 32'd3870
; 
32'd144920: dataIn1 = 32'd3933
; 
32'd144921: dataIn1 = 32'd443
; 
32'd144922: dataIn1 = 32'd2294
; 
32'd144923: dataIn1 = 32'd2295
; 
32'd144924: dataIn1 = 32'd3868
; 
32'd144925: dataIn1 = 32'd3869
; 
32'd144926: dataIn1 = 32'd3870
; 
32'd144927: dataIn1 = 32'd3871
; 
32'd144928: dataIn1 = 32'd5650
; 
32'd144929: dataIn1 = 32'd5651
; 
32'd144930: dataIn1 = 32'd5653
; 
32'd144931: dataIn1 = 32'd5655
; 
32'd144932: dataIn1 = 32'd5657
; 
32'd144933: dataIn1 = 32'd5658
; 
32'd144934: dataIn1 = 32'd2296
; 
32'd144935: dataIn1 = 32'd3872
; 
32'd144936: dataIn1 = 32'd3877
; 
32'd144937: dataIn1 = 32'd5649
; 
32'd144938: dataIn1 = 32'd5651
; 
32'd144939: dataIn1 = 32'd5654
; 
32'd144940: dataIn1 = 32'd5662
; 
32'd144941: dataIn1 = 32'd2296
; 
32'd144942: dataIn1 = 32'd3873
; 
32'd144943: dataIn1 = 32'd3879
; 
32'd144944: dataIn1 = 32'd5649
; 
32'd144945: dataIn1 = 32'd5650
; 
32'd144946: dataIn1 = 32'd5652
; 
32'd144947: dataIn1 = 32'd5663
; 
32'd144948: dataIn1 = 32'd205
; 
32'd144949: dataIn1 = 32'd3874
; 
32'd144950: dataIn1 = 32'd3897
; 
32'd144951: dataIn1 = 32'd5656
; 
32'd144952: dataIn1 = 32'd5658
; 
32'd144953: dataIn1 = 32'd5660
; 
32'd144954: dataIn1 = 32'd5686
; 
32'd144955: dataIn1 = 32'd205
; 
32'd144956: dataIn1 = 32'd3875
; 
32'd144957: dataIn1 = 32'd3890
; 
32'd144958: dataIn1 = 32'd5656
; 
32'd144959: dataIn1 = 32'd5657
; 
32'd144960: dataIn1 = 32'd5659
; 
32'd144961: dataIn1 = 32'd5671
; 
32'd144962: dataIn1 = 32'd444
; 
32'd144963: dataIn1 = 32'd3876
; 
32'd144964: dataIn1 = 32'd3877
; 
32'd144965: dataIn1 = 32'd3898
; 
32'd144966: dataIn1 = 32'd5661
; 
32'd144967: dataIn1 = 32'd5662
; 
32'd144968: dataIn1 = 32'd5687
; 
32'd144969: dataIn1 = 32'd444
; 
32'd144970: dataIn1 = 32'd2296
; 
32'd144971: dataIn1 = 32'd3872
; 
32'd144972: dataIn1 = 32'd3876
; 
32'd144973: dataIn1 = 32'd3877
; 
32'd144974: dataIn1 = 32'd3881
; 
32'd144975: dataIn1 = 32'd3885
; 
32'd144976: dataIn1 = 32'd5662
; 
32'd144977: dataIn1 = 32'd445
; 
32'd144978: dataIn1 = 32'd3878
; 
32'd144979: dataIn1 = 32'd3879
; 
32'd144980: dataIn1 = 32'd5663
; 
32'd144981: dataIn1 = 32'd5664
; 
32'd144982: dataIn1 = 32'd5673
; 
32'd144983: dataIn1 = 32'd5674
; 
32'd144984: dataIn1 = 32'd445
; 
32'd144985: dataIn1 = 32'd2296
; 
32'd144986: dataIn1 = 32'd3873
; 
32'd144987: dataIn1 = 32'd3878
; 
32'd144988: dataIn1 = 32'd3879
; 
32'd144989: dataIn1 = 32'd3882
; 
32'd144990: dataIn1 = 32'd3886
; 
32'd144991: dataIn1 = 32'd5663
; 
32'd144992: dataIn1 = 32'd2299
; 
32'd144993: dataIn1 = 32'd2300
; 
32'd144994: dataIn1 = 32'd3880
; 
32'd144995: dataIn1 = 32'd3881
; 
32'd144996: dataIn1 = 32'd3882
; 
32'd144997: dataIn1 = 32'd3883
; 
32'd144998: dataIn1 = 32'd3884
; 
32'd144999: dataIn1 = 32'd5665
; 
32'd145000: dataIn1 = 32'd5788
; 
32'd145001: dataIn1 = 32'd2296
; 
32'd145002: dataIn1 = 32'd2300
; 
32'd145003: dataIn1 = 32'd3877
; 
32'd145004: dataIn1 = 32'd3880
; 
32'd145005: dataIn1 = 32'd3881
; 
32'd145006: dataIn1 = 32'd3882
; 
32'd145007: dataIn1 = 32'd3885
; 
32'd145008: dataIn1 = 32'd2296
; 
32'd145009: dataIn1 = 32'd2299
; 
32'd145010: dataIn1 = 32'd3879
; 
32'd145011: dataIn1 = 32'd3880
; 
32'd145012: dataIn1 = 32'd3881
; 
32'd145013: dataIn1 = 32'd3882
; 
32'd145014: dataIn1 = 32'd3886
; 
32'd145015: dataIn1 = 32'd2300
; 
32'd145016: dataIn1 = 32'd3880
; 
32'd145017: dataIn1 = 32'd3883
; 
32'd145018: dataIn1 = 32'd5665
; 
32'd145019: dataIn1 = 32'd5667
; 
32'd145020: dataIn1 = 32'd5941
; 
32'd145021: dataIn1 = 32'd5943
; 
32'd145022: dataIn1 = 32'd3880
; 
32'd145023: dataIn1 = 32'd3884
; 
32'd145024: dataIn1 = 32'd5665
; 
32'd145025: dataIn1 = 32'd5666
; 
32'd145026: dataIn1 = 32'd5784
; 
32'd145027: dataIn1 = 32'd5785
; 
32'd145028: dataIn1 = 32'd5788
; 
32'd145029: dataIn1 = 32'd444
; 
32'd145030: dataIn1 = 32'd2300
; 
32'd145031: dataIn1 = 32'd3877
; 
32'd145032: dataIn1 = 32'd3881
; 
32'd145033: dataIn1 = 32'd3885
; 
32'd145034: dataIn1 = 32'd4824
; 
32'd145035: dataIn1 = 32'd4828
; 
32'd145036: dataIn1 = 32'd445
; 
32'd145037: dataIn1 = 32'd2299
; 
32'd145038: dataIn1 = 32'd3879
; 
32'd145039: dataIn1 = 32'd3882
; 
32'd145040: dataIn1 = 32'd3886
; 
32'd145041: dataIn1 = 32'd3942
; 
32'd145042: dataIn1 = 32'd3945
; 
32'd145043: dataIn1 = 32'd5780
; 
32'd145044: dataIn1 = 32'd5795
; 
32'd145045: dataIn1 = 32'd399
; 
32'd145046: dataIn1 = 32'd3887
; 
32'd145047: dataIn1 = 32'd3888
; 
32'd145048: dataIn1 = 32'd3890
; 
32'd145049: dataIn1 = 32'd5669
; 
32'd145050: dataIn1 = 32'd5670
; 
32'd145051: dataIn1 = 32'd5671
; 
32'd145052: dataIn1 = 32'd399
; 
32'd145053: dataIn1 = 32'd2301
; 
32'd145054: dataIn1 = 32'd3887
; 
32'd145055: dataIn1 = 32'd3888
; 
32'd145056: dataIn1 = 32'd3889
; 
32'd145057: dataIn1 = 32'd3891
; 
32'd145058: dataIn1 = 32'd3892
; 
32'd145059: dataIn1 = 32'd5669
; 
32'd145060: dataIn1 = 32'd5675
; 
32'd145061: dataIn1 = 32'd3888
; 
32'd145062: dataIn1 = 32'd3889
; 
32'd145063: dataIn1 = 32'd5668
; 
32'd145064: dataIn1 = 32'd5669
; 
32'd145065: dataIn1 = 32'd5672
; 
32'd145066: dataIn1 = 32'd5673
; 
32'd145067: dataIn1 = 32'd5675
; 
32'd145068: dataIn1 = 32'd205
; 
32'd145069: dataIn1 = 32'd399
; 
32'd145070: dataIn1 = 32'd3875
; 
32'd145071: dataIn1 = 32'd3887
; 
32'd145072: dataIn1 = 32'd3890
; 
32'd145073: dataIn1 = 32'd5426
; 
32'd145074: dataIn1 = 32'd5509
; 
32'd145075: dataIn1 = 32'd5671
; 
32'd145076: dataIn1 = 32'd128
; 
32'd145077: dataIn1 = 32'd399
; 
32'd145078: dataIn1 = 32'd3888
; 
32'd145079: dataIn1 = 32'd3891
; 
32'd145080: dataIn1 = 32'd3892
; 
32'd145081: dataIn1 = 32'd5427
; 
32'd145082: dataIn1 = 32'd5510
; 
32'd145083: dataIn1 = 32'd128
; 
32'd145084: dataIn1 = 32'd2301
; 
32'd145085: dataIn1 = 32'd3888
; 
32'd145086: dataIn1 = 32'd3891
; 
32'd145087: dataIn1 = 32'd3892
; 
32'd145088: dataIn1 = 32'd3925
; 
32'd145089: dataIn1 = 32'd3949
; 
32'd145090: dataIn1 = 32'd5800
; 
32'd145091: dataIn1 = 32'd445
; 
32'd145092: dataIn1 = 32'd3893
; 
32'd145093: dataIn1 = 32'd3941
; 
32'd145094: dataIn1 = 32'd5672
; 
32'd145095: dataIn1 = 32'd5674
; 
32'd145096: dataIn1 = 32'd5676
; 
32'd145097: dataIn1 = 32'd5804
; 
32'd145098: dataIn1 = 32'd3894
; 
32'd145099: dataIn1 = 32'd3897
; 
32'd145100: dataIn1 = 32'd5678
; 
32'd145101: dataIn1 = 32'd5679
; 
32'd145102: dataIn1 = 32'd5683
; 
32'd145103: dataIn1 = 32'd5685
; 
32'd145104: dataIn1 = 32'd5686
; 
32'd145105: dataIn1 = 32'd3895
; 
32'd145106: dataIn1 = 32'd3898
; 
32'd145107: dataIn1 = 32'd5677
; 
32'd145108: dataIn1 = 32'd5679
; 
32'd145109: dataIn1 = 32'd5681
; 
32'd145110: dataIn1 = 32'd5684
; 
32'd145111: dataIn1 = 32'd5687
; 
32'd145112: dataIn1 = 32'd3896
; 
32'd145113: dataIn1 = 32'd5677
; 
32'd145114: dataIn1 = 32'd5678
; 
32'd145115: dataIn1 = 32'd5680
; 
32'd145116: dataIn1 = 32'd5682
; 
32'd145117: dataIn1 = 32'd5688
; 
32'd145118: dataIn1 = 32'd5689
; 
32'd145119: dataIn1 = 32'd205
; 
32'd145120: dataIn1 = 32'd400
; 
32'd145121: dataIn1 = 32'd2489
; 
32'd145122: dataIn1 = 32'd3874
; 
32'd145123: dataIn1 = 32'd3894
; 
32'd145124: dataIn1 = 32'd3897
; 
32'd145125: dataIn1 = 32'd4602
; 
32'd145126: dataIn1 = 32'd5683
; 
32'd145127: dataIn1 = 32'd5686
; 
32'd145128: dataIn1 = 32'd444
; 
32'd145129: dataIn1 = 32'd2302
; 
32'd145130: dataIn1 = 32'd3876
; 
32'd145131: dataIn1 = 32'd3895
; 
32'd145132: dataIn1 = 32'd3898
; 
32'd145133: dataIn1 = 32'd4823
; 
32'd145134: dataIn1 = 32'd5318
; 
32'd145135: dataIn1 = 32'd5681
; 
32'd145136: dataIn1 = 32'd5687
; 
32'd145137: dataIn1 = 32'd3899
; 
32'd145138: dataIn1 = 32'd5688
; 
32'd145139: dataIn1 = 32'd5690
; 
32'd145140: dataIn1 = 32'd5691
; 
32'd145141: dataIn1 = 32'd5947
; 
32'd145142: dataIn1 = 32'd5949
; 
32'd145143: dataIn1 = 32'd5951
; 
32'd145144: dataIn1 = 32'd2304
; 
32'd145145: dataIn1 = 32'd3900
; 
32'd145146: dataIn1 = 32'd3904
; 
32'd145147: dataIn1 = 32'd5694
; 
32'd145148: dataIn1 = 32'd5695
; 
32'd145149: dataIn1 = 32'd5699
; 
32'd145150: dataIn1 = 32'd5701
; 
32'd145151: dataIn1 = 32'd3901
; 
32'd145152: dataIn1 = 32'd5693
; 
32'd145153: dataIn1 = 32'd5695
; 
32'd145154: dataIn1 = 32'd5697
; 
32'd145155: dataIn1 = 32'd5698
; 
32'd145156: dataIn1 = 32'd5702
; 
32'd145157: dataIn1 = 32'd5704
; 
32'd145158: dataIn1 = 32'd2304
; 
32'd145159: dataIn1 = 32'd3902
; 
32'd145160: dataIn1 = 32'd3907
; 
32'd145161: dataIn1 = 32'd5693
; 
32'd145162: dataIn1 = 32'd5694
; 
32'd145163: dataIn1 = 32'd5696
; 
32'd145164: dataIn1 = 32'd5707
; 
32'd145165: dataIn1 = 32'd446
; 
32'd145166: dataIn1 = 32'd3903
; 
32'd145167: dataIn1 = 32'd3904
; 
32'd145168: dataIn1 = 32'd5700
; 
32'd145169: dataIn1 = 32'd5701
; 
32'd145170: dataIn1 = 32'd5752
; 
32'd145171: dataIn1 = 32'd5754
; 
32'd145172: dataIn1 = 32'd446
; 
32'd145173: dataIn1 = 32'd2304
; 
32'd145174: dataIn1 = 32'd3900
; 
32'd145175: dataIn1 = 32'd3903
; 
32'd145176: dataIn1 = 32'd3904
; 
32'd145177: dataIn1 = 32'd3914
; 
32'd145178: dataIn1 = 32'd3917
; 
32'd145179: dataIn1 = 32'd5701
; 
32'd145180: dataIn1 = 32'd5735
; 
32'd145181: dataIn1 = 32'd206
; 
32'd145182: dataIn1 = 32'd2293
; 
32'd145183: dataIn1 = 32'd3905
; 
32'd145184: dataIn1 = 32'd5703
; 
32'd145185: dataIn1 = 32'd5704
; 
32'd145186: dataIn1 = 32'd5706
; 
32'd145187: dataIn1 = 32'd5756
; 
32'd145188: dataIn1 = 32'd206
; 
32'd145189: dataIn1 = 32'd2527
; 
32'd145190: dataIn1 = 32'd3906
; 
32'd145191: dataIn1 = 32'd5702
; 
32'd145192: dataIn1 = 32'd5703
; 
32'd145193: dataIn1 = 32'd5705
; 
32'd145194: dataIn1 = 32'd5725
; 
32'd145195: dataIn1 = 32'd447
; 
32'd145196: dataIn1 = 32'd2304
; 
32'd145197: dataIn1 = 32'd3902
; 
32'd145198: dataIn1 = 32'd3907
; 
32'd145199: dataIn1 = 32'd3908
; 
32'd145200: dataIn1 = 32'd3916
; 
32'd145201: dataIn1 = 32'd3920
; 
32'd145202: dataIn1 = 32'd5707
; 
32'd145203: dataIn1 = 32'd5743
; 
32'd145204: dataIn1 = 32'd447
; 
32'd145205: dataIn1 = 32'd3907
; 
32'd145206: dataIn1 = 32'd3908
; 
32'd145207: dataIn1 = 32'd3913
; 
32'd145208: dataIn1 = 32'd5707
; 
32'd145209: dataIn1 = 32'd5708
; 
32'd145210: dataIn1 = 32'd5726
; 
32'd145211: dataIn1 = 32'd3909
; 
32'd145212: dataIn1 = 32'd5710
; 
32'd145213: dataIn1 = 32'd5711
; 
32'd145214: dataIn1 = 32'd5715
; 
32'd145215: dataIn1 = 32'd5717
; 
32'd145216: dataIn1 = 32'd5719
; 
32'd145217: dataIn1 = 32'd5720
; 
32'd145218: dataIn1 = 32'd2527
; 
32'd145219: dataIn1 = 32'd3910
; 
32'd145220: dataIn1 = 32'd5709
; 
32'd145221: dataIn1 = 32'd5711
; 
32'd145222: dataIn1 = 32'd5713
; 
32'd145223: dataIn1 = 32'd5716
; 
32'd145224: dataIn1 = 32'd5725
; 
32'd145225: dataIn1 = 32'd3911
; 
32'd145226: dataIn1 = 32'd3913
; 
32'd145227: dataIn1 = 32'd5709
; 
32'd145228: dataIn1 = 32'd5710
; 
32'd145229: dataIn1 = 32'd5712
; 
32'd145230: dataIn1 = 32'd5714
; 
32'd145231: dataIn1 = 32'd5726
; 
32'd145232: dataIn1 = 32'd3912
; 
32'd145233: dataIn1 = 32'd5718
; 
32'd145234: dataIn1 = 32'd5719
; 
32'd145235: dataIn1 = 32'd5721
; 
32'd145236: dataIn1 = 32'd5723
; 
32'd145237: dataIn1 = 32'd6062
; 
32'd145238: dataIn1 = 32'd6063
; 
32'd145239: dataIn1 = 32'd447
; 
32'd145240: dataIn1 = 32'd2306
; 
32'd145241: dataIn1 = 32'd3908
; 
32'd145242: dataIn1 = 32'd3911
; 
32'd145243: dataIn1 = 32'd3913
; 
32'd145244: dataIn1 = 32'd4865
; 
32'd145245: dataIn1 = 32'd4881
; 
32'd145246: dataIn1 = 32'd5714
; 
32'd145247: dataIn1 = 32'd5726
; 
32'd145248: dataIn1 = 32'd2304
; 
32'd145249: dataIn1 = 32'd3904
; 
32'd145250: dataIn1 = 32'd3914
; 
32'd145251: dataIn1 = 32'd5728
; 
32'd145252: dataIn1 = 32'd5729
; 
32'd145253: dataIn1 = 32'd5733
; 
32'd145254: dataIn1 = 32'd5735
; 
32'd145255: dataIn1 = 32'd3915
; 
32'd145256: dataIn1 = 32'd5727
; 
32'd145257: dataIn1 = 32'd5729
; 
32'd145258: dataIn1 = 32'd5731
; 
32'd145259: dataIn1 = 32'd5732
; 
32'd145260: dataIn1 = 32'd5736
; 
32'd145261: dataIn1 = 32'd5738
; 
32'd145262: dataIn1 = 32'd2304
; 
32'd145263: dataIn1 = 32'd3907
; 
32'd145264: dataIn1 = 32'd3916
; 
32'd145265: dataIn1 = 32'd5727
; 
32'd145266: dataIn1 = 32'd5728
; 
32'd145267: dataIn1 = 32'd5730
; 
32'd145268: dataIn1 = 32'd5743
; 
32'd145269: dataIn1 = 32'd446
; 
32'd145270: dataIn1 = 32'd3904
; 
32'd145271: dataIn1 = 32'd3917
; 
32'd145272: dataIn1 = 32'd5734
; 
32'd145273: dataIn1 = 32'd5735
; 
32'd145274: dataIn1 = 32'd5814
; 
32'd145275: dataIn1 = 32'd5815
; 
32'd145276: dataIn1 = 32'd3918
; 
32'd145277: dataIn1 = 32'd5737
; 
32'd145278: dataIn1 = 32'd5738
; 
32'd145279: dataIn1 = 32'd5741
; 
32'd145280: dataIn1 = 32'd5742
; 
32'd145281: dataIn1 = 32'd5823
; 
32'd145282: dataIn1 = 32'd5824
; 
32'd145283: dataIn1 = 32'd3919
; 
32'd145284: dataIn1 = 32'd5736
; 
32'd145285: dataIn1 = 32'd5737
; 
32'd145286: dataIn1 = 32'd5739
; 
32'd145287: dataIn1 = 32'd5740
; 
32'd145288: dataIn1 = 32'd6053
; 
32'd145289: dataIn1 = 32'd6054
; 
32'd145290: dataIn1 = 32'd447
; 
32'd145291: dataIn1 = 32'd3907
; 
32'd145292: dataIn1 = 32'd3920
; 
32'd145293: dataIn1 = 32'd5743
; 
32'd145294: dataIn1 = 32'd5744
; 
32'd145295: dataIn1 = 32'd6696
; 
32'd145296: dataIn1 = 32'd6732
; 
32'd145297: dataIn1 = 32'd3921
; 
32'd145298: dataIn1 = 32'd5746
; 
32'd145299: dataIn1 = 32'd5747
; 
32'd145300: dataIn1 = 32'd5749
; 
32'd145301: dataIn1 = 32'd5751
; 
32'd145302: dataIn1 = 32'd5753
; 
32'd145303: dataIn1 = 32'd5754
; 
32'd145304: dataIn1 = 32'd404
; 
32'd145305: dataIn1 = 32'd2293
; 
32'd145306: dataIn1 = 32'd3922
; 
32'd145307: dataIn1 = 32'd5745
; 
32'd145308: dataIn1 = 32'd5747
; 
32'd145309: dataIn1 = 32'd5750
; 
32'd145310: dataIn1 = 32'd5756
; 
32'd145311: dataIn1 = 32'd404
; 
32'd145312: dataIn1 = 32'd3923
; 
32'd145313: dataIn1 = 32'd3925
; 
32'd145314: dataIn1 = 32'd3926
; 
32'd145315: dataIn1 = 32'd5745
; 
32'd145316: dataIn1 = 32'd5746
; 
32'd145317: dataIn1 = 32'd5748
; 
32'd145318: dataIn1 = 32'd446
; 
32'd145319: dataIn1 = 32'd3924
; 
32'd145320: dataIn1 = 32'd3938
; 
32'd145321: dataIn1 = 32'd5752
; 
32'd145322: dataIn1 = 32'd5753
; 
32'd145323: dataIn1 = 32'd5755
; 
32'd145324: dataIn1 = 32'd5803
; 
32'd145325: dataIn1 = 32'd128
; 
32'd145326: dataIn1 = 32'd2309
; 
32'd145327: dataIn1 = 32'd3892
; 
32'd145328: dataIn1 = 32'd3923
; 
32'd145329: dataIn1 = 32'd3925
; 
32'd145330: dataIn1 = 32'd3926
; 
32'd145331: dataIn1 = 32'd3949
; 
32'd145332: dataIn1 = 32'd5748
; 
32'd145333: dataIn1 = 32'd5801
; 
32'd145334: dataIn1 = 32'd128
; 
32'd145335: dataIn1 = 32'd404
; 
32'd145336: dataIn1 = 32'd2490
; 
32'd145337: dataIn1 = 32'd3923
; 
32'd145338: dataIn1 = 32'd3925
; 
32'd145339: dataIn1 = 32'd3926
; 
32'd145340: dataIn1 = 32'd4603
; 
32'd145341: dataIn1 = 32'd2310
; 
32'd145342: dataIn1 = 32'd2311
; 
32'd145343: dataIn1 = 32'd3927
; 
32'd145344: dataIn1 = 32'd3928
; 
32'd145345: dataIn1 = 32'd3929
; 
32'd145346: dataIn1 = 32'd3930
; 
32'd145347: dataIn1 = 32'd3931
; 
32'd145348: dataIn1 = 32'd2294
; 
32'd145349: dataIn1 = 32'd2311
; 
32'd145350: dataIn1 = 32'd3927
; 
32'd145351: dataIn1 = 32'd3928
; 
32'd145352: dataIn1 = 32'd3929
; 
32'd145353: dataIn1 = 32'd3932
; 
32'd145354: dataIn1 = 32'd3933
; 
32'd145355: dataIn1 = 32'd443
; 
32'd145356: dataIn1 = 32'd2294
; 
32'd145357: dataIn1 = 32'd2310
; 
32'd145358: dataIn1 = 32'd3927
; 
32'd145359: dataIn1 = 32'd3928
; 
32'd145360: dataIn1 = 32'd3929
; 
32'd145361: dataIn1 = 32'd448
; 
32'd145362: dataIn1 = 32'd2311
; 
32'd145363: dataIn1 = 32'd3927
; 
32'd145364: dataIn1 = 32'd3930
; 
32'd145365: dataIn1 = 32'd3931
; 
32'd145366: dataIn1 = 32'd3956
; 
32'd145367: dataIn1 = 32'd3959
; 
32'd145368: dataIn1 = 32'd448
; 
32'd145369: dataIn1 = 32'd2310
; 
32'd145370: dataIn1 = 32'd3927
; 
32'd145371: dataIn1 = 32'd3930
; 
32'd145372: dataIn1 = 32'd3931
; 
32'd145373: dataIn1 = 32'd5320
; 
32'd145374: dataIn1 = 32'd154
; 
32'd145375: dataIn1 = 32'd2311
; 
32'd145376: dataIn1 = 32'd3928
; 
32'd145377: dataIn1 = 32'd3932
; 
32'd145378: dataIn1 = 32'd3933
; 
32'd145379: dataIn1 = 32'd3957
; 
32'd145380: dataIn1 = 32'd3960
; 
32'd145381: dataIn1 = 32'd154
; 
32'd145382: dataIn1 = 32'd2294
; 
32'd145383: dataIn1 = 32'd2770
; 
32'd145384: dataIn1 = 32'd3869
; 
32'd145385: dataIn1 = 32'd3928
; 
32'd145386: dataIn1 = 32'd3932
; 
32'd145387: dataIn1 = 32'd3933
; 
32'd145388: dataIn1 = 32'd2313
; 
32'd145389: dataIn1 = 32'd3934
; 
32'd145390: dataIn1 = 32'd3938
; 
32'd145391: dataIn1 = 32'd5758
; 
32'd145392: dataIn1 = 32'd5759
; 
32'd145393: dataIn1 = 32'd5763
; 
32'd145394: dataIn1 = 32'd5765
; 
32'd145395: dataIn1 = 32'd3935
; 
32'd145396: dataIn1 = 32'd5757
; 
32'd145397: dataIn1 = 32'd5759
; 
32'd145398: dataIn1 = 32'd5761
; 
32'd145399: dataIn1 = 32'd5762
; 
32'd145400: dataIn1 = 32'd5766
; 
32'd145401: dataIn1 = 32'd5768
; 
32'd145402: dataIn1 = 32'd2313
; 
32'd145403: dataIn1 = 32'd3936
; 
32'd145404: dataIn1 = 32'd3941
; 
32'd145405: dataIn1 = 32'd5757
; 
32'd145406: dataIn1 = 32'd5758
; 
32'd145407: dataIn1 = 32'd5760
; 
32'd145408: dataIn1 = 32'd5773
; 
32'd145409: dataIn1 = 32'd446
; 
32'd145410: dataIn1 = 32'd3937
; 
32'd145411: dataIn1 = 32'd3938
; 
32'd145412: dataIn1 = 32'd5764
; 
32'd145413: dataIn1 = 32'd5765
; 
32'd145414: dataIn1 = 32'd5814
; 
32'd145415: dataIn1 = 32'd5816
; 
32'd145416: dataIn1 = 32'd446
; 
32'd145417: dataIn1 = 32'd2313
; 
32'd145418: dataIn1 = 32'd3924
; 
32'd145419: dataIn1 = 32'd3934
; 
32'd145420: dataIn1 = 32'd3937
; 
32'd145421: dataIn1 = 32'd3938
; 
32'd145422: dataIn1 = 32'd3948
; 
32'd145423: dataIn1 = 32'd5765
; 
32'd145424: dataIn1 = 32'd5803
; 
32'd145425: dataIn1 = 32'd3939
; 
32'd145426: dataIn1 = 32'd5767
; 
32'd145427: dataIn1 = 32'd5768
; 
32'd145428: dataIn1 = 32'd5771
; 
32'd145429: dataIn1 = 32'd5772
; 
32'd145430: dataIn1 = 32'd5818
; 
32'd145431: dataIn1 = 32'd5819
; 
32'd145432: dataIn1 = 32'd3940
; 
32'd145433: dataIn1 = 32'd5766
; 
32'd145434: dataIn1 = 32'd5767
; 
32'd145435: dataIn1 = 32'd5769
; 
32'd145436: dataIn1 = 32'd5770
; 
32'd145437: dataIn1 = 32'd5790
; 
32'd145438: dataIn1 = 32'd5791
; 
32'd145439: dataIn1 = 32'd445
; 
32'd145440: dataIn1 = 32'd2313
; 
32'd145441: dataIn1 = 32'd3893
; 
32'd145442: dataIn1 = 32'd3936
; 
32'd145443: dataIn1 = 32'd3941
; 
32'd145444: dataIn1 = 32'd3942
; 
32'd145445: dataIn1 = 32'd3950
; 
32'd145446: dataIn1 = 32'd5773
; 
32'd145447: dataIn1 = 32'd5804
; 
32'd145448: dataIn1 = 32'd445
; 
32'd145449: dataIn1 = 32'd3886
; 
32'd145450: dataIn1 = 32'd3941
; 
32'd145451: dataIn1 = 32'd3942
; 
32'd145452: dataIn1 = 32'd5773
; 
32'd145453: dataIn1 = 32'd5774
; 
32'd145454: dataIn1 = 32'd5795
; 
32'd145455: dataIn1 = 32'd3943
; 
32'd145456: dataIn1 = 32'd5776
; 
32'd145457: dataIn1 = 32'd5777
; 
32'd145458: dataIn1 = 32'd5781
; 
32'd145459: dataIn1 = 32'd5783
; 
32'd145460: dataIn1 = 32'd5785
; 
32'd145461: dataIn1 = 32'd5786
; 
32'd145462: dataIn1 = 32'd3944
; 
32'd145463: dataIn1 = 32'd5775
; 
32'd145464: dataIn1 = 32'd5777
; 
32'd145465: dataIn1 = 32'd5779
; 
32'd145466: dataIn1 = 32'd5782
; 
32'd145467: dataIn1 = 32'd5790
; 
32'd145468: dataIn1 = 32'd5792
; 
32'd145469: dataIn1 = 32'd3886
; 
32'd145470: dataIn1 = 32'd3945
; 
32'd145471: dataIn1 = 32'd5775
; 
32'd145472: dataIn1 = 32'd5776
; 
32'd145473: dataIn1 = 32'd5778
; 
32'd145474: dataIn1 = 32'd5780
; 
32'd145475: dataIn1 = 32'd5795
; 
32'd145476: dataIn1 = 32'd3946
; 
32'd145477: dataIn1 = 32'd5784
; 
32'd145478: dataIn1 = 32'd5786
; 
32'd145479: dataIn1 = 32'd5787
; 
32'd145480: dataIn1 = 32'd5789
; 
32'd145481: dataIn1 = 32'd7030
; 
32'd145482: dataIn1 = 32'd7031
; 
32'd145483: dataIn1 = 32'd3947
; 
32'd145484: dataIn1 = 32'd5791
; 
32'd145485: dataIn1 = 32'd5792
; 
32'd145486: dataIn1 = 32'd5793
; 
32'd145487: dataIn1 = 32'd5794
; 
32'd145488: dataIn1 = 32'd7026
; 
32'd145489: dataIn1 = 32'd7028
; 
32'd145490: dataIn1 = 32'd2313
; 
32'd145491: dataIn1 = 32'd3938
; 
32'd145492: dataIn1 = 32'd3948
; 
32'd145493: dataIn1 = 32'd5797
; 
32'd145494: dataIn1 = 32'd5798
; 
32'd145495: dataIn1 = 32'd5802
; 
32'd145496: dataIn1 = 32'd5803
; 
32'd145497: dataIn1 = 32'd3892
; 
32'd145498: dataIn1 = 32'd3925
; 
32'd145499: dataIn1 = 32'd3949
; 
32'd145500: dataIn1 = 32'd5796
; 
32'd145501: dataIn1 = 32'd5798
; 
32'd145502: dataIn1 = 32'd5800
; 
32'd145503: dataIn1 = 32'd5801
; 
32'd145504: dataIn1 = 32'd2313
; 
32'd145505: dataIn1 = 32'd3941
; 
32'd145506: dataIn1 = 32'd3950
; 
32'd145507: dataIn1 = 32'd5796
; 
32'd145508: dataIn1 = 32'd5797
; 
32'd145509: dataIn1 = 32'd5799
; 
32'd145510: dataIn1 = 32'd5804
; 
32'd145511: dataIn1 = 32'd3951
; 
32'd145512: dataIn1 = 32'd5806
; 
32'd145513: dataIn1 = 32'd5807
; 
32'd145514: dataIn1 = 32'd5811
; 
32'd145515: dataIn1 = 32'd5813
; 
32'd145516: dataIn1 = 32'd5815
; 
32'd145517: dataIn1 = 32'd5816
; 
32'd145518: dataIn1 = 32'd3952
; 
32'd145519: dataIn1 = 32'd5805
; 
32'd145520: dataIn1 = 32'd5807
; 
32'd145521: dataIn1 = 32'd5809
; 
32'd145522: dataIn1 = 32'd5812
; 
32'd145523: dataIn1 = 32'd5817
; 
32'd145524: dataIn1 = 32'd5819
; 
32'd145525: dataIn1 = 32'd3953
; 
32'd145526: dataIn1 = 32'd5805
; 
32'd145527: dataIn1 = 32'd5806
; 
32'd145528: dataIn1 = 32'd5808
; 
32'd145529: dataIn1 = 32'd5810
; 
32'd145530: dataIn1 = 32'd5822
; 
32'd145531: dataIn1 = 32'd5823
; 
32'd145532: dataIn1 = 32'd3954
; 
32'd145533: dataIn1 = 32'd5817
; 
32'd145534: dataIn1 = 32'd5818
; 
32'd145535: dataIn1 = 32'd5820
; 
32'd145536: dataIn1 = 32'd5821
; 
32'd145537: dataIn1 = 32'd7044
; 
32'd145538: dataIn1 = 32'd7045
; 
32'd145539: dataIn1 = 32'd3955
; 
32'd145540: dataIn1 = 32'd5822
; 
32'd145541: dataIn1 = 32'd5824
; 
32'd145542: dataIn1 = 32'd5825
; 
32'd145543: dataIn1 = 32'd5826
; 
32'd145544: dataIn1 = 32'd7052
; 
32'd145545: dataIn1 = 32'd7053
; 
32'd145546: dataIn1 = 32'd2311
; 
32'd145547: dataIn1 = 32'd2318
; 
32'd145548: dataIn1 = 32'd3930
; 
32'd145549: dataIn1 = 32'd3956
; 
32'd145550: dataIn1 = 32'd3957
; 
32'd145551: dataIn1 = 32'd3958
; 
32'd145552: dataIn1 = 32'd3959
; 
32'd145553: dataIn1 = 32'd2311
; 
32'd145554: dataIn1 = 32'd2317
; 
32'd145555: dataIn1 = 32'd3932
; 
32'd145556: dataIn1 = 32'd3956
; 
32'd145557: dataIn1 = 32'd3957
; 
32'd145558: dataIn1 = 32'd3958
; 
32'd145559: dataIn1 = 32'd3960
; 
32'd145560: dataIn1 = 32'd2317
; 
32'd145561: dataIn1 = 32'd2318
; 
32'd145562: dataIn1 = 32'd3956
; 
32'd145563: dataIn1 = 32'd3957
; 
32'd145564: dataIn1 = 32'd3958
; 
32'd145565: dataIn1 = 32'd3961
; 
32'd145566: dataIn1 = 32'd3962
; 
32'd145567: dataIn1 = 32'd448
; 
32'd145568: dataIn1 = 32'd2318
; 
32'd145569: dataIn1 = 32'd3930
; 
32'd145570: dataIn1 = 32'd3956
; 
32'd145571: dataIn1 = 32'd3959
; 
32'd145572: dataIn1 = 32'd5322
; 
32'd145573: dataIn1 = 32'd154
; 
32'd145574: dataIn1 = 32'd2317
; 
32'd145575: dataIn1 = 32'd3052
; 
32'd145576: dataIn1 = 32'd3932
; 
32'd145577: dataIn1 = 32'd3957
; 
32'd145578: dataIn1 = 32'd3960
; 
32'd145579: dataIn1 = 32'd3996
; 
32'd145580: dataIn1 = 32'd450
; 
32'd145581: dataIn1 = 32'd2318
; 
32'd145582: dataIn1 = 32'd3958
; 
32'd145583: dataIn1 = 32'd3961
; 
32'd145584: dataIn1 = 32'd3962
; 
32'd145585: dataIn1 = 32'd5321
; 
32'd145586: dataIn1 = 32'd450
; 
32'd145587: dataIn1 = 32'd2317
; 
32'd145588: dataIn1 = 32'd3958
; 
32'd145589: dataIn1 = 32'd3961
; 
32'd145590: dataIn1 = 32'd3962
; 
32'd145591: dataIn1 = 32'd3993
; 
32'd145592: dataIn1 = 32'd3997
; 
32'd145593: dataIn1 = 32'd3963
; 
32'd145594: dataIn1 = 32'd3967
; 
32'd145595: dataIn1 = 32'd5835
; 
32'd145596: dataIn1 = 32'd6854
; 
32'd145597: dataIn1 = 32'd6855
; 
32'd145598: dataIn1 = 32'd6870
; 
32'd145599: dataIn1 = 32'd9271
; 
32'd145600: dataIn1 = 32'd3964
; 
32'd145601: dataIn1 = 32'd6856
; 
32'd145602: dataIn1 = 32'd6857
; 
32'd145603: dataIn1 = 32'd6865
; 
32'd145604: dataIn1 = 32'd6871
; 
32'd145605: dataIn1 = 32'd6879
; 
32'd145606: dataIn1 = 32'd6880
; 
32'd145607: dataIn1 = 32'd3965
; 
32'd145608: dataIn1 = 32'd5844
; 
32'd145609: dataIn1 = 32'd6858
; 
32'd145610: dataIn1 = 32'd6859
; 
32'd145611: dataIn1 = 32'd6866
; 
32'd145612: dataIn1 = 32'd6906
; 
32'd145613: dataIn1 = 32'd9270
; 
32'd145614: dataIn1 = 32'd451
; 
32'd145615: dataIn1 = 32'd3966
; 
32'd145616: dataIn1 = 32'd3967
; 
32'd145617: dataIn1 = 32'd5834
; 
32'd145618: dataIn1 = 32'd5835
; 
32'd145619: dataIn1 = 32'd5880
; 
32'd145620: dataIn1 = 32'd9320
; 
32'd145621: dataIn1 = 32'd451
; 
32'd145622: dataIn1 = 32'd2320
; 
32'd145623: dataIn1 = 32'd3963
; 
32'd145624: dataIn1 = 32'd3966
; 
32'd145625: dataIn1 = 32'd3967
; 
32'd145626: dataIn1 = 32'd3977
; 
32'd145627: dataIn1 = 32'd5323
; 
32'd145628: dataIn1 = 32'd5835
; 
32'd145629: dataIn1 = 32'd9271
; 
32'd145630: dataIn1 = 32'd3968
; 
32'd145631: dataIn1 = 32'd6877
; 
32'd145632: dataIn1 = 32'd6878
; 
32'd145633: dataIn1 = 32'd6891
; 
32'd145634: dataIn1 = 32'd6898
; 
32'd145635: dataIn1 = 32'd7020
; 
32'd145636: dataIn1 = 32'd7021
; 
32'd145637: dataIn1 = 32'd3969
; 
32'd145638: dataIn1 = 32'd6881
; 
32'd145639: dataIn1 = 32'd6882
; 
32'd145640: dataIn1 = 32'd6887
; 
32'd145641: dataIn1 = 32'd6894
; 
32'd145642: dataIn1 = 32'd6959
; 
32'd145643: dataIn1 = 32'd6960
; 
32'd145644: dataIn1 = 32'd3970
; 
32'd145645: dataIn1 = 32'd3979
; 
32'd145646: dataIn1 = 32'd3980
; 
32'd145647: dataIn1 = 32'd5844
; 
32'd145648: dataIn1 = 32'd5845
; 
32'd145649: dataIn1 = 32'd5848
; 
32'd145650: dataIn1 = 32'd9319
; 
32'd145651: dataIn1 = 32'd3971
; 
32'd145652: dataIn1 = 32'd5845
; 
32'd145653: dataIn1 = 32'd5847
; 
32'd145654: dataIn1 = 32'd6904
; 
32'd145655: dataIn1 = 32'd6905
; 
32'd145656: dataIn1 = 32'd6977
; 
32'd145657: dataIn1 = 32'd6978
; 
32'd145658: dataIn1 = 32'd3972
; 
32'd145659: dataIn1 = 32'd6910
; 
32'd145660: dataIn1 = 32'd6911
; 
32'd145661: dataIn1 = 32'd6926
; 
32'd145662: dataIn1 = 32'd6933
; 
32'd145663: dataIn1 = 32'd6940
; 
32'd145664: dataIn1 = 32'd6941
; 
32'd145665: dataIn1 = 32'd3973
; 
32'd145666: dataIn1 = 32'd6912
; 
32'd145667: dataIn1 = 32'd6913
; 
32'd145668: dataIn1 = 32'd6921
; 
32'd145669: dataIn1 = 32'd6934
; 
32'd145670: dataIn1 = 32'd6957
; 
32'd145671: dataIn1 = 32'd6958
; 
32'd145672: dataIn1 = 32'd3974
; 
32'd145673: dataIn1 = 32'd6914
; 
32'd145674: dataIn1 = 32'd6915
; 
32'd145675: dataIn1 = 32'd6922
; 
32'd145676: dataIn1 = 32'd6929
; 
32'd145677: dataIn1 = 32'd6979
; 
32'd145678: dataIn1 = 32'd6980
; 
32'd145679: dataIn1 = 32'd3975
; 
32'd145680: dataIn1 = 32'd6942
; 
32'd145681: dataIn1 = 32'd6943
; 
32'd145682: dataIn1 = 32'd6944
; 
32'd145683: dataIn1 = 32'd6950
; 
32'd145684: dataIn1 = 32'd8898
; 
32'd145685: dataIn1 = 32'd8899
; 
32'd145686: dataIn1 = 32'd3976
; 
32'd145687: dataIn1 = 32'd5870
; 
32'd145688: dataIn1 = 32'd6586
; 
32'd145689: dataIn1 = 32'd6975
; 
32'd145690: dataIn1 = 32'd6976
; 
32'd145691: dataIn1 = 32'd6987
; 
32'd145692: dataIn1 = 32'd8914
; 
32'd145693: dataIn1 = 32'd2320
; 
32'd145694: dataIn1 = 32'd2324
; 
32'd145695: dataIn1 = 32'd3967
; 
32'd145696: dataIn1 = 32'd3977
; 
32'd145697: dataIn1 = 32'd3978
; 
32'd145698: dataIn1 = 32'd3979
; 
32'd145699: dataIn1 = 32'd5323
; 
32'd145700: dataIn1 = 32'd15
; 
32'd145701: dataIn1 = 32'd2323
; 
32'd145702: dataIn1 = 32'd2324
; 
32'd145703: dataIn1 = 32'd3977
; 
32'd145704: dataIn1 = 32'd3978
; 
32'd145705: dataIn1 = 32'd3979
; 
32'd145706: dataIn1 = 32'd2320
; 
32'd145707: dataIn1 = 32'd2323
; 
32'd145708: dataIn1 = 32'd3970
; 
32'd145709: dataIn1 = 32'd3977
; 
32'd145710: dataIn1 = 32'd3978
; 
32'd145711: dataIn1 = 32'd3979
; 
32'd145712: dataIn1 = 32'd3980
; 
32'd145713: dataIn1 = 32'd9319
; 
32'd145714: dataIn1 = 32'd452
; 
32'd145715: dataIn1 = 32'd2323
; 
32'd145716: dataIn1 = 32'd3970
; 
32'd145717: dataIn1 = 32'd3979
; 
32'd145718: dataIn1 = 32'd3980
; 
32'd145719: dataIn1 = 32'd5848
; 
32'd145720: dataIn1 = 32'd6717
; 
32'd145721: dataIn1 = 32'd6742
; 
32'd145722: dataIn1 = 32'd3981
; 
32'd145723: dataIn1 = 32'd5880
; 
32'd145724: dataIn1 = 32'd6992
; 
32'd145725: dataIn1 = 32'd6993
; 
32'd145726: dataIn1 = 32'd7008
; 
32'd145727: dataIn1 = 32'd7013
; 
32'd145728: dataIn1 = 32'd9273
; 
32'd145729: dataIn1 = 32'd3982
; 
32'd145730: dataIn1 = 32'd6994
; 
32'd145731: dataIn1 = 32'd6995
; 
32'd145732: dataIn1 = 32'd7003
; 
32'd145733: dataIn1 = 32'd7014
; 
32'd145734: dataIn1 = 32'd7022
; 
32'd145735: dataIn1 = 32'd7023
; 
32'd145736: dataIn1 = 32'd3983
; 
32'd145737: dataIn1 = 32'd6996
; 
32'd145738: dataIn1 = 32'd6997
; 
32'd145739: dataIn1 = 32'd7004
; 
32'd145740: dataIn1 = 32'd7009
; 
32'd145741: dataIn1 = 32'd7042
; 
32'd145742: dataIn1 = 32'd7043
; 
32'd145743: dataIn1 = 32'd451
; 
32'd145744: dataIn1 = 32'd3984
; 
32'd145745: dataIn1 = 32'd5271
; 
32'd145746: dataIn1 = 32'd5273
; 
32'd145747: dataIn1 = 32'd9272
; 
32'd145748: dataIn1 = 32'd9273
; 
32'd145749: dataIn1 = 32'd9320
; 
32'd145750: dataIn1 = 32'd3985
; 
32'd145751: dataIn1 = 32'd7038
; 
32'd145752: dataIn1 = 32'd7039
; 
32'd145753: dataIn1 = 32'd7050
; 
32'd145754: dataIn1 = 32'd7054
; 
32'd145755: dataIn1 = 32'd8926
; 
32'd145756: dataIn1 = 32'd9768
; 
32'd145757: dataIn1 = 32'd2327
; 
32'd145758: dataIn1 = 32'd2328
; 
32'd145759: dataIn1 = 32'd3986
; 
32'd145760: dataIn1 = 32'd3987
; 
32'd145761: dataIn1 = 32'd3988
; 
32'd145762: dataIn1 = 32'd3989
; 
32'd145763: dataIn1 = 32'd3990
; 
32'd145764: dataIn1 = 32'd2326
; 
32'd145765: dataIn1 = 32'd2328
; 
32'd145766: dataIn1 = 32'd3986
; 
32'd145767: dataIn1 = 32'd3987
; 
32'd145768: dataIn1 = 32'd3988
; 
32'd145769: dataIn1 = 32'd3991
; 
32'd145770: dataIn1 = 32'd3992
; 
32'd145771: dataIn1 = 32'd2326
; 
32'd145772: dataIn1 = 32'd2327
; 
32'd145773: dataIn1 = 32'd3986
; 
32'd145774: dataIn1 = 32'd3987
; 
32'd145775: dataIn1 = 32'd3988
; 
32'd145776: dataIn1 = 32'd3993
; 
32'd145777: dataIn1 = 32'd3994
; 
32'd145778: dataIn1 = 32'd279
; 
32'd145779: dataIn1 = 32'd2328
; 
32'd145780: dataIn1 = 32'd3044
; 
32'd145781: dataIn1 = 32'd3986
; 
32'd145782: dataIn1 = 32'd3989
; 
32'd145783: dataIn1 = 32'd3990
; 
32'd145784: dataIn1 = 32'd3998
; 
32'd145785: dataIn1 = 32'd279
; 
32'd145786: dataIn1 = 32'd2327
; 
32'd145787: dataIn1 = 32'd3051
; 
32'd145788: dataIn1 = 32'd3986
; 
32'd145789: dataIn1 = 32'd3989
; 
32'd145790: dataIn1 = 32'd3990
; 
32'd145791: dataIn1 = 32'd3995
; 
32'd145792: dataIn1 = 32'd453
; 
32'd145793: dataIn1 = 32'd2328
; 
32'd145794: dataIn1 = 32'd3987
; 
32'd145795: dataIn1 = 32'd3991
; 
32'd145796: dataIn1 = 32'd3992
; 
32'd145797: dataIn1 = 32'd3999
; 
32'd145798: dataIn1 = 32'd4001
; 
32'd145799: dataIn1 = 32'd453
; 
32'd145800: dataIn1 = 32'd2326
; 
32'd145801: dataIn1 = 32'd3987
; 
32'd145802: dataIn1 = 32'd3991
; 
32'd145803: dataIn1 = 32'd3992
; 
32'd145804: dataIn1 = 32'd5325
; 
32'd145805: dataIn1 = 32'd450
; 
32'd145806: dataIn1 = 32'd2327
; 
32'd145807: dataIn1 = 32'd3962
; 
32'd145808: dataIn1 = 32'd3988
; 
32'd145809: dataIn1 = 32'd3993
; 
32'd145810: dataIn1 = 32'd3994
; 
32'd145811: dataIn1 = 32'd3997
; 
32'd145812: dataIn1 = 32'd450
; 
32'd145813: dataIn1 = 32'd2326
; 
32'd145814: dataIn1 = 32'd3988
; 
32'd145815: dataIn1 = 32'd3993
; 
32'd145816: dataIn1 = 32'd3994
; 
32'd145817: dataIn1 = 32'd5324
; 
32'd145818: dataIn1 = 32'd1978
; 
32'd145819: dataIn1 = 32'd2327
; 
32'd145820: dataIn1 = 32'd3051
; 
32'd145821: dataIn1 = 32'd3990
; 
32'd145822: dataIn1 = 32'd3995
; 
32'd145823: dataIn1 = 32'd3996
; 
32'd145824: dataIn1 = 32'd3997
; 
32'd145825: dataIn1 = 32'd1978
; 
32'd145826: dataIn1 = 32'd2317
; 
32'd145827: dataIn1 = 32'd3052
; 
32'd145828: dataIn1 = 32'd3960
; 
32'd145829: dataIn1 = 32'd3995
; 
32'd145830: dataIn1 = 32'd3996
; 
32'd145831: dataIn1 = 32'd3997
; 
32'd145832: dataIn1 = 32'd2317
; 
32'd145833: dataIn1 = 32'd2327
; 
32'd145834: dataIn1 = 32'd3962
; 
32'd145835: dataIn1 = 32'd3993
; 
32'd145836: dataIn1 = 32'd3995
; 
32'd145837: dataIn1 = 32'd3996
; 
32'd145838: dataIn1 = 32'd3997
; 
32'd145839: dataIn1 = 32'd1977
; 
32'd145840: dataIn1 = 32'd2328
; 
32'd145841: dataIn1 = 32'd3044
; 
32'd145842: dataIn1 = 32'd3989
; 
32'd145843: dataIn1 = 32'd3998
; 
32'd145844: dataIn1 = 32'd3999
; 
32'd145845: dataIn1 = 32'd4000
; 
32'd145846: dataIn1 = 32'd2328
; 
32'd145847: dataIn1 = 32'd2329
; 
32'd145848: dataIn1 = 32'd3991
; 
32'd145849: dataIn1 = 32'd3998
; 
32'd145850: dataIn1 = 32'd3999
; 
32'd145851: dataIn1 = 32'd4000
; 
32'd145852: dataIn1 = 32'd4001
; 
32'd145853: dataIn1 = 32'd1977
; 
32'd145854: dataIn1 = 32'd2329
; 
32'd145855: dataIn1 = 32'd3047
; 
32'd145856: dataIn1 = 32'd3998
; 
32'd145857: dataIn1 = 32'd3999
; 
32'd145858: dataIn1 = 32'd4000
; 
32'd145859: dataIn1 = 32'd4009
; 
32'd145860: dataIn1 = 32'd453
; 
32'd145861: dataIn1 = 32'd2329
; 
32'd145862: dataIn1 = 32'd3991
; 
32'd145863: dataIn1 = 32'd3999
; 
32'd145864: dataIn1 = 32'd4001
; 
32'd145865: dataIn1 = 32'd4003
; 
32'd145866: dataIn1 = 32'd4007
; 
32'd145867: dataIn1 = 32'd2330
; 
32'd145868: dataIn1 = 32'd2331
; 
32'd145869: dataIn1 = 32'd4002
; 
32'd145870: dataIn1 = 32'd4003
; 
32'd145871: dataIn1 = 32'd4004
; 
32'd145872: dataIn1 = 32'd4005
; 
32'd145873: dataIn1 = 32'd4006
; 
32'd145874: dataIn1 = 32'd2329
; 
32'd145875: dataIn1 = 32'd2331
; 
32'd145876: dataIn1 = 32'd4001
; 
32'd145877: dataIn1 = 32'd4002
; 
32'd145878: dataIn1 = 32'd4003
; 
32'd145879: dataIn1 = 32'd4004
; 
32'd145880: dataIn1 = 32'd4007
; 
32'd145881: dataIn1 = 32'd2329
; 
32'd145882: dataIn1 = 32'd2330
; 
32'd145883: dataIn1 = 32'd4002
; 
32'd145884: dataIn1 = 32'd4003
; 
32'd145885: dataIn1 = 32'd4004
; 
32'd145886: dataIn1 = 32'd4008
; 
32'd145887: dataIn1 = 32'd4009
; 
32'd145888: dataIn1 = 32'd454
; 
32'd145889: dataIn1 = 32'd2331
; 
32'd145890: dataIn1 = 32'd4002
; 
32'd145891: dataIn1 = 32'd4005
; 
32'd145892: dataIn1 = 32'd4006
; 
32'd145893: dataIn1 = 32'd5327
; 
32'd145894: dataIn1 = 32'd454
; 
32'd145895: dataIn1 = 32'd2330
; 
32'd145896: dataIn1 = 32'd4002
; 
32'd145897: dataIn1 = 32'd4005
; 
32'd145898: dataIn1 = 32'd4006
; 
32'd145899: dataIn1 = 32'd4013
; 
32'd145900: dataIn1 = 32'd4023
; 
32'd145901: dataIn1 = 32'd453
; 
32'd145902: dataIn1 = 32'd2331
; 
32'd145903: dataIn1 = 32'd4001
; 
32'd145904: dataIn1 = 32'd4003
; 
32'd145905: dataIn1 = 32'd4007
; 
32'd145906: dataIn1 = 32'd5326
; 
32'd145907: dataIn1 = 32'd155
; 
32'd145908: dataIn1 = 32'd2330
; 
32'd145909: dataIn1 = 32'd3061
; 
32'd145910: dataIn1 = 32'd4004
; 
32'd145911: dataIn1 = 32'd4008
; 
32'd145912: dataIn1 = 32'd4009
; 
32'd145913: dataIn1 = 32'd4025
; 
32'd145914: dataIn1 = 32'd155
; 
32'd145915: dataIn1 = 32'd2329
; 
32'd145916: dataIn1 = 32'd3047
; 
32'd145917: dataIn1 = 32'd4000
; 
32'd145918: dataIn1 = 32'd4004
; 
32'd145919: dataIn1 = 32'd4008
; 
32'd145920: dataIn1 = 32'd4009
; 
32'd145921: dataIn1 = 32'd2333
; 
32'd145922: dataIn1 = 32'd2334
; 
32'd145923: dataIn1 = 32'd4010
; 
32'd145924: dataIn1 = 32'd4011
; 
32'd145925: dataIn1 = 32'd4012
; 
32'd145926: dataIn1 = 32'd4013
; 
32'd145927: dataIn1 = 32'd4014
; 
32'd145928: dataIn1 = 32'd2332
; 
32'd145929: dataIn1 = 32'd2334
; 
32'd145930: dataIn1 = 32'd4010
; 
32'd145931: dataIn1 = 32'd4011
; 
32'd145932: dataIn1 = 32'd4012
; 
32'd145933: dataIn1 = 32'd4015
; 
32'd145934: dataIn1 = 32'd4016
; 
32'd145935: dataIn1 = 32'd2332
; 
32'd145936: dataIn1 = 32'd2333
; 
32'd145937: dataIn1 = 32'd4010
; 
32'd145938: dataIn1 = 32'd4011
; 
32'd145939: dataIn1 = 32'd4012
; 
32'd145940: dataIn1 = 32'd4017
; 
32'd145941: dataIn1 = 32'd4018
; 
32'd145942: dataIn1 = 32'd454
; 
32'd145943: dataIn1 = 32'd2334
; 
32'd145944: dataIn1 = 32'd4006
; 
32'd145945: dataIn1 = 32'd4010
; 
32'd145946: dataIn1 = 32'd4013
; 
32'd145947: dataIn1 = 32'd4014
; 
32'd145948: dataIn1 = 32'd4023
; 
32'd145949: dataIn1 = 32'd454
; 
32'd145950: dataIn1 = 32'd2333
; 
32'd145951: dataIn1 = 32'd4010
; 
32'd145952: dataIn1 = 32'd4013
; 
32'd145953: dataIn1 = 32'd4014
; 
32'd145954: dataIn1 = 32'd5329
; 
32'd145955: dataIn1 = 32'd286
; 
32'd145956: dataIn1 = 32'd2334
; 
32'd145957: dataIn1 = 32'd3060
; 
32'd145958: dataIn1 = 32'd4011
; 
32'd145959: dataIn1 = 32'd4015
; 
32'd145960: dataIn1 = 32'd4016
; 
32'd145961: dataIn1 = 32'd4024
; 
32'd145962: dataIn1 = 32'd286
; 
32'd145963: dataIn1 = 32'd2332
; 
32'd145964: dataIn1 = 32'd3066
; 
32'd145965: dataIn1 = 32'd4011
; 
32'd145966: dataIn1 = 32'd4015
; 
32'd145967: dataIn1 = 32'd4016
; 
32'd145968: dataIn1 = 32'd4020
; 
32'd145969: dataIn1 = 32'd455
; 
32'd145970: dataIn1 = 32'd2333
; 
32'd145971: dataIn1 = 32'd4012
; 
32'd145972: dataIn1 = 32'd4017
; 
32'd145973: dataIn1 = 32'd4018
; 
32'd145974: dataIn1 = 32'd5328
; 
32'd145975: dataIn1 = 32'd455
; 
32'd145976: dataIn1 = 32'd2332
; 
32'd145977: dataIn1 = 32'd4012
; 
32'd145978: dataIn1 = 32'd4017
; 
32'd145979: dataIn1 = 32'd4018
; 
32'd145980: dataIn1 = 32'd4021
; 
32'd145981: dataIn1 = 32'd4022
; 
32'd145982: dataIn1 = 32'd1980
; 
32'd145983: dataIn1 = 32'd2335
; 
32'd145984: dataIn1 = 32'd3065
; 
32'd145985: dataIn1 = 32'd4019
; 
32'd145986: dataIn1 = 32'd4020
; 
32'd145987: dataIn1 = 32'd4021
; 
32'd145988: dataIn1 = 32'd4029
; 
32'd145989: dataIn1 = 32'd1980
; 
32'd145990: dataIn1 = 32'd2332
; 
32'd145991: dataIn1 = 32'd3066
; 
32'd145992: dataIn1 = 32'd4016
; 
32'd145993: dataIn1 = 32'd4019
; 
32'd145994: dataIn1 = 32'd4020
; 
32'd145995: dataIn1 = 32'd4021
; 
32'd145996: dataIn1 = 32'd2332
; 
32'd145997: dataIn1 = 32'd2335
; 
32'd145998: dataIn1 = 32'd4018
; 
32'd145999: dataIn1 = 32'd4019
; 
32'd146000: dataIn1 = 32'd4020
; 
32'd146001: dataIn1 = 32'd4021
; 
32'd146002: dataIn1 = 32'd4022
; 
32'd146003: dataIn1 = 32'd455
; 
32'd146004: dataIn1 = 32'd2335
; 
32'd146005: dataIn1 = 32'd4018
; 
32'd146006: dataIn1 = 32'd4021
; 
32'd146007: dataIn1 = 32'd4022
; 
32'd146008: dataIn1 = 32'd4027
; 
32'd146009: dataIn1 = 32'd4031
; 
32'd146010: dataIn1 = 32'd2330
; 
32'd146011: dataIn1 = 32'd2334
; 
32'd146012: dataIn1 = 32'd4006
; 
32'd146013: dataIn1 = 32'd4013
; 
32'd146014: dataIn1 = 32'd4023
; 
32'd146015: dataIn1 = 32'd4024
; 
32'd146016: dataIn1 = 32'd4025
; 
32'd146017: dataIn1 = 32'd1979
; 
32'd146018: dataIn1 = 32'd2334
; 
32'd146019: dataIn1 = 32'd3060
; 
32'd146020: dataIn1 = 32'd4015
; 
32'd146021: dataIn1 = 32'd4023
; 
32'd146022: dataIn1 = 32'd4024
; 
32'd146023: dataIn1 = 32'd4025
; 
32'd146024: dataIn1 = 32'd1979
; 
32'd146025: dataIn1 = 32'd2330
; 
32'd146026: dataIn1 = 32'd3061
; 
32'd146027: dataIn1 = 32'd4008
; 
32'd146028: dataIn1 = 32'd4023
; 
32'd146029: dataIn1 = 32'd4024
; 
32'd146030: dataIn1 = 32'd4025
; 
32'd146031: dataIn1 = 32'd2335
; 
32'd146032: dataIn1 = 32'd2337
; 
32'd146033: dataIn1 = 32'd4026
; 
32'd146034: dataIn1 = 32'd4027
; 
32'd146035: dataIn1 = 32'd4028
; 
32'd146036: dataIn1 = 32'd4029
; 
32'd146037: dataIn1 = 32'd4030
; 
32'd146038: dataIn1 = 32'd2335
; 
32'd146039: dataIn1 = 32'd2336
; 
32'd146040: dataIn1 = 32'd4022
; 
32'd146041: dataIn1 = 32'd4026
; 
32'd146042: dataIn1 = 32'd4027
; 
32'd146043: dataIn1 = 32'd4028
; 
32'd146044: dataIn1 = 32'd4031
; 
32'd146045: dataIn1 = 32'd2336
; 
32'd146046: dataIn1 = 32'd2337
; 
32'd146047: dataIn1 = 32'd4026
; 
32'd146048: dataIn1 = 32'd4027
; 
32'd146049: dataIn1 = 32'd4028
; 
32'd146050: dataIn1 = 32'd4032
; 
32'd146051: dataIn1 = 32'd4033
; 
32'd146052: dataIn1 = 32'd157
; 
32'd146053: dataIn1 = 32'd2335
; 
32'd146054: dataIn1 = 32'd3065
; 
32'd146055: dataIn1 = 32'd4019
; 
32'd146056: dataIn1 = 32'd4026
; 
32'd146057: dataIn1 = 32'd4029
; 
32'd146058: dataIn1 = 32'd4030
; 
32'd146059: dataIn1 = 32'd157
; 
32'd146060: dataIn1 = 32'd2337
; 
32'd146061: dataIn1 = 32'd3072
; 
32'd146062: dataIn1 = 32'd4026
; 
32'd146063: dataIn1 = 32'd4029
; 
32'd146064: dataIn1 = 32'd4030
; 
32'd146065: dataIn1 = 32'd4043
; 
32'd146066: dataIn1 = 32'd455
; 
32'd146067: dataIn1 = 32'd2336
; 
32'd146068: dataIn1 = 32'd4022
; 
32'd146069: dataIn1 = 32'd4027
; 
32'd146070: dataIn1 = 32'd4031
; 
32'd146071: dataIn1 = 32'd5331
; 
32'd146072: dataIn1 = 32'd456
; 
32'd146073: dataIn1 = 32'd2337
; 
32'd146074: dataIn1 = 32'd4028
; 
32'd146075: dataIn1 = 32'd4032
; 
32'd146076: dataIn1 = 32'd4033
; 
32'd146077: dataIn1 = 32'd4042
; 
32'd146078: dataIn1 = 32'd4045
; 
32'd146079: dataIn1 = 32'd456
; 
32'd146080: dataIn1 = 32'd2336
; 
32'd146081: dataIn1 = 32'd4028
; 
32'd146082: dataIn1 = 32'd4032
; 
32'd146083: dataIn1 = 32'd4033
; 
32'd146084: dataIn1 = 32'd5330
; 
32'd146085: dataIn1 = 32'd2339
; 
32'd146086: dataIn1 = 32'd2340
; 
32'd146087: dataIn1 = 32'd4034
; 
32'd146088: dataIn1 = 32'd4035
; 
32'd146089: dataIn1 = 32'd4036
; 
32'd146090: dataIn1 = 32'd4037
; 
32'd146091: dataIn1 = 32'd4038
; 
32'd146092: dataIn1 = 32'd2338
; 
32'd146093: dataIn1 = 32'd2340
; 
32'd146094: dataIn1 = 32'd4034
; 
32'd146095: dataIn1 = 32'd4035
; 
32'd146096: dataIn1 = 32'd4036
; 
32'd146097: dataIn1 = 32'd4039
; 
32'd146098: dataIn1 = 32'd4040
; 
32'd146099: dataIn1 = 32'd2338
; 
32'd146100: dataIn1 = 32'd2339
; 
32'd146101: dataIn1 = 32'd4034
; 
32'd146102: dataIn1 = 32'd4035
; 
32'd146103: dataIn1 = 32'd4036
; 
32'd146104: dataIn1 = 32'd4041
; 
32'd146105: dataIn1 = 32'd4042
; 
32'd146106: dataIn1 = 32'd457
; 
32'd146107: dataIn1 = 32'd2340
; 
32'd146108: dataIn1 = 32'd4034
; 
32'd146109: dataIn1 = 32'd4037
; 
32'd146110: dataIn1 = 32'd4038
; 
32'd146111: dataIn1 = 32'd4046
; 
32'd146112: dataIn1 = 32'd4049
; 
32'd146113: dataIn1 = 32'd457
; 
32'd146114: dataIn1 = 32'd2339
; 
32'd146115: dataIn1 = 32'd4034
; 
32'd146116: dataIn1 = 32'd4037
; 
32'd146117: dataIn1 = 32'd4038
; 
32'd146118: dataIn1 = 32'd5333
; 
32'd146119: dataIn1 = 32'd293
; 
32'd146120: dataIn1 = 32'd2340
; 
32'd146121: dataIn1 = 32'd3081
; 
32'd146122: dataIn1 = 32'd4035
; 
32'd146123: dataIn1 = 32'd4039
; 
32'd146124: dataIn1 = 32'd4040
; 
32'd146125: dataIn1 = 32'd4047
; 
32'd146126: dataIn1 = 32'd293
; 
32'd146127: dataIn1 = 32'd2338
; 
32'd146128: dataIn1 = 32'd3073
; 
32'd146129: dataIn1 = 32'd4035
; 
32'd146130: dataIn1 = 32'd4039
; 
32'd146131: dataIn1 = 32'd4040
; 
32'd146132: dataIn1 = 32'd4044
; 
32'd146133: dataIn1 = 32'd456
; 
32'd146134: dataIn1 = 32'd2339
; 
32'd146135: dataIn1 = 32'd4036
; 
32'd146136: dataIn1 = 32'd4041
; 
32'd146137: dataIn1 = 32'd4042
; 
32'd146138: dataIn1 = 32'd5332
; 
32'd146139: dataIn1 = 32'd456
; 
32'd146140: dataIn1 = 32'd2338
; 
32'd146141: dataIn1 = 32'd4032
; 
32'd146142: dataIn1 = 32'd4036
; 
32'd146143: dataIn1 = 32'd4041
; 
32'd146144: dataIn1 = 32'd4042
; 
32'd146145: dataIn1 = 32'd4045
; 
32'd146146: dataIn1 = 32'd1981
; 
32'd146147: dataIn1 = 32'd2337
; 
32'd146148: dataIn1 = 32'd3072
; 
32'd146149: dataIn1 = 32'd4030
; 
32'd146150: dataIn1 = 32'd4043
; 
32'd146151: dataIn1 = 32'd4044
; 
32'd146152: dataIn1 = 32'd4045
; 
32'd146153: dataIn1 = 32'd1981
; 
32'd146154: dataIn1 = 32'd2338
; 
32'd146155: dataIn1 = 32'd3073
; 
32'd146156: dataIn1 = 32'd4040
; 
32'd146157: dataIn1 = 32'd4043
; 
32'd146158: dataIn1 = 32'd4044
; 
32'd146159: dataIn1 = 32'd4045
; 
32'd146160: dataIn1 = 32'd2337
; 
32'd146161: dataIn1 = 32'd2338
; 
32'd146162: dataIn1 = 32'd4032
; 
32'd146163: dataIn1 = 32'd4042
; 
32'd146164: dataIn1 = 32'd4043
; 
32'd146165: dataIn1 = 32'd4044
; 
32'd146166: dataIn1 = 32'd4045
; 
32'd146167: dataIn1 = 32'd2340
; 
32'd146168: dataIn1 = 32'd2341
; 
32'd146169: dataIn1 = 32'd4037
; 
32'd146170: dataIn1 = 32'd4046
; 
32'd146171: dataIn1 = 32'd4047
; 
32'd146172: dataIn1 = 32'd4048
; 
32'd146173: dataIn1 = 32'd4049
; 
32'd146174: dataIn1 = 32'd1982
; 
32'd146175: dataIn1 = 32'd2340
; 
32'd146176: dataIn1 = 32'd3081
; 
32'd146177: dataIn1 = 32'd4039
; 
32'd146178: dataIn1 = 32'd4046
; 
32'd146179: dataIn1 = 32'd4047
; 
32'd146180: dataIn1 = 32'd4048
; 
32'd146181: dataIn1 = 32'd1982
; 
32'd146182: dataIn1 = 32'd2341
; 
32'd146183: dataIn1 = 32'd3082
; 
32'd146184: dataIn1 = 32'd4046
; 
32'd146185: dataIn1 = 32'd4047
; 
32'd146186: dataIn1 = 32'd4048
; 
32'd146187: dataIn1 = 32'd4056
; 
32'd146188: dataIn1 = 32'd457
; 
32'd146189: dataIn1 = 32'd2341
; 
32'd146190: dataIn1 = 32'd4037
; 
32'd146191: dataIn1 = 32'd4046
; 
32'd146192: dataIn1 = 32'd4049
; 
32'd146193: dataIn1 = 32'd4050
; 
32'd146194: dataIn1 = 32'd4053
; 
32'd146195: dataIn1 = 32'd2341
; 
32'd146196: dataIn1 = 32'd2343
; 
32'd146197: dataIn1 = 32'd4049
; 
32'd146198: dataIn1 = 32'd4050
; 
32'd146199: dataIn1 = 32'd4051
; 
32'd146200: dataIn1 = 32'd4052
; 
32'd146201: dataIn1 = 32'd4053
; 
32'd146202: dataIn1 = 32'd2342
; 
32'd146203: dataIn1 = 32'd2343
; 
32'd146204: dataIn1 = 32'd4050
; 
32'd146205: dataIn1 = 32'd4051
; 
32'd146206: dataIn1 = 32'd4052
; 
32'd146207: dataIn1 = 32'd4054
; 
32'd146208: dataIn1 = 32'd4055
; 
32'd146209: dataIn1 = 32'd2341
; 
32'd146210: dataIn1 = 32'd2342
; 
32'd146211: dataIn1 = 32'd4050
; 
32'd146212: dataIn1 = 32'd4051
; 
32'd146213: dataIn1 = 32'd4052
; 
32'd146214: dataIn1 = 32'd4056
; 
32'd146215: dataIn1 = 32'd4057
; 
32'd146216: dataIn1 = 32'd457
; 
32'd146217: dataIn1 = 32'd2343
; 
32'd146218: dataIn1 = 32'd4049
; 
32'd146219: dataIn1 = 32'd4050
; 
32'd146220: dataIn1 = 32'd4053
; 
32'd146221: dataIn1 = 32'd5335
; 
32'd146222: dataIn1 = 32'd458
; 
32'd146223: dataIn1 = 32'd2343
; 
32'd146224: dataIn1 = 32'd4051
; 
32'd146225: dataIn1 = 32'd4054
; 
32'd146226: dataIn1 = 32'd4055
; 
32'd146227: dataIn1 = 32'd5334
; 
32'd146228: dataIn1 = 32'd458
; 
32'd146229: dataIn1 = 32'd2342
; 
32'd146230: dataIn1 = 32'd4051
; 
32'd146231: dataIn1 = 32'd4054
; 
32'd146232: dataIn1 = 32'd4055
; 
32'd146233: dataIn1 = 32'd4064
; 
32'd146234: dataIn1 = 32'd4068
; 
32'd146235: dataIn1 = 32'd159
; 
32'd146236: dataIn1 = 32'd2341
; 
32'd146237: dataIn1 = 32'd3082
; 
32'd146238: dataIn1 = 32'd4048
; 
32'd146239: dataIn1 = 32'd4052
; 
32'd146240: dataIn1 = 32'd4056
; 
32'd146241: dataIn1 = 32'd4057
; 
32'd146242: dataIn1 = 32'd159
; 
32'd146243: dataIn1 = 32'd2342
; 
32'd146244: dataIn1 = 32'd3107
; 
32'd146245: dataIn1 = 32'd4052
; 
32'd146246: dataIn1 = 32'd4056
; 
32'd146247: dataIn1 = 32'd4057
; 
32'd146248: dataIn1 = 32'd4067
; 
32'd146249: dataIn1 = 32'd2345
; 
32'd146250: dataIn1 = 32'd2346
; 
32'd146251: dataIn1 = 32'd4058
; 
32'd146252: dataIn1 = 32'd4059
; 
32'd146253: dataIn1 = 32'd4060
; 
32'd146254: dataIn1 = 32'd4061
; 
32'd146255: dataIn1 = 32'd4062
; 
32'd146256: dataIn1 = 32'd2344
; 
32'd146257: dataIn1 = 32'd2346
; 
32'd146258: dataIn1 = 32'd4058
; 
32'd146259: dataIn1 = 32'd4059
; 
32'd146260: dataIn1 = 32'd4060
; 
32'd146261: dataIn1 = 32'd4063
; 
32'd146262: dataIn1 = 32'd4064
; 
32'd146263: dataIn1 = 32'd2344
; 
32'd146264: dataIn1 = 32'd2345
; 
32'd146265: dataIn1 = 32'd4058
; 
32'd146266: dataIn1 = 32'd4059
; 
32'd146267: dataIn1 = 32'd4060
; 
32'd146268: dataIn1 = 32'd4065
; 
32'd146269: dataIn1 = 32'd4066
; 
32'd146270: dataIn1 = 32'd459
; 
32'd146271: dataIn1 = 32'd2346
; 
32'd146272: dataIn1 = 32'd4058
; 
32'd146273: dataIn1 = 32'd4061
; 
32'd146274: dataIn1 = 32'd4062
; 
32'd146275: dataIn1 = 32'd5337
; 
32'd146276: dataIn1 = 32'd459
; 
32'd146277: dataIn1 = 32'd2345
; 
32'd146278: dataIn1 = 32'd4058
; 
32'd146279: dataIn1 = 32'd4061
; 
32'd146280: dataIn1 = 32'd4062
; 
32'd146281: dataIn1 = 32'd4070
; 
32'd146282: dataIn1 = 32'd4073
; 
32'd146283: dataIn1 = 32'd458
; 
32'd146284: dataIn1 = 32'd2346
; 
32'd146285: dataIn1 = 32'd4059
; 
32'd146286: dataIn1 = 32'd4063
; 
32'd146287: dataIn1 = 32'd4064
; 
32'd146288: dataIn1 = 32'd5336
; 
32'd146289: dataIn1 = 32'd458
; 
32'd146290: dataIn1 = 32'd2344
; 
32'd146291: dataIn1 = 32'd4055
; 
32'd146292: dataIn1 = 32'd4059
; 
32'd146293: dataIn1 = 32'd4063
; 
32'd146294: dataIn1 = 32'd4064
; 
32'd146295: dataIn1 = 32'd4068
; 
32'd146296: dataIn1 = 32'd301
; 
32'd146297: dataIn1 = 32'd2345
; 
32'd146298: dataIn1 = 32'd3103
; 
32'd146299: dataIn1 = 32'd4060
; 
32'd146300: dataIn1 = 32'd4065
; 
32'd146301: dataIn1 = 32'd4066
; 
32'd146302: dataIn1 = 32'd4072
; 
32'd146303: dataIn1 = 32'd301
; 
32'd146304: dataIn1 = 32'd2344
; 
32'd146305: dataIn1 = 32'd3110
; 
32'd146306: dataIn1 = 32'd4060
; 
32'd146307: dataIn1 = 32'd4065
; 
32'd146308: dataIn1 = 32'd4066
; 
32'd146309: dataIn1 = 32'd4069
; 
32'd146310: dataIn1 = 32'd1986
; 
32'd146311: dataIn1 = 32'd2342
; 
32'd146312: dataIn1 = 32'd3107
; 
32'd146313: dataIn1 = 32'd4057
; 
32'd146314: dataIn1 = 32'd4067
; 
32'd146315: dataIn1 = 32'd4068
; 
32'd146316: dataIn1 = 32'd4069
; 
32'd146317: dataIn1 = 32'd2342
; 
32'd146318: dataIn1 = 32'd2344
; 
32'd146319: dataIn1 = 32'd4055
; 
32'd146320: dataIn1 = 32'd4064
; 
32'd146321: dataIn1 = 32'd4067
; 
32'd146322: dataIn1 = 32'd4068
; 
32'd146323: dataIn1 = 32'd4069
; 
32'd146324: dataIn1 = 32'd1986
; 
32'd146325: dataIn1 = 32'd2344
; 
32'd146326: dataIn1 = 32'd3110
; 
32'd146327: dataIn1 = 32'd4066
; 
32'd146328: dataIn1 = 32'd4067
; 
32'd146329: dataIn1 = 32'd4068
; 
32'd146330: dataIn1 = 32'd4069
; 
32'd146331: dataIn1 = 32'd2345
; 
32'd146332: dataIn1 = 32'd2347
; 
32'd146333: dataIn1 = 32'd4062
; 
32'd146334: dataIn1 = 32'd4070
; 
32'd146335: dataIn1 = 32'd4071
; 
32'd146336: dataIn1 = 32'd4072
; 
32'd146337: dataIn1 = 32'd4073
; 
32'd146338: dataIn1 = 32'd1985
; 
32'd146339: dataIn1 = 32'd2347
; 
32'd146340: dataIn1 = 32'd3102
; 
32'd146341: dataIn1 = 32'd4070
; 
32'd146342: dataIn1 = 32'd4071
; 
32'd146343: dataIn1 = 32'd4072
; 
32'd146344: dataIn1 = 32'd4078
; 
32'd146345: dataIn1 = 32'd1985
; 
32'd146346: dataIn1 = 32'd2345
; 
32'd146347: dataIn1 = 32'd3103
; 
32'd146348: dataIn1 = 32'd4065
; 
32'd146349: dataIn1 = 32'd4070
; 
32'd146350: dataIn1 = 32'd4071
; 
32'd146351: dataIn1 = 32'd4072
; 
32'd146352: dataIn1 = 32'd459
; 
32'd146353: dataIn1 = 32'd2347
; 
32'd146354: dataIn1 = 32'd4062
; 
32'd146355: dataIn1 = 32'd4070
; 
32'd146356: dataIn1 = 32'd4073
; 
32'd146357: dataIn1 = 32'd4074
; 
32'd146358: dataIn1 = 32'd4077
; 
32'd146359: dataIn1 = 32'd2347
; 
32'd146360: dataIn1 = 32'd2349
; 
32'd146361: dataIn1 = 32'd4073
; 
32'd146362: dataIn1 = 32'd4074
; 
32'd146363: dataIn1 = 32'd4075
; 
32'd146364: dataIn1 = 32'd4076
; 
32'd146365: dataIn1 = 32'd4077
; 
32'd146366: dataIn1 = 32'd2347
; 
32'd146367: dataIn1 = 32'd2348
; 
32'd146368: dataIn1 = 32'd4074
; 
32'd146369: dataIn1 = 32'd4075
; 
32'd146370: dataIn1 = 32'd4076
; 
32'd146371: dataIn1 = 32'd4078
; 
32'd146372: dataIn1 = 32'd4079
; 
32'd146373: dataIn1 = 32'd2348
; 
32'd146374: dataIn1 = 32'd2349
; 
32'd146375: dataIn1 = 32'd4074
; 
32'd146376: dataIn1 = 32'd4075
; 
32'd146377: dataIn1 = 32'd4076
; 
32'd146378: dataIn1 = 32'd4080
; 
32'd146379: dataIn1 = 32'd4081
; 
32'd146380: dataIn1 = 32'd459
; 
32'd146381: dataIn1 = 32'd2349
; 
32'd146382: dataIn1 = 32'd4073
; 
32'd146383: dataIn1 = 32'd4074
; 
32'd146384: dataIn1 = 32'd4077
; 
32'd146385: dataIn1 = 32'd5339
; 
32'd146386: dataIn1 = 32'd161
; 
32'd146387: dataIn1 = 32'd2347
; 
32'd146388: dataIn1 = 32'd3102
; 
32'd146389: dataIn1 = 32'd4071
; 
32'd146390: dataIn1 = 32'd4075
; 
32'd146391: dataIn1 = 32'd4078
; 
32'd146392: dataIn1 = 32'd4079
; 
32'd146393: dataIn1 = 32'd161
; 
32'd146394: dataIn1 = 32'd2348
; 
32'd146395: dataIn1 = 32'd3094
; 
32'd146396: dataIn1 = 32'd4075
; 
32'd146397: dataIn1 = 32'd4078
; 
32'd146398: dataIn1 = 32'd4079
; 
32'd146399: dataIn1 = 32'd4092
; 
32'd146400: dataIn1 = 32'd460
; 
32'd146401: dataIn1 = 32'd2349
; 
32'd146402: dataIn1 = 32'd4076
; 
32'd146403: dataIn1 = 32'd4080
; 
32'd146404: dataIn1 = 32'd4081
; 
32'd146405: dataIn1 = 32'd5338
; 
32'd146406: dataIn1 = 32'd460
; 
32'd146407: dataIn1 = 32'd2348
; 
32'd146408: dataIn1 = 32'd4076
; 
32'd146409: dataIn1 = 32'd4080
; 
32'd146410: dataIn1 = 32'd4081
; 
32'd146411: dataIn1 = 32'd4089
; 
32'd146412: dataIn1 = 32'd4093
; 
32'd146413: dataIn1 = 32'd2351
; 
32'd146414: dataIn1 = 32'd2352
; 
32'd146415: dataIn1 = 32'd4082
; 
32'd146416: dataIn1 = 32'd4083
; 
32'd146417: dataIn1 = 32'd4084
; 
32'd146418: dataIn1 = 32'd4085
; 
32'd146419: dataIn1 = 32'd4086
; 
32'd146420: dataIn1 = 32'd2350
; 
32'd146421: dataIn1 = 32'd2352
; 
32'd146422: dataIn1 = 32'd4082
; 
32'd146423: dataIn1 = 32'd4083
; 
32'd146424: dataIn1 = 32'd4084
; 
32'd146425: dataIn1 = 32'd4087
; 
32'd146426: dataIn1 = 32'd4088
; 
32'd146427: dataIn1 = 32'd2350
; 
32'd146428: dataIn1 = 32'd2351
; 
32'd146429: dataIn1 = 32'd4082
; 
32'd146430: dataIn1 = 32'd4083
; 
32'd146431: dataIn1 = 32'd4084
; 
32'd146432: dataIn1 = 32'd4089
; 
32'd146433: dataIn1 = 32'd4090
; 
32'd146434: dataIn1 = 32'd295
; 
32'd146435: dataIn1 = 32'd2352
; 
32'd146436: dataIn1 = 32'd3086
; 
32'd146437: dataIn1 = 32'd4082
; 
32'd146438: dataIn1 = 32'd4085
; 
32'd146439: dataIn1 = 32'd4086
; 
32'd146440: dataIn1 = 32'd4094
; 
32'd146441: dataIn1 = 32'd295
; 
32'd146442: dataIn1 = 32'd2351
; 
32'd146443: dataIn1 = 32'd3093
; 
32'd146444: dataIn1 = 32'd4082
; 
32'd146445: dataIn1 = 32'd4085
; 
32'd146446: dataIn1 = 32'd4086
; 
32'd146447: dataIn1 = 32'd4091
; 
32'd146448: dataIn1 = 32'd461
; 
32'd146449: dataIn1 = 32'd2352
; 
32'd146450: dataIn1 = 32'd4083
; 
32'd146451: dataIn1 = 32'd4087
; 
32'd146452: dataIn1 = 32'd4088
; 
32'd146453: dataIn1 = 32'd4095
; 
32'd146454: dataIn1 = 32'd4097
; 
32'd146455: dataIn1 = 32'd461
; 
32'd146456: dataIn1 = 32'd2350
; 
32'd146457: dataIn1 = 32'd4083
; 
32'd146458: dataIn1 = 32'd4087
; 
32'd146459: dataIn1 = 32'd4088
; 
32'd146460: dataIn1 = 32'd5341
; 
32'd146461: dataIn1 = 32'd460
; 
32'd146462: dataIn1 = 32'd2351
; 
32'd146463: dataIn1 = 32'd4081
; 
32'd146464: dataIn1 = 32'd4084
; 
32'd146465: dataIn1 = 32'd4089
; 
32'd146466: dataIn1 = 32'd4090
; 
32'd146467: dataIn1 = 32'd4093
; 
32'd146468: dataIn1 = 32'd460
; 
32'd146469: dataIn1 = 32'd2350
; 
32'd146470: dataIn1 = 32'd4084
; 
32'd146471: dataIn1 = 32'd4089
; 
32'd146472: dataIn1 = 32'd4090
; 
32'd146473: dataIn1 = 32'd5340
; 
32'd146474: dataIn1 = 32'd1984
; 
32'd146475: dataIn1 = 32'd2351
; 
32'd146476: dataIn1 = 32'd3093
; 
32'd146477: dataIn1 = 32'd4086
; 
32'd146478: dataIn1 = 32'd4091
; 
32'd146479: dataIn1 = 32'd4092
; 
32'd146480: dataIn1 = 32'd4093
; 
32'd146481: dataIn1 = 32'd1984
; 
32'd146482: dataIn1 = 32'd2348
; 
32'd146483: dataIn1 = 32'd3094
; 
32'd146484: dataIn1 = 32'd4079
; 
32'd146485: dataIn1 = 32'd4091
; 
32'd146486: dataIn1 = 32'd4092
; 
32'd146487: dataIn1 = 32'd4093
; 
32'd146488: dataIn1 = 32'd2348
; 
32'd146489: dataIn1 = 32'd2351
; 
32'd146490: dataIn1 = 32'd4081
; 
32'd146491: dataIn1 = 32'd4089
; 
32'd146492: dataIn1 = 32'd4091
; 
32'd146493: dataIn1 = 32'd4092
; 
32'd146494: dataIn1 = 32'd4093
; 
32'd146495: dataIn1 = 32'd1983
; 
32'd146496: dataIn1 = 32'd2352
; 
32'd146497: dataIn1 = 32'd3086
; 
32'd146498: dataIn1 = 32'd4085
; 
32'd146499: dataIn1 = 32'd4094
; 
32'd146500: dataIn1 = 32'd4095
; 
32'd146501: dataIn1 = 32'd4096
; 
32'd146502: dataIn1 = 32'd2352
; 
32'd146503: dataIn1 = 32'd2353
; 
32'd146504: dataIn1 = 32'd4087
; 
32'd146505: dataIn1 = 32'd4094
; 
32'd146506: dataIn1 = 32'd4095
; 
32'd146507: dataIn1 = 32'd4096
; 
32'd146508: dataIn1 = 32'd4097
; 
32'd146509: dataIn1 = 32'd1983
; 
32'd146510: dataIn1 = 32'd2353
; 
32'd146511: dataIn1 = 32'd3089
; 
32'd146512: dataIn1 = 32'd4094
; 
32'd146513: dataIn1 = 32'd4095
; 
32'd146514: dataIn1 = 32'd4096
; 
32'd146515: dataIn1 = 32'd4105
; 
32'd146516: dataIn1 = 32'd461
; 
32'd146517: dataIn1 = 32'd2353
; 
32'd146518: dataIn1 = 32'd4087
; 
32'd146519: dataIn1 = 32'd4095
; 
32'd146520: dataIn1 = 32'd4097
; 
32'd146521: dataIn1 = 32'd4099
; 
32'd146522: dataIn1 = 32'd4103
; 
32'd146523: dataIn1 = 32'd2354
; 
32'd146524: dataIn1 = 32'd2355
; 
32'd146525: dataIn1 = 32'd4098
; 
32'd146526: dataIn1 = 32'd4099
; 
32'd146527: dataIn1 = 32'd4100
; 
32'd146528: dataIn1 = 32'd4101
; 
32'd146529: dataIn1 = 32'd4102
; 
32'd146530: dataIn1 = 32'd2353
; 
32'd146531: dataIn1 = 32'd2355
; 
32'd146532: dataIn1 = 32'd4097
; 
32'd146533: dataIn1 = 32'd4098
; 
32'd146534: dataIn1 = 32'd4099
; 
32'd146535: dataIn1 = 32'd4100
; 
32'd146536: dataIn1 = 32'd4103
; 
32'd146537: dataIn1 = 32'd2353
; 
32'd146538: dataIn1 = 32'd2354
; 
32'd146539: dataIn1 = 32'd4098
; 
32'd146540: dataIn1 = 32'd4099
; 
32'd146541: dataIn1 = 32'd4100
; 
32'd146542: dataIn1 = 32'd4104
; 
32'd146543: dataIn1 = 32'd4105
; 
32'd146544: dataIn1 = 32'd462
; 
32'd146545: dataIn1 = 32'd2355
; 
32'd146546: dataIn1 = 32'd4098
; 
32'd146547: dataIn1 = 32'd4101
; 
32'd146548: dataIn1 = 32'd4102
; 
32'd146549: dataIn1 = 32'd5343
; 
32'd146550: dataIn1 = 32'd462
; 
32'd146551: dataIn1 = 32'd2354
; 
32'd146552: dataIn1 = 32'd4098
; 
32'd146553: dataIn1 = 32'd4101
; 
32'd146554: dataIn1 = 32'd4102
; 
32'd146555: dataIn1 = 32'd4109
; 
32'd146556: dataIn1 = 32'd4119
; 
32'd146557: dataIn1 = 32'd461
; 
32'd146558: dataIn1 = 32'd2355
; 
32'd146559: dataIn1 = 32'd4097
; 
32'd146560: dataIn1 = 32'd4099
; 
32'd146561: dataIn1 = 32'd4103
; 
32'd146562: dataIn1 = 32'd5342
; 
32'd146563: dataIn1 = 32'd162
; 
32'd146564: dataIn1 = 32'd2354
; 
32'd146565: dataIn1 = 32'd3117
; 
32'd146566: dataIn1 = 32'd4100
; 
32'd146567: dataIn1 = 32'd4104
; 
32'd146568: dataIn1 = 32'd4105
; 
32'd146569: dataIn1 = 32'd4121
; 
32'd146570: dataIn1 = 32'd162
; 
32'd146571: dataIn1 = 32'd2353
; 
32'd146572: dataIn1 = 32'd3089
; 
32'd146573: dataIn1 = 32'd4096
; 
32'd146574: dataIn1 = 32'd4100
; 
32'd146575: dataIn1 = 32'd4104
; 
32'd146576: dataIn1 = 32'd4105
; 
32'd146577: dataIn1 = 32'd2357
; 
32'd146578: dataIn1 = 32'd2358
; 
32'd146579: dataIn1 = 32'd4106
; 
32'd146580: dataIn1 = 32'd4107
; 
32'd146581: dataIn1 = 32'd4108
; 
32'd146582: dataIn1 = 32'd4109
; 
32'd146583: dataIn1 = 32'd4110
; 
32'd146584: dataIn1 = 32'd2356
; 
32'd146585: dataIn1 = 32'd2358
; 
32'd146586: dataIn1 = 32'd4106
; 
32'd146587: dataIn1 = 32'd4107
; 
32'd146588: dataIn1 = 32'd4108
; 
32'd146589: dataIn1 = 32'd4111
; 
32'd146590: dataIn1 = 32'd4112
; 
32'd146591: dataIn1 = 32'd2356
; 
32'd146592: dataIn1 = 32'd2357
; 
32'd146593: dataIn1 = 32'd4106
; 
32'd146594: dataIn1 = 32'd4107
; 
32'd146595: dataIn1 = 32'd4108
; 
32'd146596: dataIn1 = 32'd4113
; 
32'd146597: dataIn1 = 32'd4114
; 
32'd146598: dataIn1 = 32'd462
; 
32'd146599: dataIn1 = 32'd2358
; 
32'd146600: dataIn1 = 32'd4102
; 
32'd146601: dataIn1 = 32'd4106
; 
32'd146602: dataIn1 = 32'd4109
; 
32'd146603: dataIn1 = 32'd4110
; 
32'd146604: dataIn1 = 32'd4119
; 
32'd146605: dataIn1 = 32'd462
; 
32'd146606: dataIn1 = 32'd2357
; 
32'd146607: dataIn1 = 32'd4106
; 
32'd146608: dataIn1 = 32'd4109
; 
32'd146609: dataIn1 = 32'd4110
; 
32'd146610: dataIn1 = 32'd5345
; 
32'd146611: dataIn1 = 32'd302
; 
32'd146612: dataIn1 = 32'd2358
; 
32'd146613: dataIn1 = 32'd3116
; 
32'd146614: dataIn1 = 32'd4107
; 
32'd146615: dataIn1 = 32'd4111
; 
32'd146616: dataIn1 = 32'd4112
; 
32'd146617: dataIn1 = 32'd4120
; 
32'd146618: dataIn1 = 32'd302
; 
32'd146619: dataIn1 = 32'd2356
; 
32'd146620: dataIn1 = 32'd3122
; 
32'd146621: dataIn1 = 32'd4107
; 
32'd146622: dataIn1 = 32'd4111
; 
32'd146623: dataIn1 = 32'd4112
; 
32'd146624: dataIn1 = 32'd4116
; 
32'd146625: dataIn1 = 32'd463
; 
32'd146626: dataIn1 = 32'd2357
; 
32'd146627: dataIn1 = 32'd4108
; 
32'd146628: dataIn1 = 32'd4113
; 
32'd146629: dataIn1 = 32'd4114
; 
32'd146630: dataIn1 = 32'd5344
; 
32'd146631: dataIn1 = 32'd463
; 
32'd146632: dataIn1 = 32'd2356
; 
32'd146633: dataIn1 = 32'd4108
; 
32'd146634: dataIn1 = 32'd4113
; 
32'd146635: dataIn1 = 32'd4114
; 
32'd146636: dataIn1 = 32'd4117
; 
32'd146637: dataIn1 = 32'd4118
; 
32'd146638: dataIn1 = 32'd1988
; 
32'd146639: dataIn1 = 32'd2359
; 
32'd146640: dataIn1 = 32'd3121
; 
32'd146641: dataIn1 = 32'd4115
; 
32'd146642: dataIn1 = 32'd4116
; 
32'd146643: dataIn1 = 32'd4117
; 
32'd146644: dataIn1 = 32'd4125
; 
32'd146645: dataIn1 = 32'd1988
; 
32'd146646: dataIn1 = 32'd2356
; 
32'd146647: dataIn1 = 32'd3122
; 
32'd146648: dataIn1 = 32'd4112
; 
32'd146649: dataIn1 = 32'd4115
; 
32'd146650: dataIn1 = 32'd4116
; 
32'd146651: dataIn1 = 32'd4117
; 
32'd146652: dataIn1 = 32'd2356
; 
32'd146653: dataIn1 = 32'd2359
; 
32'd146654: dataIn1 = 32'd4114
; 
32'd146655: dataIn1 = 32'd4115
; 
32'd146656: dataIn1 = 32'd4116
; 
32'd146657: dataIn1 = 32'd4117
; 
32'd146658: dataIn1 = 32'd4118
; 
32'd146659: dataIn1 = 32'd463
; 
32'd146660: dataIn1 = 32'd2359
; 
32'd146661: dataIn1 = 32'd4114
; 
32'd146662: dataIn1 = 32'd4117
; 
32'd146663: dataIn1 = 32'd4118
; 
32'd146664: dataIn1 = 32'd4123
; 
32'd146665: dataIn1 = 32'd4127
; 
32'd146666: dataIn1 = 32'd2354
; 
32'd146667: dataIn1 = 32'd2358
; 
32'd146668: dataIn1 = 32'd4102
; 
32'd146669: dataIn1 = 32'd4109
; 
32'd146670: dataIn1 = 32'd4119
; 
32'd146671: dataIn1 = 32'd4120
; 
32'd146672: dataIn1 = 32'd4121
; 
32'd146673: dataIn1 = 32'd1987
; 
32'd146674: dataIn1 = 32'd2358
; 
32'd146675: dataIn1 = 32'd3116
; 
32'd146676: dataIn1 = 32'd4111
; 
32'd146677: dataIn1 = 32'd4119
; 
32'd146678: dataIn1 = 32'd4120
; 
32'd146679: dataIn1 = 32'd4121
; 
32'd146680: dataIn1 = 32'd1987
; 
32'd146681: dataIn1 = 32'd2354
; 
32'd146682: dataIn1 = 32'd3117
; 
32'd146683: dataIn1 = 32'd4104
; 
32'd146684: dataIn1 = 32'd4119
; 
32'd146685: dataIn1 = 32'd4120
; 
32'd146686: dataIn1 = 32'd4121
; 
32'd146687: dataIn1 = 32'd2359
; 
32'd146688: dataIn1 = 32'd2361
; 
32'd146689: dataIn1 = 32'd4122
; 
32'd146690: dataIn1 = 32'd4123
; 
32'd146691: dataIn1 = 32'd4124
; 
32'd146692: dataIn1 = 32'd4125
; 
32'd146693: dataIn1 = 32'd4126
; 
32'd146694: dataIn1 = 32'd2359
; 
32'd146695: dataIn1 = 32'd2360
; 
32'd146696: dataIn1 = 32'd4118
; 
32'd146697: dataIn1 = 32'd4122
; 
32'd146698: dataIn1 = 32'd4123
; 
32'd146699: dataIn1 = 32'd4124
; 
32'd146700: dataIn1 = 32'd4127
; 
32'd146701: dataIn1 = 32'd2360
; 
32'd146702: dataIn1 = 32'd2361
; 
32'd146703: dataIn1 = 32'd4122
; 
32'd146704: dataIn1 = 32'd4123
; 
32'd146705: dataIn1 = 32'd4124
; 
32'd146706: dataIn1 = 32'd4128
; 
32'd146707: dataIn1 = 32'd4129
; 
32'd146708: dataIn1 = 32'd163
; 
32'd146709: dataIn1 = 32'd2359
; 
32'd146710: dataIn1 = 32'd3121
; 
32'd146711: dataIn1 = 32'd4115
; 
32'd146712: dataIn1 = 32'd4122
; 
32'd146713: dataIn1 = 32'd4125
; 
32'd146714: dataIn1 = 32'd4126
; 
32'd146715: dataIn1 = 32'd163
; 
32'd146716: dataIn1 = 32'd2361
; 
32'd146717: dataIn1 = 32'd3128
; 
32'd146718: dataIn1 = 32'd4122
; 
32'd146719: dataIn1 = 32'd4125
; 
32'd146720: dataIn1 = 32'd4126
; 
32'd146721: dataIn1 = 32'd4139
; 
32'd146722: dataIn1 = 32'd463
; 
32'd146723: dataIn1 = 32'd2360
; 
32'd146724: dataIn1 = 32'd4118
; 
32'd146725: dataIn1 = 32'd4123
; 
32'd146726: dataIn1 = 32'd4127
; 
32'd146727: dataIn1 = 32'd5347
; 
32'd146728: dataIn1 = 32'd464
; 
32'd146729: dataIn1 = 32'd2361
; 
32'd146730: dataIn1 = 32'd4124
; 
32'd146731: dataIn1 = 32'd4128
; 
32'd146732: dataIn1 = 32'd4129
; 
32'd146733: dataIn1 = 32'd4138
; 
32'd146734: dataIn1 = 32'd4141
; 
32'd146735: dataIn1 = 32'd464
; 
32'd146736: dataIn1 = 32'd2360
; 
32'd146737: dataIn1 = 32'd4124
; 
32'd146738: dataIn1 = 32'd4128
; 
32'd146739: dataIn1 = 32'd4129
; 
32'd146740: dataIn1 = 32'd5346
; 
32'd146741: dataIn1 = 32'd2363
; 
32'd146742: dataIn1 = 32'd2364
; 
32'd146743: dataIn1 = 32'd4130
; 
32'd146744: dataIn1 = 32'd4131
; 
32'd146745: dataIn1 = 32'd4132
; 
32'd146746: dataIn1 = 32'd4133
; 
32'd146747: dataIn1 = 32'd4134
; 
32'd146748: dataIn1 = 32'd2362
; 
32'd146749: dataIn1 = 32'd2364
; 
32'd146750: dataIn1 = 32'd4130
; 
32'd146751: dataIn1 = 32'd4131
; 
32'd146752: dataIn1 = 32'd4132
; 
32'd146753: dataIn1 = 32'd4135
; 
32'd146754: dataIn1 = 32'd4136
; 
32'd146755: dataIn1 = 32'd2362
; 
32'd146756: dataIn1 = 32'd2363
; 
32'd146757: dataIn1 = 32'd4130
; 
32'd146758: dataIn1 = 32'd4131
; 
32'd146759: dataIn1 = 32'd4132
; 
32'd146760: dataIn1 = 32'd4137
; 
32'd146761: dataIn1 = 32'd4138
; 
32'd146762: dataIn1 = 32'd465
; 
32'd146763: dataIn1 = 32'd2364
; 
32'd146764: dataIn1 = 32'd4130
; 
32'd146765: dataIn1 = 32'd4133
; 
32'd146766: dataIn1 = 32'd4134
; 
32'd146767: dataIn1 = 32'd4142
; 
32'd146768: dataIn1 = 32'd4145
; 
32'd146769: dataIn1 = 32'd465
; 
32'd146770: dataIn1 = 32'd2363
; 
32'd146771: dataIn1 = 32'd4130
; 
32'd146772: dataIn1 = 32'd4133
; 
32'd146773: dataIn1 = 32'd4134
; 
32'd146774: dataIn1 = 32'd5349
; 
32'd146775: dataIn1 = 32'd309
; 
32'd146776: dataIn1 = 32'd2364
; 
32'd146777: dataIn1 = 32'd3137
; 
32'd146778: dataIn1 = 32'd4131
; 
32'd146779: dataIn1 = 32'd4135
; 
32'd146780: dataIn1 = 32'd4136
; 
32'd146781: dataIn1 = 32'd4143
; 
32'd146782: dataIn1 = 32'd309
; 
32'd146783: dataIn1 = 32'd2362
; 
32'd146784: dataIn1 = 32'd3129
; 
32'd146785: dataIn1 = 32'd4131
; 
32'd146786: dataIn1 = 32'd4135
; 
32'd146787: dataIn1 = 32'd4136
; 
32'd146788: dataIn1 = 32'd4140
; 
32'd146789: dataIn1 = 32'd464
; 
32'd146790: dataIn1 = 32'd2363
; 
32'd146791: dataIn1 = 32'd4132
; 
32'd146792: dataIn1 = 32'd4137
; 
32'd146793: dataIn1 = 32'd4138
; 
32'd146794: dataIn1 = 32'd5348
; 
32'd146795: dataIn1 = 32'd464
; 
32'd146796: dataIn1 = 32'd2362
; 
32'd146797: dataIn1 = 32'd4128
; 
32'd146798: dataIn1 = 32'd4132
; 
32'd146799: dataIn1 = 32'd4137
; 
32'd146800: dataIn1 = 32'd4138
; 
32'd146801: dataIn1 = 32'd4141
; 
32'd146802: dataIn1 = 32'd1989
; 
32'd146803: dataIn1 = 32'd2361
; 
32'd146804: dataIn1 = 32'd3128
; 
32'd146805: dataIn1 = 32'd4126
; 
32'd146806: dataIn1 = 32'd4139
; 
32'd146807: dataIn1 = 32'd4140
; 
32'd146808: dataIn1 = 32'd4141
; 
32'd146809: dataIn1 = 32'd1989
; 
32'd146810: dataIn1 = 32'd2362
; 
32'd146811: dataIn1 = 32'd3129
; 
32'd146812: dataIn1 = 32'd4136
; 
32'd146813: dataIn1 = 32'd4139
; 
32'd146814: dataIn1 = 32'd4140
; 
32'd146815: dataIn1 = 32'd4141
; 
32'd146816: dataIn1 = 32'd2361
; 
32'd146817: dataIn1 = 32'd2362
; 
32'd146818: dataIn1 = 32'd4128
; 
32'd146819: dataIn1 = 32'd4138
; 
32'd146820: dataIn1 = 32'd4139
; 
32'd146821: dataIn1 = 32'd4140
; 
32'd146822: dataIn1 = 32'd4141
; 
32'd146823: dataIn1 = 32'd2364
; 
32'd146824: dataIn1 = 32'd2365
; 
32'd146825: dataIn1 = 32'd4133
; 
32'd146826: dataIn1 = 32'd4142
; 
32'd146827: dataIn1 = 32'd4143
; 
32'd146828: dataIn1 = 32'd4144
; 
32'd146829: dataIn1 = 32'd4145
; 
32'd146830: dataIn1 = 32'd1990
; 
32'd146831: dataIn1 = 32'd2364
; 
32'd146832: dataIn1 = 32'd3137
; 
32'd146833: dataIn1 = 32'd4135
; 
32'd146834: dataIn1 = 32'd4142
; 
32'd146835: dataIn1 = 32'd4143
; 
32'd146836: dataIn1 = 32'd4144
; 
32'd146837: dataIn1 = 32'd1990
; 
32'd146838: dataIn1 = 32'd2365
; 
32'd146839: dataIn1 = 32'd3138
; 
32'd146840: dataIn1 = 32'd4142
; 
32'd146841: dataIn1 = 32'd4143
; 
32'd146842: dataIn1 = 32'd4144
; 
32'd146843: dataIn1 = 32'd4152
; 
32'd146844: dataIn1 = 32'd465
; 
32'd146845: dataIn1 = 32'd2365
; 
32'd146846: dataIn1 = 32'd4133
; 
32'd146847: dataIn1 = 32'd4142
; 
32'd146848: dataIn1 = 32'd4145
; 
32'd146849: dataIn1 = 32'd4146
; 
32'd146850: dataIn1 = 32'd4149
; 
32'd146851: dataIn1 = 32'd2365
; 
32'd146852: dataIn1 = 32'd2367
; 
32'd146853: dataIn1 = 32'd4145
; 
32'd146854: dataIn1 = 32'd4146
; 
32'd146855: dataIn1 = 32'd4147
; 
32'd146856: dataIn1 = 32'd4148
; 
32'd146857: dataIn1 = 32'd4149
; 
32'd146858: dataIn1 = 32'd2366
; 
32'd146859: dataIn1 = 32'd2367
; 
32'd146860: dataIn1 = 32'd4146
; 
32'd146861: dataIn1 = 32'd4147
; 
32'd146862: dataIn1 = 32'd4148
; 
32'd146863: dataIn1 = 32'd4150
; 
32'd146864: dataIn1 = 32'd4151
; 
32'd146865: dataIn1 = 32'd2365
; 
32'd146866: dataIn1 = 32'd2366
; 
32'd146867: dataIn1 = 32'd4146
; 
32'd146868: dataIn1 = 32'd4147
; 
32'd146869: dataIn1 = 32'd4148
; 
32'd146870: dataIn1 = 32'd4152
; 
32'd146871: dataIn1 = 32'd4153
; 
32'd146872: dataIn1 = 32'd465
; 
32'd146873: dataIn1 = 32'd2367
; 
32'd146874: dataIn1 = 32'd4145
; 
32'd146875: dataIn1 = 32'd4146
; 
32'd146876: dataIn1 = 32'd4149
; 
32'd146877: dataIn1 = 32'd5351
; 
32'd146878: dataIn1 = 32'd466
; 
32'd146879: dataIn1 = 32'd2367
; 
32'd146880: dataIn1 = 32'd4147
; 
32'd146881: dataIn1 = 32'd4150
; 
32'd146882: dataIn1 = 32'd4151
; 
32'd146883: dataIn1 = 32'd5350
; 
32'd146884: dataIn1 = 32'd466
; 
32'd146885: dataIn1 = 32'd2366
; 
32'd146886: dataIn1 = 32'd4147
; 
32'd146887: dataIn1 = 32'd4150
; 
32'd146888: dataIn1 = 32'd4151
; 
32'd146889: dataIn1 = 32'd4160
; 
32'd146890: dataIn1 = 32'd4164
; 
32'd146891: dataIn1 = 32'd165
; 
32'd146892: dataIn1 = 32'd2365
; 
32'd146893: dataIn1 = 32'd3138
; 
32'd146894: dataIn1 = 32'd4144
; 
32'd146895: dataIn1 = 32'd4148
; 
32'd146896: dataIn1 = 32'd4152
; 
32'd146897: dataIn1 = 32'd4153
; 
32'd146898: dataIn1 = 32'd165
; 
32'd146899: dataIn1 = 32'd2366
; 
32'd146900: dataIn1 = 32'd3163
; 
32'd146901: dataIn1 = 32'd4148
; 
32'd146902: dataIn1 = 32'd4152
; 
32'd146903: dataIn1 = 32'd4153
; 
32'd146904: dataIn1 = 32'd4163
; 
32'd146905: dataIn1 = 32'd2369
; 
32'd146906: dataIn1 = 32'd2370
; 
32'd146907: dataIn1 = 32'd4154
; 
32'd146908: dataIn1 = 32'd4155
; 
32'd146909: dataIn1 = 32'd4156
; 
32'd146910: dataIn1 = 32'd4157
; 
32'd146911: dataIn1 = 32'd4158
; 
32'd146912: dataIn1 = 32'd2368
; 
32'd146913: dataIn1 = 32'd2370
; 
32'd146914: dataIn1 = 32'd4154
; 
32'd146915: dataIn1 = 32'd4155
; 
32'd146916: dataIn1 = 32'd4156
; 
32'd146917: dataIn1 = 32'd4159
; 
32'd146918: dataIn1 = 32'd4160
; 
32'd146919: dataIn1 = 32'd2368
; 
32'd146920: dataIn1 = 32'd2369
; 
32'd146921: dataIn1 = 32'd4154
; 
32'd146922: dataIn1 = 32'd4155
; 
32'd146923: dataIn1 = 32'd4156
; 
32'd146924: dataIn1 = 32'd4161
; 
32'd146925: dataIn1 = 32'd4162
; 
32'd146926: dataIn1 = 32'd467
; 
32'd146927: dataIn1 = 32'd2370
; 
32'd146928: dataIn1 = 32'd4154
; 
32'd146929: dataIn1 = 32'd4157
; 
32'd146930: dataIn1 = 32'd4158
; 
32'd146931: dataIn1 = 32'd5353
; 
32'd146932: dataIn1 = 32'd467
; 
32'd146933: dataIn1 = 32'd2369
; 
32'd146934: dataIn1 = 32'd4154
; 
32'd146935: dataIn1 = 32'd4157
; 
32'd146936: dataIn1 = 32'd4158
; 
32'd146937: dataIn1 = 32'd4166
; 
32'd146938: dataIn1 = 32'd4169
; 
32'd146939: dataIn1 = 32'd466
; 
32'd146940: dataIn1 = 32'd2370
; 
32'd146941: dataIn1 = 32'd4155
; 
32'd146942: dataIn1 = 32'd4159
; 
32'd146943: dataIn1 = 32'd4160
; 
32'd146944: dataIn1 = 32'd5352
; 
32'd146945: dataIn1 = 32'd466
; 
32'd146946: dataIn1 = 32'd2368
; 
32'd146947: dataIn1 = 32'd4151
; 
32'd146948: dataIn1 = 32'd4155
; 
32'd146949: dataIn1 = 32'd4159
; 
32'd146950: dataIn1 = 32'd4160
; 
32'd146951: dataIn1 = 32'd4164
; 
32'd146952: dataIn1 = 32'd317
; 
32'd146953: dataIn1 = 32'd2369
; 
32'd146954: dataIn1 = 32'd3159
; 
32'd146955: dataIn1 = 32'd4156
; 
32'd146956: dataIn1 = 32'd4161
; 
32'd146957: dataIn1 = 32'd4162
; 
32'd146958: dataIn1 = 32'd4168
; 
32'd146959: dataIn1 = 32'd317
; 
32'd146960: dataIn1 = 32'd2368
; 
32'd146961: dataIn1 = 32'd3166
; 
32'd146962: dataIn1 = 32'd4156
; 
32'd146963: dataIn1 = 32'd4161
; 
32'd146964: dataIn1 = 32'd4162
; 
32'd146965: dataIn1 = 32'd4165
; 
32'd146966: dataIn1 = 32'd1994
; 
32'd146967: dataIn1 = 32'd2366
; 
32'd146968: dataIn1 = 32'd3163
; 
32'd146969: dataIn1 = 32'd4153
; 
32'd146970: dataIn1 = 32'd4163
; 
32'd146971: dataIn1 = 32'd4164
; 
32'd146972: dataIn1 = 32'd4165
; 
32'd146973: dataIn1 = 32'd2366
; 
32'd146974: dataIn1 = 32'd2368
; 
32'd146975: dataIn1 = 32'd4151
; 
32'd146976: dataIn1 = 32'd4160
; 
32'd146977: dataIn1 = 32'd4163
; 
32'd146978: dataIn1 = 32'd4164
; 
32'd146979: dataIn1 = 32'd4165
; 
32'd146980: dataIn1 = 32'd1994
; 
32'd146981: dataIn1 = 32'd2368
; 
32'd146982: dataIn1 = 32'd3166
; 
32'd146983: dataIn1 = 32'd4162
; 
32'd146984: dataIn1 = 32'd4163
; 
32'd146985: dataIn1 = 32'd4164
; 
32'd146986: dataIn1 = 32'd4165
; 
32'd146987: dataIn1 = 32'd2369
; 
32'd146988: dataIn1 = 32'd2371
; 
32'd146989: dataIn1 = 32'd4158
; 
32'd146990: dataIn1 = 32'd4166
; 
32'd146991: dataIn1 = 32'd4167
; 
32'd146992: dataIn1 = 32'd4168
; 
32'd146993: dataIn1 = 32'd4169
; 
32'd146994: dataIn1 = 32'd1993
; 
32'd146995: dataIn1 = 32'd2371
; 
32'd146996: dataIn1 = 32'd3158
; 
32'd146997: dataIn1 = 32'd4166
; 
32'd146998: dataIn1 = 32'd4167
; 
32'd146999: dataIn1 = 32'd4168
; 
32'd147000: dataIn1 = 32'd4174
; 
32'd147001: dataIn1 = 32'd1993
; 
32'd147002: dataIn1 = 32'd2369
; 
32'd147003: dataIn1 = 32'd3159
; 
32'd147004: dataIn1 = 32'd4161
; 
32'd147005: dataIn1 = 32'd4166
; 
32'd147006: dataIn1 = 32'd4167
; 
32'd147007: dataIn1 = 32'd4168
; 
32'd147008: dataIn1 = 32'd467
; 
32'd147009: dataIn1 = 32'd2371
; 
32'd147010: dataIn1 = 32'd4158
; 
32'd147011: dataIn1 = 32'd4166
; 
32'd147012: dataIn1 = 32'd4169
; 
32'd147013: dataIn1 = 32'd4170
; 
32'd147014: dataIn1 = 32'd4173
; 
32'd147015: dataIn1 = 32'd2371
; 
32'd147016: dataIn1 = 32'd2373
; 
32'd147017: dataIn1 = 32'd4169
; 
32'd147018: dataIn1 = 32'd4170
; 
32'd147019: dataIn1 = 32'd4171
; 
32'd147020: dataIn1 = 32'd4172
; 
32'd147021: dataIn1 = 32'd4173
; 
32'd147022: dataIn1 = 32'd2371
; 
32'd147023: dataIn1 = 32'd2372
; 
32'd147024: dataIn1 = 32'd4170
; 
32'd147025: dataIn1 = 32'd4171
; 
32'd147026: dataIn1 = 32'd4172
; 
32'd147027: dataIn1 = 32'd4174
; 
32'd147028: dataIn1 = 32'd4175
; 
32'd147029: dataIn1 = 32'd2372
; 
32'd147030: dataIn1 = 32'd2373
; 
32'd147031: dataIn1 = 32'd4170
; 
32'd147032: dataIn1 = 32'd4171
; 
32'd147033: dataIn1 = 32'd4172
; 
32'd147034: dataIn1 = 32'd4176
; 
32'd147035: dataIn1 = 32'd4177
; 
32'd147036: dataIn1 = 32'd467
; 
32'd147037: dataIn1 = 32'd2373
; 
32'd147038: dataIn1 = 32'd4169
; 
32'd147039: dataIn1 = 32'd4170
; 
32'd147040: dataIn1 = 32'd4173
; 
32'd147041: dataIn1 = 32'd5355
; 
32'd147042: dataIn1 = 32'd167
; 
32'd147043: dataIn1 = 32'd2371
; 
32'd147044: dataIn1 = 32'd3158
; 
32'd147045: dataIn1 = 32'd4167
; 
32'd147046: dataIn1 = 32'd4171
; 
32'd147047: dataIn1 = 32'd4174
; 
32'd147048: dataIn1 = 32'd4175
; 
32'd147049: dataIn1 = 32'd167
; 
32'd147050: dataIn1 = 32'd2372
; 
32'd147051: dataIn1 = 32'd3150
; 
32'd147052: dataIn1 = 32'd4171
; 
32'd147053: dataIn1 = 32'd4174
; 
32'd147054: dataIn1 = 32'd4175
; 
32'd147055: dataIn1 = 32'd4188
; 
32'd147056: dataIn1 = 32'd468
; 
32'd147057: dataIn1 = 32'd2373
; 
32'd147058: dataIn1 = 32'd4172
; 
32'd147059: dataIn1 = 32'd4176
; 
32'd147060: dataIn1 = 32'd4177
; 
32'd147061: dataIn1 = 32'd5354
; 
32'd147062: dataIn1 = 32'd468
; 
32'd147063: dataIn1 = 32'd2372
; 
32'd147064: dataIn1 = 32'd4172
; 
32'd147065: dataIn1 = 32'd4176
; 
32'd147066: dataIn1 = 32'd4177
; 
32'd147067: dataIn1 = 32'd4185
; 
32'd147068: dataIn1 = 32'd4189
; 
32'd147069: dataIn1 = 32'd2375
; 
32'd147070: dataIn1 = 32'd2376
; 
32'd147071: dataIn1 = 32'd4178
; 
32'd147072: dataIn1 = 32'd4179
; 
32'd147073: dataIn1 = 32'd4180
; 
32'd147074: dataIn1 = 32'd4181
; 
32'd147075: dataIn1 = 32'd4182
; 
32'd147076: dataIn1 = 32'd2374
; 
32'd147077: dataIn1 = 32'd2376
; 
32'd147078: dataIn1 = 32'd4178
; 
32'd147079: dataIn1 = 32'd4179
; 
32'd147080: dataIn1 = 32'd4180
; 
32'd147081: dataIn1 = 32'd4183
; 
32'd147082: dataIn1 = 32'd4184
; 
32'd147083: dataIn1 = 32'd2374
; 
32'd147084: dataIn1 = 32'd2375
; 
32'd147085: dataIn1 = 32'd4178
; 
32'd147086: dataIn1 = 32'd4179
; 
32'd147087: dataIn1 = 32'd4180
; 
32'd147088: dataIn1 = 32'd4185
; 
32'd147089: dataIn1 = 32'd4186
; 
32'd147090: dataIn1 = 32'd311
; 
32'd147091: dataIn1 = 32'd2376
; 
32'd147092: dataIn1 = 32'd3142
; 
32'd147093: dataIn1 = 32'd4178
; 
32'd147094: dataIn1 = 32'd4181
; 
32'd147095: dataIn1 = 32'd4182
; 
32'd147096: dataIn1 = 32'd4190
; 
32'd147097: dataIn1 = 32'd311
; 
32'd147098: dataIn1 = 32'd2375
; 
32'd147099: dataIn1 = 32'd3149
; 
32'd147100: dataIn1 = 32'd4178
; 
32'd147101: dataIn1 = 32'd4181
; 
32'd147102: dataIn1 = 32'd4182
; 
32'd147103: dataIn1 = 32'd4187
; 
32'd147104: dataIn1 = 32'd469
; 
32'd147105: dataIn1 = 32'd2376
; 
32'd147106: dataIn1 = 32'd4179
; 
32'd147107: dataIn1 = 32'd4183
; 
32'd147108: dataIn1 = 32'd4184
; 
32'd147109: dataIn1 = 32'd4191
; 
32'd147110: dataIn1 = 32'd4193
; 
32'd147111: dataIn1 = 32'd469
; 
32'd147112: dataIn1 = 32'd2374
; 
32'd147113: dataIn1 = 32'd4179
; 
32'd147114: dataIn1 = 32'd4183
; 
32'd147115: dataIn1 = 32'd4184
; 
32'd147116: dataIn1 = 32'd5357
; 
32'd147117: dataIn1 = 32'd468
; 
32'd147118: dataIn1 = 32'd2375
; 
32'd147119: dataIn1 = 32'd4177
; 
32'd147120: dataIn1 = 32'd4180
; 
32'd147121: dataIn1 = 32'd4185
; 
32'd147122: dataIn1 = 32'd4186
; 
32'd147123: dataIn1 = 32'd4189
; 
32'd147124: dataIn1 = 32'd468
; 
32'd147125: dataIn1 = 32'd2374
; 
32'd147126: dataIn1 = 32'd4180
; 
32'd147127: dataIn1 = 32'd4185
; 
32'd147128: dataIn1 = 32'd4186
; 
32'd147129: dataIn1 = 32'd5356
; 
32'd147130: dataIn1 = 32'd1992
; 
32'd147131: dataIn1 = 32'd2375
; 
32'd147132: dataIn1 = 32'd3149
; 
32'd147133: dataIn1 = 32'd4182
; 
32'd147134: dataIn1 = 32'd4187
; 
32'd147135: dataIn1 = 32'd4188
; 
32'd147136: dataIn1 = 32'd4189
; 
32'd147137: dataIn1 = 32'd1992
; 
32'd147138: dataIn1 = 32'd2372
; 
32'd147139: dataIn1 = 32'd3150
; 
32'd147140: dataIn1 = 32'd4175
; 
32'd147141: dataIn1 = 32'd4187
; 
32'd147142: dataIn1 = 32'd4188
; 
32'd147143: dataIn1 = 32'd4189
; 
32'd147144: dataIn1 = 32'd2372
; 
32'd147145: dataIn1 = 32'd2375
; 
32'd147146: dataIn1 = 32'd4177
; 
32'd147147: dataIn1 = 32'd4185
; 
32'd147148: dataIn1 = 32'd4187
; 
32'd147149: dataIn1 = 32'd4188
; 
32'd147150: dataIn1 = 32'd4189
; 
32'd147151: dataIn1 = 32'd1991
; 
32'd147152: dataIn1 = 32'd2376
; 
32'd147153: dataIn1 = 32'd3142
; 
32'd147154: dataIn1 = 32'd4181
; 
32'd147155: dataIn1 = 32'd4190
; 
32'd147156: dataIn1 = 32'd4191
; 
32'd147157: dataIn1 = 32'd4192
; 
32'd147158: dataIn1 = 32'd2376
; 
32'd147159: dataIn1 = 32'd2377
; 
32'd147160: dataIn1 = 32'd4183
; 
32'd147161: dataIn1 = 32'd4190
; 
32'd147162: dataIn1 = 32'd4191
; 
32'd147163: dataIn1 = 32'd4192
; 
32'd147164: dataIn1 = 32'd4193
; 
32'd147165: dataIn1 = 32'd1991
; 
32'd147166: dataIn1 = 32'd2377
; 
32'd147167: dataIn1 = 32'd3145
; 
32'd147168: dataIn1 = 32'd4190
; 
32'd147169: dataIn1 = 32'd4191
; 
32'd147170: dataIn1 = 32'd4192
; 
32'd147171: dataIn1 = 32'd4201
; 
32'd147172: dataIn1 = 32'd469
; 
32'd147173: dataIn1 = 32'd2377
; 
32'd147174: dataIn1 = 32'd4183
; 
32'd147175: dataIn1 = 32'd4191
; 
32'd147176: dataIn1 = 32'd4193
; 
32'd147177: dataIn1 = 32'd4195
; 
32'd147178: dataIn1 = 32'd4199
; 
32'd147179: dataIn1 = 32'd2378
; 
32'd147180: dataIn1 = 32'd2379
; 
32'd147181: dataIn1 = 32'd4194
; 
32'd147182: dataIn1 = 32'd4195
; 
32'd147183: dataIn1 = 32'd4196
; 
32'd147184: dataIn1 = 32'd4197
; 
32'd147185: dataIn1 = 32'd4198
; 
32'd147186: dataIn1 = 32'd2377
; 
32'd147187: dataIn1 = 32'd2379
; 
32'd147188: dataIn1 = 32'd4193
; 
32'd147189: dataIn1 = 32'd4194
; 
32'd147190: dataIn1 = 32'd4195
; 
32'd147191: dataIn1 = 32'd4196
; 
32'd147192: dataIn1 = 32'd4199
; 
32'd147193: dataIn1 = 32'd2377
; 
32'd147194: dataIn1 = 32'd2378
; 
32'd147195: dataIn1 = 32'd4194
; 
32'd147196: dataIn1 = 32'd4195
; 
32'd147197: dataIn1 = 32'd4196
; 
32'd147198: dataIn1 = 32'd4200
; 
32'd147199: dataIn1 = 32'd4201
; 
32'd147200: dataIn1 = 32'd470
; 
32'd147201: dataIn1 = 32'd2379
; 
32'd147202: dataIn1 = 32'd4194
; 
32'd147203: dataIn1 = 32'd4197
; 
32'd147204: dataIn1 = 32'd4198
; 
32'd147205: dataIn1 = 32'd5359
; 
32'd147206: dataIn1 = 32'd470
; 
32'd147207: dataIn1 = 32'd2378
; 
32'd147208: dataIn1 = 32'd4194
; 
32'd147209: dataIn1 = 32'd4197
; 
32'd147210: dataIn1 = 32'd4198
; 
32'd147211: dataIn1 = 32'd4205
; 
32'd147212: dataIn1 = 32'd4215
; 
32'd147213: dataIn1 = 32'd469
; 
32'd147214: dataIn1 = 32'd2379
; 
32'd147215: dataIn1 = 32'd4193
; 
32'd147216: dataIn1 = 32'd4195
; 
32'd147217: dataIn1 = 32'd4199
; 
32'd147218: dataIn1 = 32'd5358
; 
32'd147219: dataIn1 = 32'd168
; 
32'd147220: dataIn1 = 32'd2378
; 
32'd147221: dataIn1 = 32'd3173
; 
32'd147222: dataIn1 = 32'd4196
; 
32'd147223: dataIn1 = 32'd4200
; 
32'd147224: dataIn1 = 32'd4201
; 
32'd147225: dataIn1 = 32'd4217
; 
32'd147226: dataIn1 = 32'd168
; 
32'd147227: dataIn1 = 32'd2377
; 
32'd147228: dataIn1 = 32'd3145
; 
32'd147229: dataIn1 = 32'd4192
; 
32'd147230: dataIn1 = 32'd4196
; 
32'd147231: dataIn1 = 32'd4200
; 
32'd147232: dataIn1 = 32'd4201
; 
32'd147233: dataIn1 = 32'd2381
; 
32'd147234: dataIn1 = 32'd2382
; 
32'd147235: dataIn1 = 32'd4202
; 
32'd147236: dataIn1 = 32'd4203
; 
32'd147237: dataIn1 = 32'd4204
; 
32'd147238: dataIn1 = 32'd4205
; 
32'd147239: dataIn1 = 32'd4206
; 
32'd147240: dataIn1 = 32'd2380
; 
32'd147241: dataIn1 = 32'd2382
; 
32'd147242: dataIn1 = 32'd4202
; 
32'd147243: dataIn1 = 32'd4203
; 
32'd147244: dataIn1 = 32'd4204
; 
32'd147245: dataIn1 = 32'd4207
; 
32'd147246: dataIn1 = 32'd4208
; 
32'd147247: dataIn1 = 32'd2380
; 
32'd147248: dataIn1 = 32'd2381
; 
32'd147249: dataIn1 = 32'd4202
; 
32'd147250: dataIn1 = 32'd4203
; 
32'd147251: dataIn1 = 32'd4204
; 
32'd147252: dataIn1 = 32'd4209
; 
32'd147253: dataIn1 = 32'd4210
; 
32'd147254: dataIn1 = 32'd470
; 
32'd147255: dataIn1 = 32'd2382
; 
32'd147256: dataIn1 = 32'd4198
; 
32'd147257: dataIn1 = 32'd4202
; 
32'd147258: dataIn1 = 32'd4205
; 
32'd147259: dataIn1 = 32'd4206
; 
32'd147260: dataIn1 = 32'd4215
; 
32'd147261: dataIn1 = 32'd470
; 
32'd147262: dataIn1 = 32'd2381
; 
32'd147263: dataIn1 = 32'd4202
; 
32'd147264: dataIn1 = 32'd4205
; 
32'd147265: dataIn1 = 32'd4206
; 
32'd147266: dataIn1 = 32'd5361
; 
32'd147267: dataIn1 = 32'd318
; 
32'd147268: dataIn1 = 32'd2382
; 
32'd147269: dataIn1 = 32'd3172
; 
32'd147270: dataIn1 = 32'd4203
; 
32'd147271: dataIn1 = 32'd4207
; 
32'd147272: dataIn1 = 32'd4208
; 
32'd147273: dataIn1 = 32'd4216
; 
32'd147274: dataIn1 = 32'd318
; 
32'd147275: dataIn1 = 32'd2380
; 
32'd147276: dataIn1 = 32'd3178
; 
32'd147277: dataIn1 = 32'd4203
; 
32'd147278: dataIn1 = 32'd4207
; 
32'd147279: dataIn1 = 32'd4208
; 
32'd147280: dataIn1 = 32'd4212
; 
32'd147281: dataIn1 = 32'd471
; 
32'd147282: dataIn1 = 32'd2381
; 
32'd147283: dataIn1 = 32'd4204
; 
32'd147284: dataIn1 = 32'd4209
; 
32'd147285: dataIn1 = 32'd4210
; 
32'd147286: dataIn1 = 32'd5360
; 
32'd147287: dataIn1 = 32'd471
; 
32'd147288: dataIn1 = 32'd2380
; 
32'd147289: dataIn1 = 32'd4204
; 
32'd147290: dataIn1 = 32'd4209
; 
32'd147291: dataIn1 = 32'd4210
; 
32'd147292: dataIn1 = 32'd4213
; 
32'd147293: dataIn1 = 32'd4214
; 
32'd147294: dataIn1 = 32'd1996
; 
32'd147295: dataIn1 = 32'd2383
; 
32'd147296: dataIn1 = 32'd3177
; 
32'd147297: dataIn1 = 32'd4211
; 
32'd147298: dataIn1 = 32'd4212
; 
32'd147299: dataIn1 = 32'd4213
; 
32'd147300: dataIn1 = 32'd4221
; 
32'd147301: dataIn1 = 32'd1996
; 
32'd147302: dataIn1 = 32'd2380
; 
32'd147303: dataIn1 = 32'd3178
; 
32'd147304: dataIn1 = 32'd4208
; 
32'd147305: dataIn1 = 32'd4211
; 
32'd147306: dataIn1 = 32'd4212
; 
32'd147307: dataIn1 = 32'd4213
; 
32'd147308: dataIn1 = 32'd2380
; 
32'd147309: dataIn1 = 32'd2383
; 
32'd147310: dataIn1 = 32'd4210
; 
32'd147311: dataIn1 = 32'd4211
; 
32'd147312: dataIn1 = 32'd4212
; 
32'd147313: dataIn1 = 32'd4213
; 
32'd147314: dataIn1 = 32'd4214
; 
32'd147315: dataIn1 = 32'd471
; 
32'd147316: dataIn1 = 32'd2383
; 
32'd147317: dataIn1 = 32'd4210
; 
32'd147318: dataIn1 = 32'd4213
; 
32'd147319: dataIn1 = 32'd4214
; 
32'd147320: dataIn1 = 32'd4219
; 
32'd147321: dataIn1 = 32'd4223
; 
32'd147322: dataIn1 = 32'd2378
; 
32'd147323: dataIn1 = 32'd2382
; 
32'd147324: dataIn1 = 32'd4198
; 
32'd147325: dataIn1 = 32'd4205
; 
32'd147326: dataIn1 = 32'd4215
; 
32'd147327: dataIn1 = 32'd4216
; 
32'd147328: dataIn1 = 32'd4217
; 
32'd147329: dataIn1 = 32'd1995
; 
32'd147330: dataIn1 = 32'd2382
; 
32'd147331: dataIn1 = 32'd3172
; 
32'd147332: dataIn1 = 32'd4207
; 
32'd147333: dataIn1 = 32'd4215
; 
32'd147334: dataIn1 = 32'd4216
; 
32'd147335: dataIn1 = 32'd4217
; 
32'd147336: dataIn1 = 32'd1995
; 
32'd147337: dataIn1 = 32'd2378
; 
32'd147338: dataIn1 = 32'd3173
; 
32'd147339: dataIn1 = 32'd4200
; 
32'd147340: dataIn1 = 32'd4215
; 
32'd147341: dataIn1 = 32'd4216
; 
32'd147342: dataIn1 = 32'd4217
; 
32'd147343: dataIn1 = 32'd2383
; 
32'd147344: dataIn1 = 32'd2385
; 
32'd147345: dataIn1 = 32'd4218
; 
32'd147346: dataIn1 = 32'd4219
; 
32'd147347: dataIn1 = 32'd4220
; 
32'd147348: dataIn1 = 32'd4221
; 
32'd147349: dataIn1 = 32'd4222
; 
32'd147350: dataIn1 = 32'd2383
; 
32'd147351: dataIn1 = 32'd2384
; 
32'd147352: dataIn1 = 32'd4214
; 
32'd147353: dataIn1 = 32'd4218
; 
32'd147354: dataIn1 = 32'd4219
; 
32'd147355: dataIn1 = 32'd4220
; 
32'd147356: dataIn1 = 32'd4223
; 
32'd147357: dataIn1 = 32'd2384
; 
32'd147358: dataIn1 = 32'd2385
; 
32'd147359: dataIn1 = 32'd4218
; 
32'd147360: dataIn1 = 32'd4219
; 
32'd147361: dataIn1 = 32'd4220
; 
32'd147362: dataIn1 = 32'd4224
; 
32'd147363: dataIn1 = 32'd4225
; 
32'd147364: dataIn1 = 32'd169
; 
32'd147365: dataIn1 = 32'd2383
; 
32'd147366: dataIn1 = 32'd3177
; 
32'd147367: dataIn1 = 32'd4211
; 
32'd147368: dataIn1 = 32'd4218
; 
32'd147369: dataIn1 = 32'd4221
; 
32'd147370: dataIn1 = 32'd4222
; 
32'd147371: dataIn1 = 32'd169
; 
32'd147372: dataIn1 = 32'd2385
; 
32'd147373: dataIn1 = 32'd3184
; 
32'd147374: dataIn1 = 32'd4218
; 
32'd147375: dataIn1 = 32'd4221
; 
32'd147376: dataIn1 = 32'd4222
; 
32'd147377: dataIn1 = 32'd4235
; 
32'd147378: dataIn1 = 32'd471
; 
32'd147379: dataIn1 = 32'd2384
; 
32'd147380: dataIn1 = 32'd4214
; 
32'd147381: dataIn1 = 32'd4219
; 
32'd147382: dataIn1 = 32'd4223
; 
32'd147383: dataIn1 = 32'd5363
; 
32'd147384: dataIn1 = 32'd472
; 
32'd147385: dataIn1 = 32'd2385
; 
32'd147386: dataIn1 = 32'd4220
; 
32'd147387: dataIn1 = 32'd4224
; 
32'd147388: dataIn1 = 32'd4225
; 
32'd147389: dataIn1 = 32'd4234
; 
32'd147390: dataIn1 = 32'd4237
; 
32'd147391: dataIn1 = 32'd472
; 
32'd147392: dataIn1 = 32'd2384
; 
32'd147393: dataIn1 = 32'd4220
; 
32'd147394: dataIn1 = 32'd4224
; 
32'd147395: dataIn1 = 32'd4225
; 
32'd147396: dataIn1 = 32'd5362
; 
32'd147397: dataIn1 = 32'd2387
; 
32'd147398: dataIn1 = 32'd2388
; 
32'd147399: dataIn1 = 32'd4226
; 
32'd147400: dataIn1 = 32'd4227
; 
32'd147401: dataIn1 = 32'd4228
; 
32'd147402: dataIn1 = 32'd4229
; 
32'd147403: dataIn1 = 32'd4230
; 
32'd147404: dataIn1 = 32'd2386
; 
32'd147405: dataIn1 = 32'd2388
; 
32'd147406: dataIn1 = 32'd4226
; 
32'd147407: dataIn1 = 32'd4227
; 
32'd147408: dataIn1 = 32'd4228
; 
32'd147409: dataIn1 = 32'd4231
; 
32'd147410: dataIn1 = 32'd4232
; 
32'd147411: dataIn1 = 32'd2386
; 
32'd147412: dataIn1 = 32'd2387
; 
32'd147413: dataIn1 = 32'd4226
; 
32'd147414: dataIn1 = 32'd4227
; 
32'd147415: dataIn1 = 32'd4228
; 
32'd147416: dataIn1 = 32'd4233
; 
32'd147417: dataIn1 = 32'd4234
; 
32'd147418: dataIn1 = 32'd473
; 
32'd147419: dataIn1 = 32'd2388
; 
32'd147420: dataIn1 = 32'd4226
; 
32'd147421: dataIn1 = 32'd4229
; 
32'd147422: dataIn1 = 32'd4230
; 
32'd147423: dataIn1 = 32'd4238
; 
32'd147424: dataIn1 = 32'd4241
; 
32'd147425: dataIn1 = 32'd473
; 
32'd147426: dataIn1 = 32'd2387
; 
32'd147427: dataIn1 = 32'd4226
; 
32'd147428: dataIn1 = 32'd4229
; 
32'd147429: dataIn1 = 32'd4230
; 
32'd147430: dataIn1 = 32'd5365
; 
32'd147431: dataIn1 = 32'd325
; 
32'd147432: dataIn1 = 32'd2388
; 
32'd147433: dataIn1 = 32'd3193
; 
32'd147434: dataIn1 = 32'd4227
; 
32'd147435: dataIn1 = 32'd4231
; 
32'd147436: dataIn1 = 32'd4232
; 
32'd147437: dataIn1 = 32'd4239
; 
32'd147438: dataIn1 = 32'd325
; 
32'd147439: dataIn1 = 32'd2386
; 
32'd147440: dataIn1 = 32'd3185
; 
32'd147441: dataIn1 = 32'd4227
; 
32'd147442: dataIn1 = 32'd4231
; 
32'd147443: dataIn1 = 32'd4232
; 
32'd147444: dataIn1 = 32'd4236
; 
32'd147445: dataIn1 = 32'd472
; 
32'd147446: dataIn1 = 32'd2387
; 
32'd147447: dataIn1 = 32'd4228
; 
32'd147448: dataIn1 = 32'd4233
; 
32'd147449: dataIn1 = 32'd4234
; 
32'd147450: dataIn1 = 32'd5364
; 
32'd147451: dataIn1 = 32'd472
; 
32'd147452: dataIn1 = 32'd2386
; 
32'd147453: dataIn1 = 32'd4224
; 
32'd147454: dataIn1 = 32'd4228
; 
32'd147455: dataIn1 = 32'd4233
; 
32'd147456: dataIn1 = 32'd4234
; 
32'd147457: dataIn1 = 32'd4237
; 
32'd147458: dataIn1 = 32'd1997
; 
32'd147459: dataIn1 = 32'd2385
; 
32'd147460: dataIn1 = 32'd3184
; 
32'd147461: dataIn1 = 32'd4222
; 
32'd147462: dataIn1 = 32'd4235
; 
32'd147463: dataIn1 = 32'd4236
; 
32'd147464: dataIn1 = 32'd4237
; 
32'd147465: dataIn1 = 32'd1997
; 
32'd147466: dataIn1 = 32'd2386
; 
32'd147467: dataIn1 = 32'd3185
; 
32'd147468: dataIn1 = 32'd4232
; 
32'd147469: dataIn1 = 32'd4235
; 
32'd147470: dataIn1 = 32'd4236
; 
32'd147471: dataIn1 = 32'd4237
; 
32'd147472: dataIn1 = 32'd2385
; 
32'd147473: dataIn1 = 32'd2386
; 
32'd147474: dataIn1 = 32'd4224
; 
32'd147475: dataIn1 = 32'd4234
; 
32'd147476: dataIn1 = 32'd4235
; 
32'd147477: dataIn1 = 32'd4236
; 
32'd147478: dataIn1 = 32'd4237
; 
32'd147479: dataIn1 = 32'd2388
; 
32'd147480: dataIn1 = 32'd2389
; 
32'd147481: dataIn1 = 32'd4229
; 
32'd147482: dataIn1 = 32'd4238
; 
32'd147483: dataIn1 = 32'd4239
; 
32'd147484: dataIn1 = 32'd4240
; 
32'd147485: dataIn1 = 32'd4241
; 
32'd147486: dataIn1 = 32'd1998
; 
32'd147487: dataIn1 = 32'd2388
; 
32'd147488: dataIn1 = 32'd3193
; 
32'd147489: dataIn1 = 32'd4231
; 
32'd147490: dataIn1 = 32'd4238
; 
32'd147491: dataIn1 = 32'd4239
; 
32'd147492: dataIn1 = 32'd4240
; 
32'd147493: dataIn1 = 32'd1998
; 
32'd147494: dataIn1 = 32'd2389
; 
32'd147495: dataIn1 = 32'd3194
; 
32'd147496: dataIn1 = 32'd4238
; 
32'd147497: dataIn1 = 32'd4239
; 
32'd147498: dataIn1 = 32'd4240
; 
32'd147499: dataIn1 = 32'd4248
; 
32'd147500: dataIn1 = 32'd473
; 
32'd147501: dataIn1 = 32'd2389
; 
32'd147502: dataIn1 = 32'd4229
; 
32'd147503: dataIn1 = 32'd4238
; 
32'd147504: dataIn1 = 32'd4241
; 
32'd147505: dataIn1 = 32'd4242
; 
32'd147506: dataIn1 = 32'd4245
; 
32'd147507: dataIn1 = 32'd2389
; 
32'd147508: dataIn1 = 32'd2391
; 
32'd147509: dataIn1 = 32'd4241
; 
32'd147510: dataIn1 = 32'd4242
; 
32'd147511: dataIn1 = 32'd4243
; 
32'd147512: dataIn1 = 32'd4244
; 
32'd147513: dataIn1 = 32'd4245
; 
32'd147514: dataIn1 = 32'd2390
; 
32'd147515: dataIn1 = 32'd2391
; 
32'd147516: dataIn1 = 32'd4242
; 
32'd147517: dataIn1 = 32'd4243
; 
32'd147518: dataIn1 = 32'd4244
; 
32'd147519: dataIn1 = 32'd4246
; 
32'd147520: dataIn1 = 32'd4247
; 
32'd147521: dataIn1 = 32'd2389
; 
32'd147522: dataIn1 = 32'd2390
; 
32'd147523: dataIn1 = 32'd4242
; 
32'd147524: dataIn1 = 32'd4243
; 
32'd147525: dataIn1 = 32'd4244
; 
32'd147526: dataIn1 = 32'd4248
; 
32'd147527: dataIn1 = 32'd4249
; 
32'd147528: dataIn1 = 32'd473
; 
32'd147529: dataIn1 = 32'd2391
; 
32'd147530: dataIn1 = 32'd4241
; 
32'd147531: dataIn1 = 32'd4242
; 
32'd147532: dataIn1 = 32'd4245
; 
32'd147533: dataIn1 = 32'd5367
; 
32'd147534: dataIn1 = 32'd474
; 
32'd147535: dataIn1 = 32'd2391
; 
32'd147536: dataIn1 = 32'd4243
; 
32'd147537: dataIn1 = 32'd4246
; 
32'd147538: dataIn1 = 32'd4247
; 
32'd147539: dataIn1 = 32'd5366
; 
32'd147540: dataIn1 = 32'd474
; 
32'd147541: dataIn1 = 32'd2390
; 
32'd147542: dataIn1 = 32'd4243
; 
32'd147543: dataIn1 = 32'd4246
; 
32'd147544: dataIn1 = 32'd4247
; 
32'd147545: dataIn1 = 32'd4256
; 
32'd147546: dataIn1 = 32'd4260
; 
32'd147547: dataIn1 = 32'd171
; 
32'd147548: dataIn1 = 32'd2389
; 
32'd147549: dataIn1 = 32'd3194
; 
32'd147550: dataIn1 = 32'd4240
; 
32'd147551: dataIn1 = 32'd4244
; 
32'd147552: dataIn1 = 32'd4248
; 
32'd147553: dataIn1 = 32'd4249
; 
32'd147554: dataIn1 = 32'd171
; 
32'd147555: dataIn1 = 32'd2390
; 
32'd147556: dataIn1 = 32'd3219
; 
32'd147557: dataIn1 = 32'd4244
; 
32'd147558: dataIn1 = 32'd4248
; 
32'd147559: dataIn1 = 32'd4249
; 
32'd147560: dataIn1 = 32'd4259
; 
32'd147561: dataIn1 = 32'd2393
; 
32'd147562: dataIn1 = 32'd2394
; 
32'd147563: dataIn1 = 32'd4250
; 
32'd147564: dataIn1 = 32'd4251
; 
32'd147565: dataIn1 = 32'd4252
; 
32'd147566: dataIn1 = 32'd4253
; 
32'd147567: dataIn1 = 32'd4254
; 
32'd147568: dataIn1 = 32'd2392
; 
32'd147569: dataIn1 = 32'd2394
; 
32'd147570: dataIn1 = 32'd4250
; 
32'd147571: dataIn1 = 32'd4251
; 
32'd147572: dataIn1 = 32'd4252
; 
32'd147573: dataIn1 = 32'd4255
; 
32'd147574: dataIn1 = 32'd4256
; 
32'd147575: dataIn1 = 32'd2392
; 
32'd147576: dataIn1 = 32'd2393
; 
32'd147577: dataIn1 = 32'd4250
; 
32'd147578: dataIn1 = 32'd4251
; 
32'd147579: dataIn1 = 32'd4252
; 
32'd147580: dataIn1 = 32'd4257
; 
32'd147581: dataIn1 = 32'd4258
; 
32'd147582: dataIn1 = 32'd475
; 
32'd147583: dataIn1 = 32'd2394
; 
32'd147584: dataIn1 = 32'd4250
; 
32'd147585: dataIn1 = 32'd4253
; 
32'd147586: dataIn1 = 32'd4254
; 
32'd147587: dataIn1 = 32'd5369
; 
32'd147588: dataIn1 = 32'd475
; 
32'd147589: dataIn1 = 32'd2393
; 
32'd147590: dataIn1 = 32'd4250
; 
32'd147591: dataIn1 = 32'd4253
; 
32'd147592: dataIn1 = 32'd4254
; 
32'd147593: dataIn1 = 32'd4262
; 
32'd147594: dataIn1 = 32'd4265
; 
32'd147595: dataIn1 = 32'd474
; 
32'd147596: dataIn1 = 32'd2394
; 
32'd147597: dataIn1 = 32'd4251
; 
32'd147598: dataIn1 = 32'd4255
; 
32'd147599: dataIn1 = 32'd4256
; 
32'd147600: dataIn1 = 32'd5368
; 
32'd147601: dataIn1 = 32'd474
; 
32'd147602: dataIn1 = 32'd2392
; 
32'd147603: dataIn1 = 32'd4247
; 
32'd147604: dataIn1 = 32'd4251
; 
32'd147605: dataIn1 = 32'd4255
; 
32'd147606: dataIn1 = 32'd4256
; 
32'd147607: dataIn1 = 32'd4260
; 
32'd147608: dataIn1 = 32'd333
; 
32'd147609: dataIn1 = 32'd2393
; 
32'd147610: dataIn1 = 32'd3215
; 
32'd147611: dataIn1 = 32'd4252
; 
32'd147612: dataIn1 = 32'd4257
; 
32'd147613: dataIn1 = 32'd4258
; 
32'd147614: dataIn1 = 32'd4264
; 
32'd147615: dataIn1 = 32'd333
; 
32'd147616: dataIn1 = 32'd2392
; 
32'd147617: dataIn1 = 32'd3222
; 
32'd147618: dataIn1 = 32'd4252
; 
32'd147619: dataIn1 = 32'd4257
; 
32'd147620: dataIn1 = 32'd4258
; 
32'd147621: dataIn1 = 32'd4261
; 
32'd147622: dataIn1 = 32'd2002
; 
32'd147623: dataIn1 = 32'd2390
; 
32'd147624: dataIn1 = 32'd3219
; 
32'd147625: dataIn1 = 32'd4249
; 
32'd147626: dataIn1 = 32'd4259
; 
32'd147627: dataIn1 = 32'd4260
; 
32'd147628: dataIn1 = 32'd4261
; 
32'd147629: dataIn1 = 32'd2390
; 
32'd147630: dataIn1 = 32'd2392
; 
32'd147631: dataIn1 = 32'd4247
; 
32'd147632: dataIn1 = 32'd4256
; 
32'd147633: dataIn1 = 32'd4259
; 
32'd147634: dataIn1 = 32'd4260
; 
32'd147635: dataIn1 = 32'd4261
; 
32'd147636: dataIn1 = 32'd2002
; 
32'd147637: dataIn1 = 32'd2392
; 
32'd147638: dataIn1 = 32'd3222
; 
32'd147639: dataIn1 = 32'd4258
; 
32'd147640: dataIn1 = 32'd4259
; 
32'd147641: dataIn1 = 32'd4260
; 
32'd147642: dataIn1 = 32'd4261
; 
32'd147643: dataIn1 = 32'd2393
; 
32'd147644: dataIn1 = 32'd2395
; 
32'd147645: dataIn1 = 32'd4254
; 
32'd147646: dataIn1 = 32'd4262
; 
32'd147647: dataIn1 = 32'd4263
; 
32'd147648: dataIn1 = 32'd4264
; 
32'd147649: dataIn1 = 32'd4265
; 
32'd147650: dataIn1 = 32'd2001
; 
32'd147651: dataIn1 = 32'd2395
; 
32'd147652: dataIn1 = 32'd3214
; 
32'd147653: dataIn1 = 32'd4262
; 
32'd147654: dataIn1 = 32'd4263
; 
32'd147655: dataIn1 = 32'd4264
; 
32'd147656: dataIn1 = 32'd4270
; 
32'd147657: dataIn1 = 32'd2001
; 
32'd147658: dataIn1 = 32'd2393
; 
32'd147659: dataIn1 = 32'd3215
; 
32'd147660: dataIn1 = 32'd4257
; 
32'd147661: dataIn1 = 32'd4262
; 
32'd147662: dataIn1 = 32'd4263
; 
32'd147663: dataIn1 = 32'd4264
; 
32'd147664: dataIn1 = 32'd475
; 
32'd147665: dataIn1 = 32'd2395
; 
32'd147666: dataIn1 = 32'd4254
; 
32'd147667: dataIn1 = 32'd4262
; 
32'd147668: dataIn1 = 32'd4265
; 
32'd147669: dataIn1 = 32'd4266
; 
32'd147670: dataIn1 = 32'd4269
; 
32'd147671: dataIn1 = 32'd2395
; 
32'd147672: dataIn1 = 32'd2397
; 
32'd147673: dataIn1 = 32'd4265
; 
32'd147674: dataIn1 = 32'd4266
; 
32'd147675: dataIn1 = 32'd4267
; 
32'd147676: dataIn1 = 32'd4268
; 
32'd147677: dataIn1 = 32'd4269
; 
32'd147678: dataIn1 = 32'd2395
; 
32'd147679: dataIn1 = 32'd2396
; 
32'd147680: dataIn1 = 32'd4266
; 
32'd147681: dataIn1 = 32'd4267
; 
32'd147682: dataIn1 = 32'd4268
; 
32'd147683: dataIn1 = 32'd4270
; 
32'd147684: dataIn1 = 32'd4271
; 
32'd147685: dataIn1 = 32'd2396
; 
32'd147686: dataIn1 = 32'd2397
; 
32'd147687: dataIn1 = 32'd4266
; 
32'd147688: dataIn1 = 32'd4267
; 
32'd147689: dataIn1 = 32'd4268
; 
32'd147690: dataIn1 = 32'd4272
; 
32'd147691: dataIn1 = 32'd4273
; 
32'd147692: dataIn1 = 32'd475
; 
32'd147693: dataIn1 = 32'd2397
; 
32'd147694: dataIn1 = 32'd4265
; 
32'd147695: dataIn1 = 32'd4266
; 
32'd147696: dataIn1 = 32'd4269
; 
32'd147697: dataIn1 = 32'd5371
; 
32'd147698: dataIn1 = 32'd173
; 
32'd147699: dataIn1 = 32'd2395
; 
32'd147700: dataIn1 = 32'd3214
; 
32'd147701: dataIn1 = 32'd4263
; 
32'd147702: dataIn1 = 32'd4267
; 
32'd147703: dataIn1 = 32'd4270
; 
32'd147704: dataIn1 = 32'd4271
; 
32'd147705: dataIn1 = 32'd173
; 
32'd147706: dataIn1 = 32'd2396
; 
32'd147707: dataIn1 = 32'd3206
; 
32'd147708: dataIn1 = 32'd4267
; 
32'd147709: dataIn1 = 32'd4270
; 
32'd147710: dataIn1 = 32'd4271
; 
32'd147711: dataIn1 = 32'd4284
; 
32'd147712: dataIn1 = 32'd476
; 
32'd147713: dataIn1 = 32'd2397
; 
32'd147714: dataIn1 = 32'd4268
; 
32'd147715: dataIn1 = 32'd4272
; 
32'd147716: dataIn1 = 32'd4273
; 
32'd147717: dataIn1 = 32'd5370
; 
32'd147718: dataIn1 = 32'd476
; 
32'd147719: dataIn1 = 32'd2396
; 
32'd147720: dataIn1 = 32'd4268
; 
32'd147721: dataIn1 = 32'd4272
; 
32'd147722: dataIn1 = 32'd4273
; 
32'd147723: dataIn1 = 32'd4281
; 
32'd147724: dataIn1 = 32'd4285
; 
32'd147725: dataIn1 = 32'd2399
; 
32'd147726: dataIn1 = 32'd2400
; 
32'd147727: dataIn1 = 32'd4274
; 
32'd147728: dataIn1 = 32'd4275
; 
32'd147729: dataIn1 = 32'd4276
; 
32'd147730: dataIn1 = 32'd4277
; 
32'd147731: dataIn1 = 32'd4278
; 
32'd147732: dataIn1 = 32'd2398
; 
32'd147733: dataIn1 = 32'd2400
; 
32'd147734: dataIn1 = 32'd4274
; 
32'd147735: dataIn1 = 32'd4275
; 
32'd147736: dataIn1 = 32'd4276
; 
32'd147737: dataIn1 = 32'd4279
; 
32'd147738: dataIn1 = 32'd4280
; 
32'd147739: dataIn1 = 32'd2398
; 
32'd147740: dataIn1 = 32'd2399
; 
32'd147741: dataIn1 = 32'd4274
; 
32'd147742: dataIn1 = 32'd4275
; 
32'd147743: dataIn1 = 32'd4276
; 
32'd147744: dataIn1 = 32'd4281
; 
32'd147745: dataIn1 = 32'd4282
; 
32'd147746: dataIn1 = 32'd327
; 
32'd147747: dataIn1 = 32'd2400
; 
32'd147748: dataIn1 = 32'd3198
; 
32'd147749: dataIn1 = 32'd4274
; 
32'd147750: dataIn1 = 32'd4277
; 
32'd147751: dataIn1 = 32'd4278
; 
32'd147752: dataIn1 = 32'd4286
; 
32'd147753: dataIn1 = 32'd327
; 
32'd147754: dataIn1 = 32'd2399
; 
32'd147755: dataIn1 = 32'd3205
; 
32'd147756: dataIn1 = 32'd4274
; 
32'd147757: dataIn1 = 32'd4277
; 
32'd147758: dataIn1 = 32'd4278
; 
32'd147759: dataIn1 = 32'd4283
; 
32'd147760: dataIn1 = 32'd477
; 
32'd147761: dataIn1 = 32'd2400
; 
32'd147762: dataIn1 = 32'd4275
; 
32'd147763: dataIn1 = 32'd4279
; 
32'd147764: dataIn1 = 32'd4280
; 
32'd147765: dataIn1 = 32'd4287
; 
32'd147766: dataIn1 = 32'd4289
; 
32'd147767: dataIn1 = 32'd477
; 
32'd147768: dataIn1 = 32'd2398
; 
32'd147769: dataIn1 = 32'd4275
; 
32'd147770: dataIn1 = 32'd4279
; 
32'd147771: dataIn1 = 32'd4280
; 
32'd147772: dataIn1 = 32'd5373
; 
32'd147773: dataIn1 = 32'd476
; 
32'd147774: dataIn1 = 32'd2399
; 
32'd147775: dataIn1 = 32'd4273
; 
32'd147776: dataIn1 = 32'd4276
; 
32'd147777: dataIn1 = 32'd4281
; 
32'd147778: dataIn1 = 32'd4282
; 
32'd147779: dataIn1 = 32'd4285
; 
32'd147780: dataIn1 = 32'd476
; 
32'd147781: dataIn1 = 32'd2398
; 
32'd147782: dataIn1 = 32'd4276
; 
32'd147783: dataIn1 = 32'd4281
; 
32'd147784: dataIn1 = 32'd4282
; 
32'd147785: dataIn1 = 32'd5372
; 
32'd147786: dataIn1 = 32'd2000
; 
32'd147787: dataIn1 = 32'd2399
; 
32'd147788: dataIn1 = 32'd3205
; 
32'd147789: dataIn1 = 32'd4278
; 
32'd147790: dataIn1 = 32'd4283
; 
32'd147791: dataIn1 = 32'd4284
; 
32'd147792: dataIn1 = 32'd4285
; 
32'd147793: dataIn1 = 32'd2000
; 
32'd147794: dataIn1 = 32'd2396
; 
32'd147795: dataIn1 = 32'd3206
; 
32'd147796: dataIn1 = 32'd4271
; 
32'd147797: dataIn1 = 32'd4283
; 
32'd147798: dataIn1 = 32'd4284
; 
32'd147799: dataIn1 = 32'd4285
; 
32'd147800: dataIn1 = 32'd2396
; 
32'd147801: dataIn1 = 32'd2399
; 
32'd147802: dataIn1 = 32'd4273
; 
32'd147803: dataIn1 = 32'd4281
; 
32'd147804: dataIn1 = 32'd4283
; 
32'd147805: dataIn1 = 32'd4284
; 
32'd147806: dataIn1 = 32'd4285
; 
32'd147807: dataIn1 = 32'd1999
; 
32'd147808: dataIn1 = 32'd2400
; 
32'd147809: dataIn1 = 32'd3198
; 
32'd147810: dataIn1 = 32'd4277
; 
32'd147811: dataIn1 = 32'd4286
; 
32'd147812: dataIn1 = 32'd4287
; 
32'd147813: dataIn1 = 32'd4288
; 
32'd147814: dataIn1 = 32'd2400
; 
32'd147815: dataIn1 = 32'd2401
; 
32'd147816: dataIn1 = 32'd4279
; 
32'd147817: dataIn1 = 32'd4286
; 
32'd147818: dataIn1 = 32'd4287
; 
32'd147819: dataIn1 = 32'd4288
; 
32'd147820: dataIn1 = 32'd4289
; 
32'd147821: dataIn1 = 32'd1999
; 
32'd147822: dataIn1 = 32'd2401
; 
32'd147823: dataIn1 = 32'd3201
; 
32'd147824: dataIn1 = 32'd4286
; 
32'd147825: dataIn1 = 32'd4287
; 
32'd147826: dataIn1 = 32'd4288
; 
32'd147827: dataIn1 = 32'd4297
; 
32'd147828: dataIn1 = 32'd477
; 
32'd147829: dataIn1 = 32'd2401
; 
32'd147830: dataIn1 = 32'd4279
; 
32'd147831: dataIn1 = 32'd4287
; 
32'd147832: dataIn1 = 32'd4289
; 
32'd147833: dataIn1 = 32'd4291
; 
32'd147834: dataIn1 = 32'd4295
; 
32'd147835: dataIn1 = 32'd2402
; 
32'd147836: dataIn1 = 32'd2403
; 
32'd147837: dataIn1 = 32'd4290
; 
32'd147838: dataIn1 = 32'd4291
; 
32'd147839: dataIn1 = 32'd4292
; 
32'd147840: dataIn1 = 32'd4293
; 
32'd147841: dataIn1 = 32'd4294
; 
32'd147842: dataIn1 = 32'd2401
; 
32'd147843: dataIn1 = 32'd2403
; 
32'd147844: dataIn1 = 32'd4289
; 
32'd147845: dataIn1 = 32'd4290
; 
32'd147846: dataIn1 = 32'd4291
; 
32'd147847: dataIn1 = 32'd4292
; 
32'd147848: dataIn1 = 32'd4295
; 
32'd147849: dataIn1 = 32'd2401
; 
32'd147850: dataIn1 = 32'd2402
; 
32'd147851: dataIn1 = 32'd4290
; 
32'd147852: dataIn1 = 32'd4291
; 
32'd147853: dataIn1 = 32'd4292
; 
32'd147854: dataIn1 = 32'd4296
; 
32'd147855: dataIn1 = 32'd4297
; 
32'd147856: dataIn1 = 32'd478
; 
32'd147857: dataIn1 = 32'd2403
; 
32'd147858: dataIn1 = 32'd4290
; 
32'd147859: dataIn1 = 32'd4293
; 
32'd147860: dataIn1 = 32'd4294
; 
32'd147861: dataIn1 = 32'd5375
; 
32'd147862: dataIn1 = 32'd478
; 
32'd147863: dataIn1 = 32'd2402
; 
32'd147864: dataIn1 = 32'd4290
; 
32'd147865: dataIn1 = 32'd4293
; 
32'd147866: dataIn1 = 32'd4294
; 
32'd147867: dataIn1 = 32'd4301
; 
32'd147868: dataIn1 = 32'd4311
; 
32'd147869: dataIn1 = 32'd477
; 
32'd147870: dataIn1 = 32'd2403
; 
32'd147871: dataIn1 = 32'd4289
; 
32'd147872: dataIn1 = 32'd4291
; 
32'd147873: dataIn1 = 32'd4295
; 
32'd147874: dataIn1 = 32'd5374
; 
32'd147875: dataIn1 = 32'd174
; 
32'd147876: dataIn1 = 32'd2402
; 
32'd147877: dataIn1 = 32'd3229
; 
32'd147878: dataIn1 = 32'd4292
; 
32'd147879: dataIn1 = 32'd4296
; 
32'd147880: dataIn1 = 32'd4297
; 
32'd147881: dataIn1 = 32'd4313
; 
32'd147882: dataIn1 = 32'd174
; 
32'd147883: dataIn1 = 32'd2401
; 
32'd147884: dataIn1 = 32'd3201
; 
32'd147885: dataIn1 = 32'd4288
; 
32'd147886: dataIn1 = 32'd4292
; 
32'd147887: dataIn1 = 32'd4296
; 
32'd147888: dataIn1 = 32'd4297
; 
32'd147889: dataIn1 = 32'd2405
; 
32'd147890: dataIn1 = 32'd2406
; 
32'd147891: dataIn1 = 32'd4298
; 
32'd147892: dataIn1 = 32'd4299
; 
32'd147893: dataIn1 = 32'd4300
; 
32'd147894: dataIn1 = 32'd4301
; 
32'd147895: dataIn1 = 32'd4302
; 
32'd147896: dataIn1 = 32'd2404
; 
32'd147897: dataIn1 = 32'd2406
; 
32'd147898: dataIn1 = 32'd4298
; 
32'd147899: dataIn1 = 32'd4299
; 
32'd147900: dataIn1 = 32'd4300
; 
32'd147901: dataIn1 = 32'd4303
; 
32'd147902: dataIn1 = 32'd4304
; 
32'd147903: dataIn1 = 32'd2404
; 
32'd147904: dataIn1 = 32'd2405
; 
32'd147905: dataIn1 = 32'd4298
; 
32'd147906: dataIn1 = 32'd4299
; 
32'd147907: dataIn1 = 32'd4300
; 
32'd147908: dataIn1 = 32'd4305
; 
32'd147909: dataIn1 = 32'd4306
; 
32'd147910: dataIn1 = 32'd478
; 
32'd147911: dataIn1 = 32'd2406
; 
32'd147912: dataIn1 = 32'd4294
; 
32'd147913: dataIn1 = 32'd4298
; 
32'd147914: dataIn1 = 32'd4301
; 
32'd147915: dataIn1 = 32'd4302
; 
32'd147916: dataIn1 = 32'd4311
; 
32'd147917: dataIn1 = 32'd478
; 
32'd147918: dataIn1 = 32'd2405
; 
32'd147919: dataIn1 = 32'd4298
; 
32'd147920: dataIn1 = 32'd4301
; 
32'd147921: dataIn1 = 32'd4302
; 
32'd147922: dataIn1 = 32'd5377
; 
32'd147923: dataIn1 = 32'd334
; 
32'd147924: dataIn1 = 32'd2406
; 
32'd147925: dataIn1 = 32'd3228
; 
32'd147926: dataIn1 = 32'd4299
; 
32'd147927: dataIn1 = 32'd4303
; 
32'd147928: dataIn1 = 32'd4304
; 
32'd147929: dataIn1 = 32'd4312
; 
32'd147930: dataIn1 = 32'd334
; 
32'd147931: dataIn1 = 32'd2404
; 
32'd147932: dataIn1 = 32'd3234
; 
32'd147933: dataIn1 = 32'd4299
; 
32'd147934: dataIn1 = 32'd4303
; 
32'd147935: dataIn1 = 32'd4304
; 
32'd147936: dataIn1 = 32'd4308
; 
32'd147937: dataIn1 = 32'd479
; 
32'd147938: dataIn1 = 32'd2405
; 
32'd147939: dataIn1 = 32'd4300
; 
32'd147940: dataIn1 = 32'd4305
; 
32'd147941: dataIn1 = 32'd4306
; 
32'd147942: dataIn1 = 32'd5376
; 
32'd147943: dataIn1 = 32'd479
; 
32'd147944: dataIn1 = 32'd2404
; 
32'd147945: dataIn1 = 32'd4300
; 
32'd147946: dataIn1 = 32'd4305
; 
32'd147947: dataIn1 = 32'd4306
; 
32'd147948: dataIn1 = 32'd4309
; 
32'd147949: dataIn1 = 32'd4310
; 
32'd147950: dataIn1 = 32'd2004
; 
32'd147951: dataIn1 = 32'd2407
; 
32'd147952: dataIn1 = 32'd3233
; 
32'd147953: dataIn1 = 32'd4307
; 
32'd147954: dataIn1 = 32'd4308
; 
32'd147955: dataIn1 = 32'd4309
; 
32'd147956: dataIn1 = 32'd4317
; 
32'd147957: dataIn1 = 32'd2004
; 
32'd147958: dataIn1 = 32'd2404
; 
32'd147959: dataIn1 = 32'd3234
; 
32'd147960: dataIn1 = 32'd4304
; 
32'd147961: dataIn1 = 32'd4307
; 
32'd147962: dataIn1 = 32'd4308
; 
32'd147963: dataIn1 = 32'd4309
; 
32'd147964: dataIn1 = 32'd2404
; 
32'd147965: dataIn1 = 32'd2407
; 
32'd147966: dataIn1 = 32'd4306
; 
32'd147967: dataIn1 = 32'd4307
; 
32'd147968: dataIn1 = 32'd4308
; 
32'd147969: dataIn1 = 32'd4309
; 
32'd147970: dataIn1 = 32'd4310
; 
32'd147971: dataIn1 = 32'd479
; 
32'd147972: dataIn1 = 32'd2407
; 
32'd147973: dataIn1 = 32'd4306
; 
32'd147974: dataIn1 = 32'd4309
; 
32'd147975: dataIn1 = 32'd4310
; 
32'd147976: dataIn1 = 32'd4315
; 
32'd147977: dataIn1 = 32'd4319
; 
32'd147978: dataIn1 = 32'd2402
; 
32'd147979: dataIn1 = 32'd2406
; 
32'd147980: dataIn1 = 32'd4294
; 
32'd147981: dataIn1 = 32'd4301
; 
32'd147982: dataIn1 = 32'd4311
; 
32'd147983: dataIn1 = 32'd4312
; 
32'd147984: dataIn1 = 32'd4313
; 
32'd147985: dataIn1 = 32'd2003
; 
32'd147986: dataIn1 = 32'd2406
; 
32'd147987: dataIn1 = 32'd3228
; 
32'd147988: dataIn1 = 32'd4303
; 
32'd147989: dataIn1 = 32'd4311
; 
32'd147990: dataIn1 = 32'd4312
; 
32'd147991: dataIn1 = 32'd4313
; 
32'd147992: dataIn1 = 32'd2003
; 
32'd147993: dataIn1 = 32'd2402
; 
32'd147994: dataIn1 = 32'd3229
; 
32'd147995: dataIn1 = 32'd4296
; 
32'd147996: dataIn1 = 32'd4311
; 
32'd147997: dataIn1 = 32'd4312
; 
32'd147998: dataIn1 = 32'd4313
; 
32'd147999: dataIn1 = 32'd2407
; 
32'd148000: dataIn1 = 32'd2409
; 
32'd148001: dataIn1 = 32'd4314
; 
32'd148002: dataIn1 = 32'd4315
; 
32'd148003: dataIn1 = 32'd4316
; 
32'd148004: dataIn1 = 32'd4317
; 
32'd148005: dataIn1 = 32'd4318
; 
32'd148006: dataIn1 = 32'd2407
; 
32'd148007: dataIn1 = 32'd2408
; 
32'd148008: dataIn1 = 32'd4310
; 
32'd148009: dataIn1 = 32'd4314
; 
32'd148010: dataIn1 = 32'd4315
; 
32'd148011: dataIn1 = 32'd4316
; 
32'd148012: dataIn1 = 32'd4319
; 
32'd148013: dataIn1 = 32'd2408
; 
32'd148014: dataIn1 = 32'd2409
; 
32'd148015: dataIn1 = 32'd4314
; 
32'd148016: dataIn1 = 32'd4315
; 
32'd148017: dataIn1 = 32'd4316
; 
32'd148018: dataIn1 = 32'd4320
; 
32'd148019: dataIn1 = 32'd4321
; 
32'd148020: dataIn1 = 32'd175
; 
32'd148021: dataIn1 = 32'd2407
; 
32'd148022: dataIn1 = 32'd3233
; 
32'd148023: dataIn1 = 32'd4307
; 
32'd148024: dataIn1 = 32'd4314
; 
32'd148025: dataIn1 = 32'd4317
; 
32'd148026: dataIn1 = 32'd4318
; 
32'd148027: dataIn1 = 32'd175
; 
32'd148028: dataIn1 = 32'd2409
; 
32'd148029: dataIn1 = 32'd3240
; 
32'd148030: dataIn1 = 32'd4314
; 
32'd148031: dataIn1 = 32'd4317
; 
32'd148032: dataIn1 = 32'd4318
; 
32'd148033: dataIn1 = 32'd4331
; 
32'd148034: dataIn1 = 32'd479
; 
32'd148035: dataIn1 = 32'd2408
; 
32'd148036: dataIn1 = 32'd4310
; 
32'd148037: dataIn1 = 32'd4315
; 
32'd148038: dataIn1 = 32'd4319
; 
32'd148039: dataIn1 = 32'd5379
; 
32'd148040: dataIn1 = 32'd480
; 
32'd148041: dataIn1 = 32'd2409
; 
32'd148042: dataIn1 = 32'd4316
; 
32'd148043: dataIn1 = 32'd4320
; 
32'd148044: dataIn1 = 32'd4321
; 
32'd148045: dataIn1 = 32'd4330
; 
32'd148046: dataIn1 = 32'd4333
; 
32'd148047: dataIn1 = 32'd480
; 
32'd148048: dataIn1 = 32'd2408
; 
32'd148049: dataIn1 = 32'd4316
; 
32'd148050: dataIn1 = 32'd4320
; 
32'd148051: dataIn1 = 32'd4321
; 
32'd148052: dataIn1 = 32'd5378
; 
32'd148053: dataIn1 = 32'd2411
; 
32'd148054: dataIn1 = 32'd2412
; 
32'd148055: dataIn1 = 32'd4322
; 
32'd148056: dataIn1 = 32'd4323
; 
32'd148057: dataIn1 = 32'd4324
; 
32'd148058: dataIn1 = 32'd4325
; 
32'd148059: dataIn1 = 32'd4326
; 
32'd148060: dataIn1 = 32'd2410
; 
32'd148061: dataIn1 = 32'd2412
; 
32'd148062: dataIn1 = 32'd4322
; 
32'd148063: dataIn1 = 32'd4323
; 
32'd148064: dataIn1 = 32'd4324
; 
32'd148065: dataIn1 = 32'd4327
; 
32'd148066: dataIn1 = 32'd4328
; 
32'd148067: dataIn1 = 32'd2410
; 
32'd148068: dataIn1 = 32'd2411
; 
32'd148069: dataIn1 = 32'd4322
; 
32'd148070: dataIn1 = 32'd4323
; 
32'd148071: dataIn1 = 32'd4324
; 
32'd148072: dataIn1 = 32'd4329
; 
32'd148073: dataIn1 = 32'd4330
; 
32'd148074: dataIn1 = 32'd481
; 
32'd148075: dataIn1 = 32'd2412
; 
32'd148076: dataIn1 = 32'd4322
; 
32'd148077: dataIn1 = 32'd4325
; 
32'd148078: dataIn1 = 32'd4326
; 
32'd148079: dataIn1 = 32'd4334
; 
32'd148080: dataIn1 = 32'd4337
; 
32'd148081: dataIn1 = 32'd481
; 
32'd148082: dataIn1 = 32'd2411
; 
32'd148083: dataIn1 = 32'd4322
; 
32'd148084: dataIn1 = 32'd4325
; 
32'd148085: dataIn1 = 32'd4326
; 
32'd148086: dataIn1 = 32'd5381
; 
32'd148087: dataIn1 = 32'd341
; 
32'd148088: dataIn1 = 32'd2412
; 
32'd148089: dataIn1 = 32'd3249
; 
32'd148090: dataIn1 = 32'd4323
; 
32'd148091: dataIn1 = 32'd4327
; 
32'd148092: dataIn1 = 32'd4328
; 
32'd148093: dataIn1 = 32'd4335
; 
32'd148094: dataIn1 = 32'd341
; 
32'd148095: dataIn1 = 32'd2410
; 
32'd148096: dataIn1 = 32'd3241
; 
32'd148097: dataIn1 = 32'd4323
; 
32'd148098: dataIn1 = 32'd4327
; 
32'd148099: dataIn1 = 32'd4328
; 
32'd148100: dataIn1 = 32'd4332
; 
32'd148101: dataIn1 = 32'd480
; 
32'd148102: dataIn1 = 32'd2411
; 
32'd148103: dataIn1 = 32'd4324
; 
32'd148104: dataIn1 = 32'd4329
; 
32'd148105: dataIn1 = 32'd4330
; 
32'd148106: dataIn1 = 32'd5380
; 
32'd148107: dataIn1 = 32'd480
; 
32'd148108: dataIn1 = 32'd2410
; 
32'd148109: dataIn1 = 32'd4320
; 
32'd148110: dataIn1 = 32'd4324
; 
32'd148111: dataIn1 = 32'd4329
; 
32'd148112: dataIn1 = 32'd4330
; 
32'd148113: dataIn1 = 32'd4333
; 
32'd148114: dataIn1 = 32'd2005
; 
32'd148115: dataIn1 = 32'd2409
; 
32'd148116: dataIn1 = 32'd3240
; 
32'd148117: dataIn1 = 32'd4318
; 
32'd148118: dataIn1 = 32'd4331
; 
32'd148119: dataIn1 = 32'd4332
; 
32'd148120: dataIn1 = 32'd4333
; 
32'd148121: dataIn1 = 32'd2005
; 
32'd148122: dataIn1 = 32'd2410
; 
32'd148123: dataIn1 = 32'd3241
; 
32'd148124: dataIn1 = 32'd4328
; 
32'd148125: dataIn1 = 32'd4331
; 
32'd148126: dataIn1 = 32'd4332
; 
32'd148127: dataIn1 = 32'd4333
; 
32'd148128: dataIn1 = 32'd2409
; 
32'd148129: dataIn1 = 32'd2410
; 
32'd148130: dataIn1 = 32'd4320
; 
32'd148131: dataIn1 = 32'd4330
; 
32'd148132: dataIn1 = 32'd4331
; 
32'd148133: dataIn1 = 32'd4332
; 
32'd148134: dataIn1 = 32'd4333
; 
32'd148135: dataIn1 = 32'd2412
; 
32'd148136: dataIn1 = 32'd2413
; 
32'd148137: dataIn1 = 32'd4325
; 
32'd148138: dataIn1 = 32'd4334
; 
32'd148139: dataIn1 = 32'd4335
; 
32'd148140: dataIn1 = 32'd4336
; 
32'd148141: dataIn1 = 32'd4337
; 
32'd148142: dataIn1 = 32'd2006
; 
32'd148143: dataIn1 = 32'd2412
; 
32'd148144: dataIn1 = 32'd3249
; 
32'd148145: dataIn1 = 32'd4327
; 
32'd148146: dataIn1 = 32'd4334
; 
32'd148147: dataIn1 = 32'd4335
; 
32'd148148: dataIn1 = 32'd4336
; 
32'd148149: dataIn1 = 32'd2006
; 
32'd148150: dataIn1 = 32'd2413
; 
32'd148151: dataIn1 = 32'd3250
; 
32'd148152: dataIn1 = 32'd4334
; 
32'd148153: dataIn1 = 32'd4335
; 
32'd148154: dataIn1 = 32'd4336
; 
32'd148155: dataIn1 = 32'd4344
; 
32'd148156: dataIn1 = 32'd481
; 
32'd148157: dataIn1 = 32'd2413
; 
32'd148158: dataIn1 = 32'd4325
; 
32'd148159: dataIn1 = 32'd4334
; 
32'd148160: dataIn1 = 32'd4337
; 
32'd148161: dataIn1 = 32'd4338
; 
32'd148162: dataIn1 = 32'd4341
; 
32'd148163: dataIn1 = 32'd2413
; 
32'd148164: dataIn1 = 32'd2415
; 
32'd148165: dataIn1 = 32'd4337
; 
32'd148166: dataIn1 = 32'd4338
; 
32'd148167: dataIn1 = 32'd4339
; 
32'd148168: dataIn1 = 32'd4340
; 
32'd148169: dataIn1 = 32'd4341
; 
32'd148170: dataIn1 = 32'd2414
; 
32'd148171: dataIn1 = 32'd2415
; 
32'd148172: dataIn1 = 32'd4338
; 
32'd148173: dataIn1 = 32'd4339
; 
32'd148174: dataIn1 = 32'd4340
; 
32'd148175: dataIn1 = 32'd4342
; 
32'd148176: dataIn1 = 32'd4343
; 
32'd148177: dataIn1 = 32'd2413
; 
32'd148178: dataIn1 = 32'd2414
; 
32'd148179: dataIn1 = 32'd4338
; 
32'd148180: dataIn1 = 32'd4339
; 
32'd148181: dataIn1 = 32'd4340
; 
32'd148182: dataIn1 = 32'd4344
; 
32'd148183: dataIn1 = 32'd4345
; 
32'd148184: dataIn1 = 32'd481
; 
32'd148185: dataIn1 = 32'd2415
; 
32'd148186: dataIn1 = 32'd4337
; 
32'd148187: dataIn1 = 32'd4338
; 
32'd148188: dataIn1 = 32'd4341
; 
32'd148189: dataIn1 = 32'd5383
; 
32'd148190: dataIn1 = 32'd482
; 
32'd148191: dataIn1 = 32'd2415
; 
32'd148192: dataIn1 = 32'd4339
; 
32'd148193: dataIn1 = 32'd4342
; 
32'd148194: dataIn1 = 32'd4343
; 
32'd148195: dataIn1 = 32'd5382
; 
32'd148196: dataIn1 = 32'd482
; 
32'd148197: dataIn1 = 32'd2414
; 
32'd148198: dataIn1 = 32'd4339
; 
32'd148199: dataIn1 = 32'd4342
; 
32'd148200: dataIn1 = 32'd4343
; 
32'd148201: dataIn1 = 32'd4352
; 
32'd148202: dataIn1 = 32'd4356
; 
32'd148203: dataIn1 = 32'd177
; 
32'd148204: dataIn1 = 32'd2413
; 
32'd148205: dataIn1 = 32'd3250
; 
32'd148206: dataIn1 = 32'd4336
; 
32'd148207: dataIn1 = 32'd4340
; 
32'd148208: dataIn1 = 32'd4344
; 
32'd148209: dataIn1 = 32'd4345
; 
32'd148210: dataIn1 = 32'd177
; 
32'd148211: dataIn1 = 32'd2414
; 
32'd148212: dataIn1 = 32'd3275
; 
32'd148213: dataIn1 = 32'd4340
; 
32'd148214: dataIn1 = 32'd4344
; 
32'd148215: dataIn1 = 32'd4345
; 
32'd148216: dataIn1 = 32'd4355
; 
32'd148217: dataIn1 = 32'd2417
; 
32'd148218: dataIn1 = 32'd2418
; 
32'd148219: dataIn1 = 32'd4346
; 
32'd148220: dataIn1 = 32'd4347
; 
32'd148221: dataIn1 = 32'd4348
; 
32'd148222: dataIn1 = 32'd4349
; 
32'd148223: dataIn1 = 32'd4350
; 
32'd148224: dataIn1 = 32'd2416
; 
32'd148225: dataIn1 = 32'd2418
; 
32'd148226: dataIn1 = 32'd4346
; 
32'd148227: dataIn1 = 32'd4347
; 
32'd148228: dataIn1 = 32'd4348
; 
32'd148229: dataIn1 = 32'd4351
; 
32'd148230: dataIn1 = 32'd4352
; 
32'd148231: dataIn1 = 32'd2416
; 
32'd148232: dataIn1 = 32'd2417
; 
32'd148233: dataIn1 = 32'd4346
; 
32'd148234: dataIn1 = 32'd4347
; 
32'd148235: dataIn1 = 32'd4348
; 
32'd148236: dataIn1 = 32'd4353
; 
32'd148237: dataIn1 = 32'd4354
; 
32'd148238: dataIn1 = 32'd483
; 
32'd148239: dataIn1 = 32'd2418
; 
32'd148240: dataIn1 = 32'd4346
; 
32'd148241: dataIn1 = 32'd4349
; 
32'd148242: dataIn1 = 32'd4350
; 
32'd148243: dataIn1 = 32'd5385
; 
32'd148244: dataIn1 = 32'd483
; 
32'd148245: dataIn1 = 32'd2417
; 
32'd148246: dataIn1 = 32'd4346
; 
32'd148247: dataIn1 = 32'd4349
; 
32'd148248: dataIn1 = 32'd4350
; 
32'd148249: dataIn1 = 32'd4358
; 
32'd148250: dataIn1 = 32'd4361
; 
32'd148251: dataIn1 = 32'd482
; 
32'd148252: dataIn1 = 32'd2418
; 
32'd148253: dataIn1 = 32'd4347
; 
32'd148254: dataIn1 = 32'd4351
; 
32'd148255: dataIn1 = 32'd4352
; 
32'd148256: dataIn1 = 32'd5384
; 
32'd148257: dataIn1 = 32'd482
; 
32'd148258: dataIn1 = 32'd2416
; 
32'd148259: dataIn1 = 32'd4343
; 
32'd148260: dataIn1 = 32'd4347
; 
32'd148261: dataIn1 = 32'd4351
; 
32'd148262: dataIn1 = 32'd4352
; 
32'd148263: dataIn1 = 32'd4356
; 
32'd148264: dataIn1 = 32'd349
; 
32'd148265: dataIn1 = 32'd2417
; 
32'd148266: dataIn1 = 32'd3271
; 
32'd148267: dataIn1 = 32'd4348
; 
32'd148268: dataIn1 = 32'd4353
; 
32'd148269: dataIn1 = 32'd4354
; 
32'd148270: dataIn1 = 32'd4360
; 
32'd148271: dataIn1 = 32'd349
; 
32'd148272: dataIn1 = 32'd2416
; 
32'd148273: dataIn1 = 32'd3278
; 
32'd148274: dataIn1 = 32'd4348
; 
32'd148275: dataIn1 = 32'd4353
; 
32'd148276: dataIn1 = 32'd4354
; 
32'd148277: dataIn1 = 32'd4357
; 
32'd148278: dataIn1 = 32'd2010
; 
32'd148279: dataIn1 = 32'd2414
; 
32'd148280: dataIn1 = 32'd3275
; 
32'd148281: dataIn1 = 32'd4345
; 
32'd148282: dataIn1 = 32'd4355
; 
32'd148283: dataIn1 = 32'd4356
; 
32'd148284: dataIn1 = 32'd4357
; 
32'd148285: dataIn1 = 32'd2414
; 
32'd148286: dataIn1 = 32'd2416
; 
32'd148287: dataIn1 = 32'd4343
; 
32'd148288: dataIn1 = 32'd4352
; 
32'd148289: dataIn1 = 32'd4355
; 
32'd148290: dataIn1 = 32'd4356
; 
32'd148291: dataIn1 = 32'd4357
; 
32'd148292: dataIn1 = 32'd2010
; 
32'd148293: dataIn1 = 32'd2416
; 
32'd148294: dataIn1 = 32'd3278
; 
32'd148295: dataIn1 = 32'd4354
; 
32'd148296: dataIn1 = 32'd4355
; 
32'd148297: dataIn1 = 32'd4356
; 
32'd148298: dataIn1 = 32'd4357
; 
32'd148299: dataIn1 = 32'd2417
; 
32'd148300: dataIn1 = 32'd2419
; 
32'd148301: dataIn1 = 32'd4350
; 
32'd148302: dataIn1 = 32'd4358
; 
32'd148303: dataIn1 = 32'd4359
; 
32'd148304: dataIn1 = 32'd4360
; 
32'd148305: dataIn1 = 32'd4361
; 
32'd148306: dataIn1 = 32'd2009
; 
32'd148307: dataIn1 = 32'd2419
; 
32'd148308: dataIn1 = 32'd3270
; 
32'd148309: dataIn1 = 32'd4358
; 
32'd148310: dataIn1 = 32'd4359
; 
32'd148311: dataIn1 = 32'd4360
; 
32'd148312: dataIn1 = 32'd4366
; 
32'd148313: dataIn1 = 32'd2009
; 
32'd148314: dataIn1 = 32'd2417
; 
32'd148315: dataIn1 = 32'd3271
; 
32'd148316: dataIn1 = 32'd4353
; 
32'd148317: dataIn1 = 32'd4358
; 
32'd148318: dataIn1 = 32'd4359
; 
32'd148319: dataIn1 = 32'd4360
; 
32'd148320: dataIn1 = 32'd483
; 
32'd148321: dataIn1 = 32'd2419
; 
32'd148322: dataIn1 = 32'd4350
; 
32'd148323: dataIn1 = 32'd4358
; 
32'd148324: dataIn1 = 32'd4361
; 
32'd148325: dataIn1 = 32'd4362
; 
32'd148326: dataIn1 = 32'd4365
; 
32'd148327: dataIn1 = 32'd2419
; 
32'd148328: dataIn1 = 32'd2421
; 
32'd148329: dataIn1 = 32'd4361
; 
32'd148330: dataIn1 = 32'd4362
; 
32'd148331: dataIn1 = 32'd4363
; 
32'd148332: dataIn1 = 32'd4364
; 
32'd148333: dataIn1 = 32'd4365
; 
32'd148334: dataIn1 = 32'd2419
; 
32'd148335: dataIn1 = 32'd2420
; 
32'd148336: dataIn1 = 32'd4362
; 
32'd148337: dataIn1 = 32'd4363
; 
32'd148338: dataIn1 = 32'd4364
; 
32'd148339: dataIn1 = 32'd4366
; 
32'd148340: dataIn1 = 32'd4367
; 
32'd148341: dataIn1 = 32'd2420
; 
32'd148342: dataIn1 = 32'd2421
; 
32'd148343: dataIn1 = 32'd4362
; 
32'd148344: dataIn1 = 32'd4363
; 
32'd148345: dataIn1 = 32'd4364
; 
32'd148346: dataIn1 = 32'd4368
; 
32'd148347: dataIn1 = 32'd4369
; 
32'd148348: dataIn1 = 32'd483
; 
32'd148349: dataIn1 = 32'd2421
; 
32'd148350: dataIn1 = 32'd4361
; 
32'd148351: dataIn1 = 32'd4362
; 
32'd148352: dataIn1 = 32'd4365
; 
32'd148353: dataIn1 = 32'd5387
; 
32'd148354: dataIn1 = 32'd179
; 
32'd148355: dataIn1 = 32'd2419
; 
32'd148356: dataIn1 = 32'd3270
; 
32'd148357: dataIn1 = 32'd4359
; 
32'd148358: dataIn1 = 32'd4363
; 
32'd148359: dataIn1 = 32'd4366
; 
32'd148360: dataIn1 = 32'd4367
; 
32'd148361: dataIn1 = 32'd179
; 
32'd148362: dataIn1 = 32'd2420
; 
32'd148363: dataIn1 = 32'd3262
; 
32'd148364: dataIn1 = 32'd4363
; 
32'd148365: dataIn1 = 32'd4366
; 
32'd148366: dataIn1 = 32'd4367
; 
32'd148367: dataIn1 = 32'd4380
; 
32'd148368: dataIn1 = 32'd484
; 
32'd148369: dataIn1 = 32'd2421
; 
32'd148370: dataIn1 = 32'd4364
; 
32'd148371: dataIn1 = 32'd4368
; 
32'd148372: dataIn1 = 32'd4369
; 
32'd148373: dataIn1 = 32'd5386
; 
32'd148374: dataIn1 = 32'd484
; 
32'd148375: dataIn1 = 32'd2420
; 
32'd148376: dataIn1 = 32'd4364
; 
32'd148377: dataIn1 = 32'd4368
; 
32'd148378: dataIn1 = 32'd4369
; 
32'd148379: dataIn1 = 32'd4377
; 
32'd148380: dataIn1 = 32'd4381
; 
32'd148381: dataIn1 = 32'd2423
; 
32'd148382: dataIn1 = 32'd2424
; 
32'd148383: dataIn1 = 32'd4370
; 
32'd148384: dataIn1 = 32'd4371
; 
32'd148385: dataIn1 = 32'd4372
; 
32'd148386: dataIn1 = 32'd4373
; 
32'd148387: dataIn1 = 32'd4374
; 
32'd148388: dataIn1 = 32'd2422
; 
32'd148389: dataIn1 = 32'd2424
; 
32'd148390: dataIn1 = 32'd4370
; 
32'd148391: dataIn1 = 32'd4371
; 
32'd148392: dataIn1 = 32'd4372
; 
32'd148393: dataIn1 = 32'd4375
; 
32'd148394: dataIn1 = 32'd4376
; 
32'd148395: dataIn1 = 32'd2422
; 
32'd148396: dataIn1 = 32'd2423
; 
32'd148397: dataIn1 = 32'd4370
; 
32'd148398: dataIn1 = 32'd4371
; 
32'd148399: dataIn1 = 32'd4372
; 
32'd148400: dataIn1 = 32'd4377
; 
32'd148401: dataIn1 = 32'd4378
; 
32'd148402: dataIn1 = 32'd343
; 
32'd148403: dataIn1 = 32'd2424
; 
32'd148404: dataIn1 = 32'd3254
; 
32'd148405: dataIn1 = 32'd4370
; 
32'd148406: dataIn1 = 32'd4373
; 
32'd148407: dataIn1 = 32'd4374
; 
32'd148408: dataIn1 = 32'd4382
; 
32'd148409: dataIn1 = 32'd343
; 
32'd148410: dataIn1 = 32'd2423
; 
32'd148411: dataIn1 = 32'd3261
; 
32'd148412: dataIn1 = 32'd4370
; 
32'd148413: dataIn1 = 32'd4373
; 
32'd148414: dataIn1 = 32'd4374
; 
32'd148415: dataIn1 = 32'd4379
; 
32'd148416: dataIn1 = 32'd485
; 
32'd148417: dataIn1 = 32'd2424
; 
32'd148418: dataIn1 = 32'd4371
; 
32'd148419: dataIn1 = 32'd4375
; 
32'd148420: dataIn1 = 32'd4376
; 
32'd148421: dataIn1 = 32'd4383
; 
32'd148422: dataIn1 = 32'd4385
; 
32'd148423: dataIn1 = 32'd485
; 
32'd148424: dataIn1 = 32'd2422
; 
32'd148425: dataIn1 = 32'd4371
; 
32'd148426: dataIn1 = 32'd4375
; 
32'd148427: dataIn1 = 32'd4376
; 
32'd148428: dataIn1 = 32'd5389
; 
32'd148429: dataIn1 = 32'd484
; 
32'd148430: dataIn1 = 32'd2423
; 
32'd148431: dataIn1 = 32'd4369
; 
32'd148432: dataIn1 = 32'd4372
; 
32'd148433: dataIn1 = 32'd4377
; 
32'd148434: dataIn1 = 32'd4378
; 
32'd148435: dataIn1 = 32'd4381
; 
32'd148436: dataIn1 = 32'd484
; 
32'd148437: dataIn1 = 32'd2422
; 
32'd148438: dataIn1 = 32'd4372
; 
32'd148439: dataIn1 = 32'd4377
; 
32'd148440: dataIn1 = 32'd4378
; 
32'd148441: dataIn1 = 32'd5388
; 
32'd148442: dataIn1 = 32'd2008
; 
32'd148443: dataIn1 = 32'd2423
; 
32'd148444: dataIn1 = 32'd3261
; 
32'd148445: dataIn1 = 32'd4374
; 
32'd148446: dataIn1 = 32'd4379
; 
32'd148447: dataIn1 = 32'd4380
; 
32'd148448: dataIn1 = 32'd4381
; 
32'd148449: dataIn1 = 32'd2008
; 
32'd148450: dataIn1 = 32'd2420
; 
32'd148451: dataIn1 = 32'd3262
; 
32'd148452: dataIn1 = 32'd4367
; 
32'd148453: dataIn1 = 32'd4379
; 
32'd148454: dataIn1 = 32'd4380
; 
32'd148455: dataIn1 = 32'd4381
; 
32'd148456: dataIn1 = 32'd2420
; 
32'd148457: dataIn1 = 32'd2423
; 
32'd148458: dataIn1 = 32'd4369
; 
32'd148459: dataIn1 = 32'd4377
; 
32'd148460: dataIn1 = 32'd4379
; 
32'd148461: dataIn1 = 32'd4380
; 
32'd148462: dataIn1 = 32'd4381
; 
32'd148463: dataIn1 = 32'd2007
; 
32'd148464: dataIn1 = 32'd2424
; 
32'd148465: dataIn1 = 32'd3254
; 
32'd148466: dataIn1 = 32'd4373
; 
32'd148467: dataIn1 = 32'd4382
; 
32'd148468: dataIn1 = 32'd4383
; 
32'd148469: dataIn1 = 32'd4384
; 
32'd148470: dataIn1 = 32'd2424
; 
32'd148471: dataIn1 = 32'd2425
; 
32'd148472: dataIn1 = 32'd4375
; 
32'd148473: dataIn1 = 32'd4382
; 
32'd148474: dataIn1 = 32'd4383
; 
32'd148475: dataIn1 = 32'd4384
; 
32'd148476: dataIn1 = 32'd4385
; 
32'd148477: dataIn1 = 32'd2007
; 
32'd148478: dataIn1 = 32'd2425
; 
32'd148479: dataIn1 = 32'd3257
; 
32'd148480: dataIn1 = 32'd4382
; 
32'd148481: dataIn1 = 32'd4383
; 
32'd148482: dataIn1 = 32'd4384
; 
32'd148483: dataIn1 = 32'd4393
; 
32'd148484: dataIn1 = 32'd485
; 
32'd148485: dataIn1 = 32'd2425
; 
32'd148486: dataIn1 = 32'd4375
; 
32'd148487: dataIn1 = 32'd4383
; 
32'd148488: dataIn1 = 32'd4385
; 
32'd148489: dataIn1 = 32'd4387
; 
32'd148490: dataIn1 = 32'd4391
; 
32'd148491: dataIn1 = 32'd2426
; 
32'd148492: dataIn1 = 32'd2427
; 
32'd148493: dataIn1 = 32'd4386
; 
32'd148494: dataIn1 = 32'd4387
; 
32'd148495: dataIn1 = 32'd4388
; 
32'd148496: dataIn1 = 32'd4389
; 
32'd148497: dataIn1 = 32'd4390
; 
32'd148498: dataIn1 = 32'd2425
; 
32'd148499: dataIn1 = 32'd2427
; 
32'd148500: dataIn1 = 32'd4385
; 
32'd148501: dataIn1 = 32'd4386
; 
32'd148502: dataIn1 = 32'd4387
; 
32'd148503: dataIn1 = 32'd4388
; 
32'd148504: dataIn1 = 32'd4391
; 
32'd148505: dataIn1 = 32'd2425
; 
32'd148506: dataIn1 = 32'd2426
; 
32'd148507: dataIn1 = 32'd4386
; 
32'd148508: dataIn1 = 32'd4387
; 
32'd148509: dataIn1 = 32'd4388
; 
32'd148510: dataIn1 = 32'd4392
; 
32'd148511: dataIn1 = 32'd4393
; 
32'd148512: dataIn1 = 32'd486
; 
32'd148513: dataIn1 = 32'd2427
; 
32'd148514: dataIn1 = 32'd4386
; 
32'd148515: dataIn1 = 32'd4389
; 
32'd148516: dataIn1 = 32'd4390
; 
32'd148517: dataIn1 = 32'd5391
; 
32'd148518: dataIn1 = 32'd486
; 
32'd148519: dataIn1 = 32'd2426
; 
32'd148520: dataIn1 = 32'd4386
; 
32'd148521: dataIn1 = 32'd4389
; 
32'd148522: dataIn1 = 32'd4390
; 
32'd148523: dataIn1 = 32'd4397
; 
32'd148524: dataIn1 = 32'd4407
; 
32'd148525: dataIn1 = 32'd485
; 
32'd148526: dataIn1 = 32'd2427
; 
32'd148527: dataIn1 = 32'd4385
; 
32'd148528: dataIn1 = 32'd4387
; 
32'd148529: dataIn1 = 32'd4391
; 
32'd148530: dataIn1 = 32'd5390
; 
32'd148531: dataIn1 = 32'd180
; 
32'd148532: dataIn1 = 32'd2426
; 
32'd148533: dataIn1 = 32'd3285
; 
32'd148534: dataIn1 = 32'd4388
; 
32'd148535: dataIn1 = 32'd4392
; 
32'd148536: dataIn1 = 32'd4393
; 
32'd148537: dataIn1 = 32'd4409
; 
32'd148538: dataIn1 = 32'd180
; 
32'd148539: dataIn1 = 32'd2425
; 
32'd148540: dataIn1 = 32'd3257
; 
32'd148541: dataIn1 = 32'd4384
; 
32'd148542: dataIn1 = 32'd4388
; 
32'd148543: dataIn1 = 32'd4392
; 
32'd148544: dataIn1 = 32'd4393
; 
32'd148545: dataIn1 = 32'd2429
; 
32'd148546: dataIn1 = 32'd2430
; 
32'd148547: dataIn1 = 32'd4394
; 
32'd148548: dataIn1 = 32'd4395
; 
32'd148549: dataIn1 = 32'd4396
; 
32'd148550: dataIn1 = 32'd4397
; 
32'd148551: dataIn1 = 32'd4398
; 
32'd148552: dataIn1 = 32'd2428
; 
32'd148553: dataIn1 = 32'd2430
; 
32'd148554: dataIn1 = 32'd4394
; 
32'd148555: dataIn1 = 32'd4395
; 
32'd148556: dataIn1 = 32'd4396
; 
32'd148557: dataIn1 = 32'd4399
; 
32'd148558: dataIn1 = 32'd4400
; 
32'd148559: dataIn1 = 32'd2428
; 
32'd148560: dataIn1 = 32'd2429
; 
32'd148561: dataIn1 = 32'd4394
; 
32'd148562: dataIn1 = 32'd4395
; 
32'd148563: dataIn1 = 32'd4396
; 
32'd148564: dataIn1 = 32'd4401
; 
32'd148565: dataIn1 = 32'd4402
; 
32'd148566: dataIn1 = 32'd486
; 
32'd148567: dataIn1 = 32'd2430
; 
32'd148568: dataIn1 = 32'd4390
; 
32'd148569: dataIn1 = 32'd4394
; 
32'd148570: dataIn1 = 32'd4397
; 
32'd148571: dataIn1 = 32'd4398
; 
32'd148572: dataIn1 = 32'd4407
; 
32'd148573: dataIn1 = 32'd486
; 
32'd148574: dataIn1 = 32'd2429
; 
32'd148575: dataIn1 = 32'd4394
; 
32'd148576: dataIn1 = 32'd4397
; 
32'd148577: dataIn1 = 32'd4398
; 
32'd148578: dataIn1 = 32'd5393
; 
32'd148579: dataIn1 = 32'd350
; 
32'd148580: dataIn1 = 32'd2430
; 
32'd148581: dataIn1 = 32'd3284
; 
32'd148582: dataIn1 = 32'd4395
; 
32'd148583: dataIn1 = 32'd4399
; 
32'd148584: dataIn1 = 32'd4400
; 
32'd148585: dataIn1 = 32'd4408
; 
32'd148586: dataIn1 = 32'd350
; 
32'd148587: dataIn1 = 32'd2428
; 
32'd148588: dataIn1 = 32'd3290
; 
32'd148589: dataIn1 = 32'd4395
; 
32'd148590: dataIn1 = 32'd4399
; 
32'd148591: dataIn1 = 32'd4400
; 
32'd148592: dataIn1 = 32'd4404
; 
32'd148593: dataIn1 = 32'd487
; 
32'd148594: dataIn1 = 32'd2429
; 
32'd148595: dataIn1 = 32'd4396
; 
32'd148596: dataIn1 = 32'd4401
; 
32'd148597: dataIn1 = 32'd4402
; 
32'd148598: dataIn1 = 32'd5392
; 
32'd148599: dataIn1 = 32'd487
; 
32'd148600: dataIn1 = 32'd2428
; 
32'd148601: dataIn1 = 32'd4396
; 
32'd148602: dataIn1 = 32'd4401
; 
32'd148603: dataIn1 = 32'd4402
; 
32'd148604: dataIn1 = 32'd4405
; 
32'd148605: dataIn1 = 32'd4406
; 
32'd148606: dataIn1 = 32'd2012
; 
32'd148607: dataIn1 = 32'd2431
; 
32'd148608: dataIn1 = 32'd3289
; 
32'd148609: dataIn1 = 32'd4403
; 
32'd148610: dataIn1 = 32'd4404
; 
32'd148611: dataIn1 = 32'd4405
; 
32'd148612: dataIn1 = 32'd4413
; 
32'd148613: dataIn1 = 32'd2012
; 
32'd148614: dataIn1 = 32'd2428
; 
32'd148615: dataIn1 = 32'd3290
; 
32'd148616: dataIn1 = 32'd4400
; 
32'd148617: dataIn1 = 32'd4403
; 
32'd148618: dataIn1 = 32'd4404
; 
32'd148619: dataIn1 = 32'd4405
; 
32'd148620: dataIn1 = 32'd2428
; 
32'd148621: dataIn1 = 32'd2431
; 
32'd148622: dataIn1 = 32'd4402
; 
32'd148623: dataIn1 = 32'd4403
; 
32'd148624: dataIn1 = 32'd4404
; 
32'd148625: dataIn1 = 32'd4405
; 
32'd148626: dataIn1 = 32'd4406
; 
32'd148627: dataIn1 = 32'd487
; 
32'd148628: dataIn1 = 32'd2431
; 
32'd148629: dataIn1 = 32'd4402
; 
32'd148630: dataIn1 = 32'd4405
; 
32'd148631: dataIn1 = 32'd4406
; 
32'd148632: dataIn1 = 32'd4411
; 
32'd148633: dataIn1 = 32'd4415
; 
32'd148634: dataIn1 = 32'd2426
; 
32'd148635: dataIn1 = 32'd2430
; 
32'd148636: dataIn1 = 32'd4390
; 
32'd148637: dataIn1 = 32'd4397
; 
32'd148638: dataIn1 = 32'd4407
; 
32'd148639: dataIn1 = 32'd4408
; 
32'd148640: dataIn1 = 32'd4409
; 
32'd148641: dataIn1 = 32'd2011
; 
32'd148642: dataIn1 = 32'd2430
; 
32'd148643: dataIn1 = 32'd3284
; 
32'd148644: dataIn1 = 32'd4399
; 
32'd148645: dataIn1 = 32'd4407
; 
32'd148646: dataIn1 = 32'd4408
; 
32'd148647: dataIn1 = 32'd4409
; 
32'd148648: dataIn1 = 32'd2011
; 
32'd148649: dataIn1 = 32'd2426
; 
32'd148650: dataIn1 = 32'd3285
; 
32'd148651: dataIn1 = 32'd4392
; 
32'd148652: dataIn1 = 32'd4407
; 
32'd148653: dataIn1 = 32'd4408
; 
32'd148654: dataIn1 = 32'd4409
; 
32'd148655: dataIn1 = 32'd2431
; 
32'd148656: dataIn1 = 32'd2433
; 
32'd148657: dataIn1 = 32'd4410
; 
32'd148658: dataIn1 = 32'd4411
; 
32'd148659: dataIn1 = 32'd4412
; 
32'd148660: dataIn1 = 32'd4413
; 
32'd148661: dataIn1 = 32'd4414
; 
32'd148662: dataIn1 = 32'd2431
; 
32'd148663: dataIn1 = 32'd2432
; 
32'd148664: dataIn1 = 32'd4406
; 
32'd148665: dataIn1 = 32'd4410
; 
32'd148666: dataIn1 = 32'd4411
; 
32'd148667: dataIn1 = 32'd4412
; 
32'd148668: dataIn1 = 32'd4415
; 
32'd148669: dataIn1 = 32'd2432
; 
32'd148670: dataIn1 = 32'd2433
; 
32'd148671: dataIn1 = 32'd4410
; 
32'd148672: dataIn1 = 32'd4411
; 
32'd148673: dataIn1 = 32'd4412
; 
32'd148674: dataIn1 = 32'd4416
; 
32'd148675: dataIn1 = 32'd4417
; 
32'd148676: dataIn1 = 32'd181
; 
32'd148677: dataIn1 = 32'd2431
; 
32'd148678: dataIn1 = 32'd3289
; 
32'd148679: dataIn1 = 32'd4403
; 
32'd148680: dataIn1 = 32'd4410
; 
32'd148681: dataIn1 = 32'd4413
; 
32'd148682: dataIn1 = 32'd4414
; 
32'd148683: dataIn1 = 32'd181
; 
32'd148684: dataIn1 = 32'd2433
; 
32'd148685: dataIn1 = 32'd3296
; 
32'd148686: dataIn1 = 32'd4410
; 
32'd148687: dataIn1 = 32'd4413
; 
32'd148688: dataIn1 = 32'd4414
; 
32'd148689: dataIn1 = 32'd4427
; 
32'd148690: dataIn1 = 32'd487
; 
32'd148691: dataIn1 = 32'd2432
; 
32'd148692: dataIn1 = 32'd4406
; 
32'd148693: dataIn1 = 32'd4411
; 
32'd148694: dataIn1 = 32'd4415
; 
32'd148695: dataIn1 = 32'd5395
; 
32'd148696: dataIn1 = 32'd488
; 
32'd148697: dataIn1 = 32'd2433
; 
32'd148698: dataIn1 = 32'd4412
; 
32'd148699: dataIn1 = 32'd4416
; 
32'd148700: dataIn1 = 32'd4417
; 
32'd148701: dataIn1 = 32'd4426
; 
32'd148702: dataIn1 = 32'd4429
; 
32'd148703: dataIn1 = 32'd488
; 
32'd148704: dataIn1 = 32'd2432
; 
32'd148705: dataIn1 = 32'd4412
; 
32'd148706: dataIn1 = 32'd4416
; 
32'd148707: dataIn1 = 32'd4417
; 
32'd148708: dataIn1 = 32'd5394
; 
32'd148709: dataIn1 = 32'd2435
; 
32'd148710: dataIn1 = 32'd2436
; 
32'd148711: dataIn1 = 32'd4418
; 
32'd148712: dataIn1 = 32'd4419
; 
32'd148713: dataIn1 = 32'd4420
; 
32'd148714: dataIn1 = 32'd4421
; 
32'd148715: dataIn1 = 32'd4422
; 
32'd148716: dataIn1 = 32'd2434
; 
32'd148717: dataIn1 = 32'd2436
; 
32'd148718: dataIn1 = 32'd4418
; 
32'd148719: dataIn1 = 32'd4419
; 
32'd148720: dataIn1 = 32'd4420
; 
32'd148721: dataIn1 = 32'd4423
; 
32'd148722: dataIn1 = 32'd4424
; 
32'd148723: dataIn1 = 32'd2434
; 
32'd148724: dataIn1 = 32'd2435
; 
32'd148725: dataIn1 = 32'd4418
; 
32'd148726: dataIn1 = 32'd4419
; 
32'd148727: dataIn1 = 32'd4420
; 
32'd148728: dataIn1 = 32'd4425
; 
32'd148729: dataIn1 = 32'd4426
; 
32'd148730: dataIn1 = 32'd489
; 
32'd148731: dataIn1 = 32'd2436
; 
32'd148732: dataIn1 = 32'd4418
; 
32'd148733: dataIn1 = 32'd4421
; 
32'd148734: dataIn1 = 32'd4422
; 
32'd148735: dataIn1 = 32'd4430
; 
32'd148736: dataIn1 = 32'd4433
; 
32'd148737: dataIn1 = 32'd489
; 
32'd148738: dataIn1 = 32'd2435
; 
32'd148739: dataIn1 = 32'd4418
; 
32'd148740: dataIn1 = 32'd4421
; 
32'd148741: dataIn1 = 32'd4422
; 
32'd148742: dataIn1 = 32'd5397
; 
32'd148743: dataIn1 = 32'd357
; 
32'd148744: dataIn1 = 32'd2436
; 
32'd148745: dataIn1 = 32'd3305
; 
32'd148746: dataIn1 = 32'd4419
; 
32'd148747: dataIn1 = 32'd4423
; 
32'd148748: dataIn1 = 32'd4424
; 
32'd148749: dataIn1 = 32'd4431
; 
32'd148750: dataIn1 = 32'd357
; 
32'd148751: dataIn1 = 32'd2434
; 
32'd148752: dataIn1 = 32'd3297
; 
32'd148753: dataIn1 = 32'd4419
; 
32'd148754: dataIn1 = 32'd4423
; 
32'd148755: dataIn1 = 32'd4424
; 
32'd148756: dataIn1 = 32'd4428
; 
32'd148757: dataIn1 = 32'd488
; 
32'd148758: dataIn1 = 32'd2435
; 
32'd148759: dataIn1 = 32'd4420
; 
32'd148760: dataIn1 = 32'd4425
; 
32'd148761: dataIn1 = 32'd4426
; 
32'd148762: dataIn1 = 32'd5396
; 
32'd148763: dataIn1 = 32'd488
; 
32'd148764: dataIn1 = 32'd2434
; 
32'd148765: dataIn1 = 32'd4416
; 
32'd148766: dataIn1 = 32'd4420
; 
32'd148767: dataIn1 = 32'd4425
; 
32'd148768: dataIn1 = 32'd4426
; 
32'd148769: dataIn1 = 32'd4429
; 
32'd148770: dataIn1 = 32'd2013
; 
32'd148771: dataIn1 = 32'd2433
; 
32'd148772: dataIn1 = 32'd3296
; 
32'd148773: dataIn1 = 32'd4414
; 
32'd148774: dataIn1 = 32'd4427
; 
32'd148775: dataIn1 = 32'd4428
; 
32'd148776: dataIn1 = 32'd4429
; 
32'd148777: dataIn1 = 32'd2013
; 
32'd148778: dataIn1 = 32'd2434
; 
32'd148779: dataIn1 = 32'd3297
; 
32'd148780: dataIn1 = 32'd4424
; 
32'd148781: dataIn1 = 32'd4427
; 
32'd148782: dataIn1 = 32'd4428
; 
32'd148783: dataIn1 = 32'd4429
; 
32'd148784: dataIn1 = 32'd2433
; 
32'd148785: dataIn1 = 32'd2434
; 
32'd148786: dataIn1 = 32'd4416
; 
32'd148787: dataIn1 = 32'd4426
; 
32'd148788: dataIn1 = 32'd4427
; 
32'd148789: dataIn1 = 32'd4428
; 
32'd148790: dataIn1 = 32'd4429
; 
32'd148791: dataIn1 = 32'd2436
; 
32'd148792: dataIn1 = 32'd2437
; 
32'd148793: dataIn1 = 32'd4421
; 
32'd148794: dataIn1 = 32'd4430
; 
32'd148795: dataIn1 = 32'd4431
; 
32'd148796: dataIn1 = 32'd4432
; 
32'd148797: dataIn1 = 32'd4433
; 
32'd148798: dataIn1 = 32'd2014
; 
32'd148799: dataIn1 = 32'd2436
; 
32'd148800: dataIn1 = 32'd3305
; 
32'd148801: dataIn1 = 32'd4423
; 
32'd148802: dataIn1 = 32'd4430
; 
32'd148803: dataIn1 = 32'd4431
; 
32'd148804: dataIn1 = 32'd4432
; 
32'd148805: dataIn1 = 32'd2014
; 
32'd148806: dataIn1 = 32'd2437
; 
32'd148807: dataIn1 = 32'd3306
; 
32'd148808: dataIn1 = 32'd4430
; 
32'd148809: dataIn1 = 32'd4431
; 
32'd148810: dataIn1 = 32'd4432
; 
32'd148811: dataIn1 = 32'd4440
; 
32'd148812: dataIn1 = 32'd489
; 
32'd148813: dataIn1 = 32'd2437
; 
32'd148814: dataIn1 = 32'd4421
; 
32'd148815: dataIn1 = 32'd4430
; 
32'd148816: dataIn1 = 32'd4433
; 
32'd148817: dataIn1 = 32'd4434
; 
32'd148818: dataIn1 = 32'd4437
; 
32'd148819: dataIn1 = 32'd2437
; 
32'd148820: dataIn1 = 32'd2439
; 
32'd148821: dataIn1 = 32'd4433
; 
32'd148822: dataIn1 = 32'd4434
; 
32'd148823: dataIn1 = 32'd4435
; 
32'd148824: dataIn1 = 32'd4436
; 
32'd148825: dataIn1 = 32'd4437
; 
32'd148826: dataIn1 = 32'd2438
; 
32'd148827: dataIn1 = 32'd2439
; 
32'd148828: dataIn1 = 32'd4434
; 
32'd148829: dataIn1 = 32'd4435
; 
32'd148830: dataIn1 = 32'd4436
; 
32'd148831: dataIn1 = 32'd4438
; 
32'd148832: dataIn1 = 32'd4439
; 
32'd148833: dataIn1 = 32'd2437
; 
32'd148834: dataIn1 = 32'd2438
; 
32'd148835: dataIn1 = 32'd4434
; 
32'd148836: dataIn1 = 32'd4435
; 
32'd148837: dataIn1 = 32'd4436
; 
32'd148838: dataIn1 = 32'd4440
; 
32'd148839: dataIn1 = 32'd4441
; 
32'd148840: dataIn1 = 32'd489
; 
32'd148841: dataIn1 = 32'd2439
; 
32'd148842: dataIn1 = 32'd4433
; 
32'd148843: dataIn1 = 32'd4434
; 
32'd148844: dataIn1 = 32'd4437
; 
32'd148845: dataIn1 = 32'd5399
; 
32'd148846: dataIn1 = 32'd490
; 
32'd148847: dataIn1 = 32'd2439
; 
32'd148848: dataIn1 = 32'd4435
; 
32'd148849: dataIn1 = 32'd4438
; 
32'd148850: dataIn1 = 32'd4439
; 
32'd148851: dataIn1 = 32'd5398
; 
32'd148852: dataIn1 = 32'd490
; 
32'd148853: dataIn1 = 32'd2438
; 
32'd148854: dataIn1 = 32'd4435
; 
32'd148855: dataIn1 = 32'd4438
; 
32'd148856: dataIn1 = 32'd4439
; 
32'd148857: dataIn1 = 32'd4448
; 
32'd148858: dataIn1 = 32'd4452
; 
32'd148859: dataIn1 = 32'd183
; 
32'd148860: dataIn1 = 32'd2437
; 
32'd148861: dataIn1 = 32'd3306
; 
32'd148862: dataIn1 = 32'd4432
; 
32'd148863: dataIn1 = 32'd4436
; 
32'd148864: dataIn1 = 32'd4440
; 
32'd148865: dataIn1 = 32'd4441
; 
32'd148866: dataIn1 = 32'd183
; 
32'd148867: dataIn1 = 32'd2438
; 
32'd148868: dataIn1 = 32'd3331
; 
32'd148869: dataIn1 = 32'd4436
; 
32'd148870: dataIn1 = 32'd4440
; 
32'd148871: dataIn1 = 32'd4441
; 
32'd148872: dataIn1 = 32'd4451
; 
32'd148873: dataIn1 = 32'd2441
; 
32'd148874: dataIn1 = 32'd2442
; 
32'd148875: dataIn1 = 32'd4442
; 
32'd148876: dataIn1 = 32'd4443
; 
32'd148877: dataIn1 = 32'd4444
; 
32'd148878: dataIn1 = 32'd4445
; 
32'd148879: dataIn1 = 32'd4446
; 
32'd148880: dataIn1 = 32'd2440
; 
32'd148881: dataIn1 = 32'd2442
; 
32'd148882: dataIn1 = 32'd4442
; 
32'd148883: dataIn1 = 32'd4443
; 
32'd148884: dataIn1 = 32'd4444
; 
32'd148885: dataIn1 = 32'd4447
; 
32'd148886: dataIn1 = 32'd4448
; 
32'd148887: dataIn1 = 32'd2440
; 
32'd148888: dataIn1 = 32'd2441
; 
32'd148889: dataIn1 = 32'd4442
; 
32'd148890: dataIn1 = 32'd4443
; 
32'd148891: dataIn1 = 32'd4444
; 
32'd148892: dataIn1 = 32'd4449
; 
32'd148893: dataIn1 = 32'd4450
; 
32'd148894: dataIn1 = 32'd491
; 
32'd148895: dataIn1 = 32'd2442
; 
32'd148896: dataIn1 = 32'd4442
; 
32'd148897: dataIn1 = 32'd4445
; 
32'd148898: dataIn1 = 32'd4446
; 
32'd148899: dataIn1 = 32'd5401
; 
32'd148900: dataIn1 = 32'd491
; 
32'd148901: dataIn1 = 32'd2441
; 
32'd148902: dataIn1 = 32'd4442
; 
32'd148903: dataIn1 = 32'd4445
; 
32'd148904: dataIn1 = 32'd4446
; 
32'd148905: dataIn1 = 32'd4454
; 
32'd148906: dataIn1 = 32'd4457
; 
32'd148907: dataIn1 = 32'd490
; 
32'd148908: dataIn1 = 32'd2442
; 
32'd148909: dataIn1 = 32'd4443
; 
32'd148910: dataIn1 = 32'd4447
; 
32'd148911: dataIn1 = 32'd4448
; 
32'd148912: dataIn1 = 32'd5400
; 
32'd148913: dataIn1 = 32'd490
; 
32'd148914: dataIn1 = 32'd2440
; 
32'd148915: dataIn1 = 32'd4439
; 
32'd148916: dataIn1 = 32'd4443
; 
32'd148917: dataIn1 = 32'd4447
; 
32'd148918: dataIn1 = 32'd4448
; 
32'd148919: dataIn1 = 32'd4452
; 
32'd148920: dataIn1 = 32'd365
; 
32'd148921: dataIn1 = 32'd2441
; 
32'd148922: dataIn1 = 32'd3327
; 
32'd148923: dataIn1 = 32'd4444
; 
32'd148924: dataIn1 = 32'd4449
; 
32'd148925: dataIn1 = 32'd4450
; 
32'd148926: dataIn1 = 32'd4456
; 
32'd148927: dataIn1 = 32'd365
; 
32'd148928: dataIn1 = 32'd2440
; 
32'd148929: dataIn1 = 32'd3334
; 
32'd148930: dataIn1 = 32'd4444
; 
32'd148931: dataIn1 = 32'd4449
; 
32'd148932: dataIn1 = 32'd4450
; 
32'd148933: dataIn1 = 32'd4453
; 
32'd148934: dataIn1 = 32'd2018
; 
32'd148935: dataIn1 = 32'd2438
; 
32'd148936: dataIn1 = 32'd3331
; 
32'd148937: dataIn1 = 32'd4441
; 
32'd148938: dataIn1 = 32'd4451
; 
32'd148939: dataIn1 = 32'd4452
; 
32'd148940: dataIn1 = 32'd4453
; 
32'd148941: dataIn1 = 32'd2438
; 
32'd148942: dataIn1 = 32'd2440
; 
32'd148943: dataIn1 = 32'd4439
; 
32'd148944: dataIn1 = 32'd4448
; 
32'd148945: dataIn1 = 32'd4451
; 
32'd148946: dataIn1 = 32'd4452
; 
32'd148947: dataIn1 = 32'd4453
; 
32'd148948: dataIn1 = 32'd2018
; 
32'd148949: dataIn1 = 32'd2440
; 
32'd148950: dataIn1 = 32'd3334
; 
32'd148951: dataIn1 = 32'd4450
; 
32'd148952: dataIn1 = 32'd4451
; 
32'd148953: dataIn1 = 32'd4452
; 
32'd148954: dataIn1 = 32'd4453
; 
32'd148955: dataIn1 = 32'd2441
; 
32'd148956: dataIn1 = 32'd2443
; 
32'd148957: dataIn1 = 32'd4446
; 
32'd148958: dataIn1 = 32'd4454
; 
32'd148959: dataIn1 = 32'd4455
; 
32'd148960: dataIn1 = 32'd4456
; 
32'd148961: dataIn1 = 32'd4457
; 
32'd148962: dataIn1 = 32'd2017
; 
32'd148963: dataIn1 = 32'd2443
; 
32'd148964: dataIn1 = 32'd3326
; 
32'd148965: dataIn1 = 32'd4454
; 
32'd148966: dataIn1 = 32'd4455
; 
32'd148967: dataIn1 = 32'd4456
; 
32'd148968: dataIn1 = 32'd4462
; 
32'd148969: dataIn1 = 32'd2017
; 
32'd148970: dataIn1 = 32'd2441
; 
32'd148971: dataIn1 = 32'd3327
; 
32'd148972: dataIn1 = 32'd4449
; 
32'd148973: dataIn1 = 32'd4454
; 
32'd148974: dataIn1 = 32'd4455
; 
32'd148975: dataIn1 = 32'd4456
; 
32'd148976: dataIn1 = 32'd491
; 
32'd148977: dataIn1 = 32'd2443
; 
32'd148978: dataIn1 = 32'd4446
; 
32'd148979: dataIn1 = 32'd4454
; 
32'd148980: dataIn1 = 32'd4457
; 
32'd148981: dataIn1 = 32'd4458
; 
32'd148982: dataIn1 = 32'd4461
; 
32'd148983: dataIn1 = 32'd2443
; 
32'd148984: dataIn1 = 32'd2445
; 
32'd148985: dataIn1 = 32'd4457
; 
32'd148986: dataIn1 = 32'd4458
; 
32'd148987: dataIn1 = 32'd4459
; 
32'd148988: dataIn1 = 32'd4460
; 
32'd148989: dataIn1 = 32'd4461
; 
32'd148990: dataIn1 = 32'd2443
; 
32'd148991: dataIn1 = 32'd2444
; 
32'd148992: dataIn1 = 32'd4458
; 
32'd148993: dataIn1 = 32'd4459
; 
32'd148994: dataIn1 = 32'd4460
; 
32'd148995: dataIn1 = 32'd4462
; 
32'd148996: dataIn1 = 32'd4463
; 
32'd148997: dataIn1 = 32'd2444
; 
32'd148998: dataIn1 = 32'd2445
; 
32'd148999: dataIn1 = 32'd4458
; 
32'd149000: dataIn1 = 32'd4459
; 
32'd149001: dataIn1 = 32'd4460
; 
32'd149002: dataIn1 = 32'd4464
; 
32'd149003: dataIn1 = 32'd4465
; 
32'd149004: dataIn1 = 32'd491
; 
32'd149005: dataIn1 = 32'd2445
; 
32'd149006: dataIn1 = 32'd4457
; 
32'd149007: dataIn1 = 32'd4458
; 
32'd149008: dataIn1 = 32'd4461
; 
32'd149009: dataIn1 = 32'd5403
; 
32'd149010: dataIn1 = 32'd185
; 
32'd149011: dataIn1 = 32'd2443
; 
32'd149012: dataIn1 = 32'd3326
; 
32'd149013: dataIn1 = 32'd4455
; 
32'd149014: dataIn1 = 32'd4459
; 
32'd149015: dataIn1 = 32'd4462
; 
32'd149016: dataIn1 = 32'd4463
; 
32'd149017: dataIn1 = 32'd185
; 
32'd149018: dataIn1 = 32'd2444
; 
32'd149019: dataIn1 = 32'd3318
; 
32'd149020: dataIn1 = 32'd4459
; 
32'd149021: dataIn1 = 32'd4462
; 
32'd149022: dataIn1 = 32'd4463
; 
32'd149023: dataIn1 = 32'd4476
; 
32'd149024: dataIn1 = 32'd492
; 
32'd149025: dataIn1 = 32'd2445
; 
32'd149026: dataIn1 = 32'd4460
; 
32'd149027: dataIn1 = 32'd4464
; 
32'd149028: dataIn1 = 32'd4465
; 
32'd149029: dataIn1 = 32'd5402
; 
32'd149030: dataIn1 = 32'd492
; 
32'd149031: dataIn1 = 32'd2444
; 
32'd149032: dataIn1 = 32'd4460
; 
32'd149033: dataIn1 = 32'd4464
; 
32'd149034: dataIn1 = 32'd4465
; 
32'd149035: dataIn1 = 32'd4473
; 
32'd149036: dataIn1 = 32'd4477
; 
32'd149037: dataIn1 = 32'd2447
; 
32'd149038: dataIn1 = 32'd2448
; 
32'd149039: dataIn1 = 32'd4466
; 
32'd149040: dataIn1 = 32'd4467
; 
32'd149041: dataIn1 = 32'd4468
; 
32'd149042: dataIn1 = 32'd4469
; 
32'd149043: dataIn1 = 32'd4470
; 
32'd149044: dataIn1 = 32'd2446
; 
32'd149045: dataIn1 = 32'd2448
; 
32'd149046: dataIn1 = 32'd4466
; 
32'd149047: dataIn1 = 32'd4467
; 
32'd149048: dataIn1 = 32'd4468
; 
32'd149049: dataIn1 = 32'd4471
; 
32'd149050: dataIn1 = 32'd4472
; 
32'd149051: dataIn1 = 32'd2446
; 
32'd149052: dataIn1 = 32'd2447
; 
32'd149053: dataIn1 = 32'd4466
; 
32'd149054: dataIn1 = 32'd4467
; 
32'd149055: dataIn1 = 32'd4468
; 
32'd149056: dataIn1 = 32'd4473
; 
32'd149057: dataIn1 = 32'd4474
; 
32'd149058: dataIn1 = 32'd359
; 
32'd149059: dataIn1 = 32'd2448
; 
32'd149060: dataIn1 = 32'd3310
; 
32'd149061: dataIn1 = 32'd4466
; 
32'd149062: dataIn1 = 32'd4469
; 
32'd149063: dataIn1 = 32'd4470
; 
32'd149064: dataIn1 = 32'd4478
; 
32'd149065: dataIn1 = 32'd359
; 
32'd149066: dataIn1 = 32'd2447
; 
32'd149067: dataIn1 = 32'd3317
; 
32'd149068: dataIn1 = 32'd4466
; 
32'd149069: dataIn1 = 32'd4469
; 
32'd149070: dataIn1 = 32'd4470
; 
32'd149071: dataIn1 = 32'd4475
; 
32'd149072: dataIn1 = 32'd493
; 
32'd149073: dataIn1 = 32'd2448
; 
32'd149074: dataIn1 = 32'd4467
; 
32'd149075: dataIn1 = 32'd4471
; 
32'd149076: dataIn1 = 32'd4472
; 
32'd149077: dataIn1 = 32'd4479
; 
32'd149078: dataIn1 = 32'd4481
; 
32'd149079: dataIn1 = 32'd493
; 
32'd149080: dataIn1 = 32'd2446
; 
32'd149081: dataIn1 = 32'd4467
; 
32'd149082: dataIn1 = 32'd4471
; 
32'd149083: dataIn1 = 32'd4472
; 
32'd149084: dataIn1 = 32'd5405
; 
32'd149085: dataIn1 = 32'd492
; 
32'd149086: dataIn1 = 32'd2447
; 
32'd149087: dataIn1 = 32'd4465
; 
32'd149088: dataIn1 = 32'd4468
; 
32'd149089: dataIn1 = 32'd4473
; 
32'd149090: dataIn1 = 32'd4474
; 
32'd149091: dataIn1 = 32'd4477
; 
32'd149092: dataIn1 = 32'd492
; 
32'd149093: dataIn1 = 32'd2446
; 
32'd149094: dataIn1 = 32'd4468
; 
32'd149095: dataIn1 = 32'd4473
; 
32'd149096: dataIn1 = 32'd4474
; 
32'd149097: dataIn1 = 32'd5404
; 
32'd149098: dataIn1 = 32'd2016
; 
32'd149099: dataIn1 = 32'd2447
; 
32'd149100: dataIn1 = 32'd3317
; 
32'd149101: dataIn1 = 32'd4470
; 
32'd149102: dataIn1 = 32'd4475
; 
32'd149103: dataIn1 = 32'd4476
; 
32'd149104: dataIn1 = 32'd4477
; 
32'd149105: dataIn1 = 32'd2016
; 
32'd149106: dataIn1 = 32'd2444
; 
32'd149107: dataIn1 = 32'd3318
; 
32'd149108: dataIn1 = 32'd4463
; 
32'd149109: dataIn1 = 32'd4475
; 
32'd149110: dataIn1 = 32'd4476
; 
32'd149111: dataIn1 = 32'd4477
; 
32'd149112: dataIn1 = 32'd2444
; 
32'd149113: dataIn1 = 32'd2447
; 
32'd149114: dataIn1 = 32'd4465
; 
32'd149115: dataIn1 = 32'd4473
; 
32'd149116: dataIn1 = 32'd4475
; 
32'd149117: dataIn1 = 32'd4476
; 
32'd149118: dataIn1 = 32'd4477
; 
32'd149119: dataIn1 = 32'd2015
; 
32'd149120: dataIn1 = 32'd2448
; 
32'd149121: dataIn1 = 32'd3310
; 
32'd149122: dataIn1 = 32'd4469
; 
32'd149123: dataIn1 = 32'd4478
; 
32'd149124: dataIn1 = 32'd4479
; 
32'd149125: dataIn1 = 32'd4480
; 
32'd149126: dataIn1 = 32'd2448
; 
32'd149127: dataIn1 = 32'd2449
; 
32'd149128: dataIn1 = 32'd4471
; 
32'd149129: dataIn1 = 32'd4478
; 
32'd149130: dataIn1 = 32'd4479
; 
32'd149131: dataIn1 = 32'd4480
; 
32'd149132: dataIn1 = 32'd4481
; 
32'd149133: dataIn1 = 32'd2015
; 
32'd149134: dataIn1 = 32'd2449
; 
32'd149135: dataIn1 = 32'd3313
; 
32'd149136: dataIn1 = 32'd4478
; 
32'd149137: dataIn1 = 32'd4479
; 
32'd149138: dataIn1 = 32'd4480
; 
32'd149139: dataIn1 = 32'd4489
; 
32'd149140: dataIn1 = 32'd493
; 
32'd149141: dataIn1 = 32'd2449
; 
32'd149142: dataIn1 = 32'd4471
; 
32'd149143: dataIn1 = 32'd4479
; 
32'd149144: dataIn1 = 32'd4481
; 
32'd149145: dataIn1 = 32'd4483
; 
32'd149146: dataIn1 = 32'd4487
; 
32'd149147: dataIn1 = 32'd2450
; 
32'd149148: dataIn1 = 32'd2451
; 
32'd149149: dataIn1 = 32'd4482
; 
32'd149150: dataIn1 = 32'd4483
; 
32'd149151: dataIn1 = 32'd4484
; 
32'd149152: dataIn1 = 32'd4485
; 
32'd149153: dataIn1 = 32'd4486
; 
32'd149154: dataIn1 = 32'd2449
; 
32'd149155: dataIn1 = 32'd2451
; 
32'd149156: dataIn1 = 32'd4481
; 
32'd149157: dataIn1 = 32'd4482
; 
32'd149158: dataIn1 = 32'd4483
; 
32'd149159: dataIn1 = 32'd4484
; 
32'd149160: dataIn1 = 32'd4487
; 
32'd149161: dataIn1 = 32'd2449
; 
32'd149162: dataIn1 = 32'd2450
; 
32'd149163: dataIn1 = 32'd4482
; 
32'd149164: dataIn1 = 32'd4483
; 
32'd149165: dataIn1 = 32'd4484
; 
32'd149166: dataIn1 = 32'd4488
; 
32'd149167: dataIn1 = 32'd4489
; 
32'd149168: dataIn1 = 32'd494
; 
32'd149169: dataIn1 = 32'd2451
; 
32'd149170: dataIn1 = 32'd4482
; 
32'd149171: dataIn1 = 32'd4485
; 
32'd149172: dataIn1 = 32'd4486
; 
32'd149173: dataIn1 = 32'd5407
; 
32'd149174: dataIn1 = 32'd494
; 
32'd149175: dataIn1 = 32'd2450
; 
32'd149176: dataIn1 = 32'd4482
; 
32'd149177: dataIn1 = 32'd4485
; 
32'd149178: dataIn1 = 32'd4486
; 
32'd149179: dataIn1 = 32'd4493
; 
32'd149180: dataIn1 = 32'd4503
; 
32'd149181: dataIn1 = 32'd493
; 
32'd149182: dataIn1 = 32'd2451
; 
32'd149183: dataIn1 = 32'd4481
; 
32'd149184: dataIn1 = 32'd4483
; 
32'd149185: dataIn1 = 32'd4487
; 
32'd149186: dataIn1 = 32'd5406
; 
32'd149187: dataIn1 = 32'd186
; 
32'd149188: dataIn1 = 32'd2450
; 
32'd149189: dataIn1 = 32'd3341
; 
32'd149190: dataIn1 = 32'd4484
; 
32'd149191: dataIn1 = 32'd4488
; 
32'd149192: dataIn1 = 32'd4489
; 
32'd149193: dataIn1 = 32'd4505
; 
32'd149194: dataIn1 = 32'd186
; 
32'd149195: dataIn1 = 32'd2449
; 
32'd149196: dataIn1 = 32'd3313
; 
32'd149197: dataIn1 = 32'd4480
; 
32'd149198: dataIn1 = 32'd4484
; 
32'd149199: dataIn1 = 32'd4488
; 
32'd149200: dataIn1 = 32'd4489
; 
32'd149201: dataIn1 = 32'd2453
; 
32'd149202: dataIn1 = 32'd2454
; 
32'd149203: dataIn1 = 32'd4490
; 
32'd149204: dataIn1 = 32'd4491
; 
32'd149205: dataIn1 = 32'd4492
; 
32'd149206: dataIn1 = 32'd4493
; 
32'd149207: dataIn1 = 32'd4494
; 
32'd149208: dataIn1 = 32'd2452
; 
32'd149209: dataIn1 = 32'd2454
; 
32'd149210: dataIn1 = 32'd4490
; 
32'd149211: dataIn1 = 32'd4491
; 
32'd149212: dataIn1 = 32'd4492
; 
32'd149213: dataIn1 = 32'd4495
; 
32'd149214: dataIn1 = 32'd4496
; 
32'd149215: dataIn1 = 32'd2452
; 
32'd149216: dataIn1 = 32'd2453
; 
32'd149217: dataIn1 = 32'd4490
; 
32'd149218: dataIn1 = 32'd4491
; 
32'd149219: dataIn1 = 32'd4492
; 
32'd149220: dataIn1 = 32'd4497
; 
32'd149221: dataIn1 = 32'd4498
; 
32'd149222: dataIn1 = 32'd494
; 
32'd149223: dataIn1 = 32'd2454
; 
32'd149224: dataIn1 = 32'd4486
; 
32'd149225: dataIn1 = 32'd4490
; 
32'd149226: dataIn1 = 32'd4493
; 
32'd149227: dataIn1 = 32'd4494
; 
32'd149228: dataIn1 = 32'd4503
; 
32'd149229: dataIn1 = 32'd494
; 
32'd149230: dataIn1 = 32'd2453
; 
32'd149231: dataIn1 = 32'd4490
; 
32'd149232: dataIn1 = 32'd4493
; 
32'd149233: dataIn1 = 32'd4494
; 
32'd149234: dataIn1 = 32'd5409
; 
32'd149235: dataIn1 = 32'd366
; 
32'd149236: dataIn1 = 32'd2454
; 
32'd149237: dataIn1 = 32'd3340
; 
32'd149238: dataIn1 = 32'd4491
; 
32'd149239: dataIn1 = 32'd4495
; 
32'd149240: dataIn1 = 32'd4496
; 
32'd149241: dataIn1 = 32'd4504
; 
32'd149242: dataIn1 = 32'd366
; 
32'd149243: dataIn1 = 32'd2452
; 
32'd149244: dataIn1 = 32'd3346
; 
32'd149245: dataIn1 = 32'd4491
; 
32'd149246: dataIn1 = 32'd4495
; 
32'd149247: dataIn1 = 32'd4496
; 
32'd149248: dataIn1 = 32'd4500
; 
32'd149249: dataIn1 = 32'd495
; 
32'd149250: dataIn1 = 32'd2453
; 
32'd149251: dataIn1 = 32'd4492
; 
32'd149252: dataIn1 = 32'd4497
; 
32'd149253: dataIn1 = 32'd4498
; 
32'd149254: dataIn1 = 32'd5408
; 
32'd149255: dataIn1 = 32'd495
; 
32'd149256: dataIn1 = 32'd2452
; 
32'd149257: dataIn1 = 32'd4492
; 
32'd149258: dataIn1 = 32'd4497
; 
32'd149259: dataIn1 = 32'd4498
; 
32'd149260: dataIn1 = 32'd4501
; 
32'd149261: dataIn1 = 32'd4502
; 
32'd149262: dataIn1 = 32'd2020
; 
32'd149263: dataIn1 = 32'd2455
; 
32'd149264: dataIn1 = 32'd3345
; 
32'd149265: dataIn1 = 32'd4499
; 
32'd149266: dataIn1 = 32'd4500
; 
32'd149267: dataIn1 = 32'd4501
; 
32'd149268: dataIn1 = 32'd4509
; 
32'd149269: dataIn1 = 32'd2020
; 
32'd149270: dataIn1 = 32'd2452
; 
32'd149271: dataIn1 = 32'd3346
; 
32'd149272: dataIn1 = 32'd4496
; 
32'd149273: dataIn1 = 32'd4499
; 
32'd149274: dataIn1 = 32'd4500
; 
32'd149275: dataIn1 = 32'd4501
; 
32'd149276: dataIn1 = 32'd2452
; 
32'd149277: dataIn1 = 32'd2455
; 
32'd149278: dataIn1 = 32'd4498
; 
32'd149279: dataIn1 = 32'd4499
; 
32'd149280: dataIn1 = 32'd4500
; 
32'd149281: dataIn1 = 32'd4501
; 
32'd149282: dataIn1 = 32'd4502
; 
32'd149283: dataIn1 = 32'd495
; 
32'd149284: dataIn1 = 32'd2455
; 
32'd149285: dataIn1 = 32'd4498
; 
32'd149286: dataIn1 = 32'd4501
; 
32'd149287: dataIn1 = 32'd4502
; 
32'd149288: dataIn1 = 32'd4507
; 
32'd149289: dataIn1 = 32'd4511
; 
32'd149290: dataIn1 = 32'd2450
; 
32'd149291: dataIn1 = 32'd2454
; 
32'd149292: dataIn1 = 32'd4486
; 
32'd149293: dataIn1 = 32'd4493
; 
32'd149294: dataIn1 = 32'd4503
; 
32'd149295: dataIn1 = 32'd4504
; 
32'd149296: dataIn1 = 32'd4505
; 
32'd149297: dataIn1 = 32'd2019
; 
32'd149298: dataIn1 = 32'd2454
; 
32'd149299: dataIn1 = 32'd3340
; 
32'd149300: dataIn1 = 32'd4495
; 
32'd149301: dataIn1 = 32'd4503
; 
32'd149302: dataIn1 = 32'd4504
; 
32'd149303: dataIn1 = 32'd4505
; 
32'd149304: dataIn1 = 32'd2019
; 
32'd149305: dataIn1 = 32'd2450
; 
32'd149306: dataIn1 = 32'd3341
; 
32'd149307: dataIn1 = 32'd4488
; 
32'd149308: dataIn1 = 32'd4503
; 
32'd149309: dataIn1 = 32'd4504
; 
32'd149310: dataIn1 = 32'd4505
; 
32'd149311: dataIn1 = 32'd2455
; 
32'd149312: dataIn1 = 32'd2457
; 
32'd149313: dataIn1 = 32'd4506
; 
32'd149314: dataIn1 = 32'd4507
; 
32'd149315: dataIn1 = 32'd4508
; 
32'd149316: dataIn1 = 32'd4509
; 
32'd149317: dataIn1 = 32'd4510
; 
32'd149318: dataIn1 = 32'd2455
; 
32'd149319: dataIn1 = 32'd2456
; 
32'd149320: dataIn1 = 32'd4502
; 
32'd149321: dataIn1 = 32'd4506
; 
32'd149322: dataIn1 = 32'd4507
; 
32'd149323: dataIn1 = 32'd4508
; 
32'd149324: dataIn1 = 32'd4511
; 
32'd149325: dataIn1 = 32'd2456
; 
32'd149326: dataIn1 = 32'd2457
; 
32'd149327: dataIn1 = 32'd4506
; 
32'd149328: dataIn1 = 32'd4507
; 
32'd149329: dataIn1 = 32'd4508
; 
32'd149330: dataIn1 = 32'd4512
; 
32'd149331: dataIn1 = 32'd4513
; 
32'd149332: dataIn1 = 32'd187
; 
32'd149333: dataIn1 = 32'd2455
; 
32'd149334: dataIn1 = 32'd3345
; 
32'd149335: dataIn1 = 32'd4499
; 
32'd149336: dataIn1 = 32'd4506
; 
32'd149337: dataIn1 = 32'd4509
; 
32'd149338: dataIn1 = 32'd4510
; 
32'd149339: dataIn1 = 32'd187
; 
32'd149340: dataIn1 = 32'd2457
; 
32'd149341: dataIn1 = 32'd3352
; 
32'd149342: dataIn1 = 32'd4506
; 
32'd149343: dataIn1 = 32'd4509
; 
32'd149344: dataIn1 = 32'd4510
; 
32'd149345: dataIn1 = 32'd4523
; 
32'd149346: dataIn1 = 32'd495
; 
32'd149347: dataIn1 = 32'd2456
; 
32'd149348: dataIn1 = 32'd4502
; 
32'd149349: dataIn1 = 32'd4507
; 
32'd149350: dataIn1 = 32'd4511
; 
32'd149351: dataIn1 = 32'd5411
; 
32'd149352: dataIn1 = 32'd496
; 
32'd149353: dataIn1 = 32'd2457
; 
32'd149354: dataIn1 = 32'd4508
; 
32'd149355: dataIn1 = 32'd4512
; 
32'd149356: dataIn1 = 32'd4513
; 
32'd149357: dataIn1 = 32'd4522
; 
32'd149358: dataIn1 = 32'd4525
; 
32'd149359: dataIn1 = 32'd496
; 
32'd149360: dataIn1 = 32'd2456
; 
32'd149361: dataIn1 = 32'd4508
; 
32'd149362: dataIn1 = 32'd4512
; 
32'd149363: dataIn1 = 32'd4513
; 
32'd149364: dataIn1 = 32'd5410
; 
32'd149365: dataIn1 = 32'd2459
; 
32'd149366: dataIn1 = 32'd2460
; 
32'd149367: dataIn1 = 32'd4514
; 
32'd149368: dataIn1 = 32'd4515
; 
32'd149369: dataIn1 = 32'd4516
; 
32'd149370: dataIn1 = 32'd4517
; 
32'd149371: dataIn1 = 32'd4518
; 
32'd149372: dataIn1 = 32'd2458
; 
32'd149373: dataIn1 = 32'd2460
; 
32'd149374: dataIn1 = 32'd4514
; 
32'd149375: dataIn1 = 32'd4515
; 
32'd149376: dataIn1 = 32'd4516
; 
32'd149377: dataIn1 = 32'd4519
; 
32'd149378: dataIn1 = 32'd4520
; 
32'd149379: dataIn1 = 32'd2458
; 
32'd149380: dataIn1 = 32'd2459
; 
32'd149381: dataIn1 = 32'd4514
; 
32'd149382: dataIn1 = 32'd4515
; 
32'd149383: dataIn1 = 32'd4516
; 
32'd149384: dataIn1 = 32'd4521
; 
32'd149385: dataIn1 = 32'd4522
; 
32'd149386: dataIn1 = 32'd497
; 
32'd149387: dataIn1 = 32'd2460
; 
32'd149388: dataIn1 = 32'd4514
; 
32'd149389: dataIn1 = 32'd4517
; 
32'd149390: dataIn1 = 32'd4518
; 
32'd149391: dataIn1 = 32'd4526
; 
32'd149392: dataIn1 = 32'd4529
; 
32'd149393: dataIn1 = 32'd497
; 
32'd149394: dataIn1 = 32'd2459
; 
32'd149395: dataIn1 = 32'd4514
; 
32'd149396: dataIn1 = 32'd4517
; 
32'd149397: dataIn1 = 32'd4518
; 
32'd149398: dataIn1 = 32'd5413
; 
32'd149399: dataIn1 = 32'd373
; 
32'd149400: dataIn1 = 32'd2460
; 
32'd149401: dataIn1 = 32'd3361
; 
32'd149402: dataIn1 = 32'd4515
; 
32'd149403: dataIn1 = 32'd4519
; 
32'd149404: dataIn1 = 32'd4520
; 
32'd149405: dataIn1 = 32'd4527
; 
32'd149406: dataIn1 = 32'd373
; 
32'd149407: dataIn1 = 32'd2458
; 
32'd149408: dataIn1 = 32'd3353
; 
32'd149409: dataIn1 = 32'd4515
; 
32'd149410: dataIn1 = 32'd4519
; 
32'd149411: dataIn1 = 32'd4520
; 
32'd149412: dataIn1 = 32'd4524
; 
32'd149413: dataIn1 = 32'd496
; 
32'd149414: dataIn1 = 32'd2459
; 
32'd149415: dataIn1 = 32'd4516
; 
32'd149416: dataIn1 = 32'd4521
; 
32'd149417: dataIn1 = 32'd4522
; 
32'd149418: dataIn1 = 32'd5412
; 
32'd149419: dataIn1 = 32'd496
; 
32'd149420: dataIn1 = 32'd2458
; 
32'd149421: dataIn1 = 32'd4512
; 
32'd149422: dataIn1 = 32'd4516
; 
32'd149423: dataIn1 = 32'd4521
; 
32'd149424: dataIn1 = 32'd4522
; 
32'd149425: dataIn1 = 32'd4525
; 
32'd149426: dataIn1 = 32'd2021
; 
32'd149427: dataIn1 = 32'd2457
; 
32'd149428: dataIn1 = 32'd3352
; 
32'd149429: dataIn1 = 32'd4510
; 
32'd149430: dataIn1 = 32'd4523
; 
32'd149431: dataIn1 = 32'd4524
; 
32'd149432: dataIn1 = 32'd4525
; 
32'd149433: dataIn1 = 32'd2021
; 
32'd149434: dataIn1 = 32'd2458
; 
32'd149435: dataIn1 = 32'd3353
; 
32'd149436: dataIn1 = 32'd4520
; 
32'd149437: dataIn1 = 32'd4523
; 
32'd149438: dataIn1 = 32'd4524
; 
32'd149439: dataIn1 = 32'd4525
; 
32'd149440: dataIn1 = 32'd2457
; 
32'd149441: dataIn1 = 32'd2458
; 
32'd149442: dataIn1 = 32'd4512
; 
32'd149443: dataIn1 = 32'd4522
; 
32'd149444: dataIn1 = 32'd4523
; 
32'd149445: dataIn1 = 32'd4524
; 
32'd149446: dataIn1 = 32'd4525
; 
32'd149447: dataIn1 = 32'd2460
; 
32'd149448: dataIn1 = 32'd2461
; 
32'd149449: dataIn1 = 32'd4517
; 
32'd149450: dataIn1 = 32'd4526
; 
32'd149451: dataIn1 = 32'd4527
; 
32'd149452: dataIn1 = 32'd4528
; 
32'd149453: dataIn1 = 32'd4529
; 
32'd149454: dataIn1 = 32'd2022
; 
32'd149455: dataIn1 = 32'd2460
; 
32'd149456: dataIn1 = 32'd3361
; 
32'd149457: dataIn1 = 32'd4519
; 
32'd149458: dataIn1 = 32'd4526
; 
32'd149459: dataIn1 = 32'd4527
; 
32'd149460: dataIn1 = 32'd4528
; 
32'd149461: dataIn1 = 32'd2022
; 
32'd149462: dataIn1 = 32'd2461
; 
32'd149463: dataIn1 = 32'd3362
; 
32'd149464: dataIn1 = 32'd4526
; 
32'd149465: dataIn1 = 32'd4527
; 
32'd149466: dataIn1 = 32'd4528
; 
32'd149467: dataIn1 = 32'd4536
; 
32'd149468: dataIn1 = 32'd497
; 
32'd149469: dataIn1 = 32'd2461
; 
32'd149470: dataIn1 = 32'd4517
; 
32'd149471: dataIn1 = 32'd4526
; 
32'd149472: dataIn1 = 32'd4529
; 
32'd149473: dataIn1 = 32'd4530
; 
32'd149474: dataIn1 = 32'd4533
; 
32'd149475: dataIn1 = 32'd2461
; 
32'd149476: dataIn1 = 32'd2463
; 
32'd149477: dataIn1 = 32'd4529
; 
32'd149478: dataIn1 = 32'd4530
; 
32'd149479: dataIn1 = 32'd4531
; 
32'd149480: dataIn1 = 32'd4532
; 
32'd149481: dataIn1 = 32'd4533
; 
32'd149482: dataIn1 = 32'd2462
; 
32'd149483: dataIn1 = 32'd2463
; 
32'd149484: dataIn1 = 32'd4530
; 
32'd149485: dataIn1 = 32'd4531
; 
32'd149486: dataIn1 = 32'd4532
; 
32'd149487: dataIn1 = 32'd4534
; 
32'd149488: dataIn1 = 32'd4535
; 
32'd149489: dataIn1 = 32'd2461
; 
32'd149490: dataIn1 = 32'd2462
; 
32'd149491: dataIn1 = 32'd4530
; 
32'd149492: dataIn1 = 32'd4531
; 
32'd149493: dataIn1 = 32'd4532
; 
32'd149494: dataIn1 = 32'd4536
; 
32'd149495: dataIn1 = 32'd4537
; 
32'd149496: dataIn1 = 32'd497
; 
32'd149497: dataIn1 = 32'd2463
; 
32'd149498: dataIn1 = 32'd4529
; 
32'd149499: dataIn1 = 32'd4530
; 
32'd149500: dataIn1 = 32'd4533
; 
32'd149501: dataIn1 = 32'd5415
; 
32'd149502: dataIn1 = 32'd498
; 
32'd149503: dataIn1 = 32'd2463
; 
32'd149504: dataIn1 = 32'd4531
; 
32'd149505: dataIn1 = 32'd4534
; 
32'd149506: dataIn1 = 32'd4535
; 
32'd149507: dataIn1 = 32'd5414
; 
32'd149508: dataIn1 = 32'd498
; 
32'd149509: dataIn1 = 32'd2462
; 
32'd149510: dataIn1 = 32'd4531
; 
32'd149511: dataIn1 = 32'd4534
; 
32'd149512: dataIn1 = 32'd4535
; 
32'd149513: dataIn1 = 32'd4544
; 
32'd149514: dataIn1 = 32'd4548
; 
32'd149515: dataIn1 = 32'd189
; 
32'd149516: dataIn1 = 32'd2461
; 
32'd149517: dataIn1 = 32'd3362
; 
32'd149518: dataIn1 = 32'd4528
; 
32'd149519: dataIn1 = 32'd4532
; 
32'd149520: dataIn1 = 32'd4536
; 
32'd149521: dataIn1 = 32'd4537
; 
32'd149522: dataIn1 = 32'd189
; 
32'd149523: dataIn1 = 32'd2462
; 
32'd149524: dataIn1 = 32'd3387
; 
32'd149525: dataIn1 = 32'd4532
; 
32'd149526: dataIn1 = 32'd4536
; 
32'd149527: dataIn1 = 32'd4537
; 
32'd149528: dataIn1 = 32'd4547
; 
32'd149529: dataIn1 = 32'd2465
; 
32'd149530: dataIn1 = 32'd2466
; 
32'd149531: dataIn1 = 32'd4538
; 
32'd149532: dataIn1 = 32'd4539
; 
32'd149533: dataIn1 = 32'd4540
; 
32'd149534: dataIn1 = 32'd4541
; 
32'd149535: dataIn1 = 32'd4542
; 
32'd149536: dataIn1 = 32'd2464
; 
32'd149537: dataIn1 = 32'd2466
; 
32'd149538: dataIn1 = 32'd4538
; 
32'd149539: dataIn1 = 32'd4539
; 
32'd149540: dataIn1 = 32'd4540
; 
32'd149541: dataIn1 = 32'd4543
; 
32'd149542: dataIn1 = 32'd4544
; 
32'd149543: dataIn1 = 32'd2464
; 
32'd149544: dataIn1 = 32'd2465
; 
32'd149545: dataIn1 = 32'd4538
; 
32'd149546: dataIn1 = 32'd4539
; 
32'd149547: dataIn1 = 32'd4540
; 
32'd149548: dataIn1 = 32'd4545
; 
32'd149549: dataIn1 = 32'd4546
; 
32'd149550: dataIn1 = 32'd499
; 
32'd149551: dataIn1 = 32'd2466
; 
32'd149552: dataIn1 = 32'd4538
; 
32'd149553: dataIn1 = 32'd4541
; 
32'd149554: dataIn1 = 32'd4542
; 
32'd149555: dataIn1 = 32'd5416
; 
32'd149556: dataIn1 = 32'd5417
; 
32'd149557: dataIn1 = 32'd499
; 
32'd149558: dataIn1 = 32'd2465
; 
32'd149559: dataIn1 = 32'd4538
; 
32'd149560: dataIn1 = 32'd4541
; 
32'd149561: dataIn1 = 32'd4542
; 
32'd149562: dataIn1 = 32'd4550
; 
32'd149563: dataIn1 = 32'd4553
; 
32'd149564: dataIn1 = 32'd498
; 
32'd149565: dataIn1 = 32'd2466
; 
32'd149566: dataIn1 = 32'd4539
; 
32'd149567: dataIn1 = 32'd4543
; 
32'd149568: dataIn1 = 32'd4544
; 
32'd149569: dataIn1 = 32'd5416
; 
32'd149570: dataIn1 = 32'd498
; 
32'd149571: dataIn1 = 32'd2464
; 
32'd149572: dataIn1 = 32'd4535
; 
32'd149573: dataIn1 = 32'd4539
; 
32'd149574: dataIn1 = 32'd4543
; 
32'd149575: dataIn1 = 32'd4544
; 
32'd149576: dataIn1 = 32'd4548
; 
32'd149577: dataIn1 = 32'd381
; 
32'd149578: dataIn1 = 32'd2465
; 
32'd149579: dataIn1 = 32'd3383
; 
32'd149580: dataIn1 = 32'd4540
; 
32'd149581: dataIn1 = 32'd4545
; 
32'd149582: dataIn1 = 32'd4546
; 
32'd149583: dataIn1 = 32'd4552
; 
32'd149584: dataIn1 = 32'd381
; 
32'd149585: dataIn1 = 32'd2464
; 
32'd149586: dataIn1 = 32'd3390
; 
32'd149587: dataIn1 = 32'd4540
; 
32'd149588: dataIn1 = 32'd4545
; 
32'd149589: dataIn1 = 32'd4546
; 
32'd149590: dataIn1 = 32'd4549
; 
32'd149591: dataIn1 = 32'd2026
; 
32'd149592: dataIn1 = 32'd2462
; 
32'd149593: dataIn1 = 32'd3387
; 
32'd149594: dataIn1 = 32'd4537
; 
32'd149595: dataIn1 = 32'd4547
; 
32'd149596: dataIn1 = 32'd4548
; 
32'd149597: dataIn1 = 32'd4549
; 
32'd149598: dataIn1 = 32'd2462
; 
32'd149599: dataIn1 = 32'd2464
; 
32'd149600: dataIn1 = 32'd4535
; 
32'd149601: dataIn1 = 32'd4544
; 
32'd149602: dataIn1 = 32'd4547
; 
32'd149603: dataIn1 = 32'd4548
; 
32'd149604: dataIn1 = 32'd4549
; 
32'd149605: dataIn1 = 32'd2026
; 
32'd149606: dataIn1 = 32'd2464
; 
32'd149607: dataIn1 = 32'd3390
; 
32'd149608: dataIn1 = 32'd4546
; 
32'd149609: dataIn1 = 32'd4547
; 
32'd149610: dataIn1 = 32'd4548
; 
32'd149611: dataIn1 = 32'd4549
; 
32'd149612: dataIn1 = 32'd2465
; 
32'd149613: dataIn1 = 32'd2467
; 
32'd149614: dataIn1 = 32'd4542
; 
32'd149615: dataIn1 = 32'd4550
; 
32'd149616: dataIn1 = 32'd4551
; 
32'd149617: dataIn1 = 32'd4552
; 
32'd149618: dataIn1 = 32'd4553
; 
32'd149619: dataIn1 = 32'd2025
; 
32'd149620: dataIn1 = 32'd2467
; 
32'd149621: dataIn1 = 32'd3382
; 
32'd149622: dataIn1 = 32'd4550
; 
32'd149623: dataIn1 = 32'd4551
; 
32'd149624: dataIn1 = 32'd4552
; 
32'd149625: dataIn1 = 32'd4558
; 
32'd149626: dataIn1 = 32'd2025
; 
32'd149627: dataIn1 = 32'd2465
; 
32'd149628: dataIn1 = 32'd3383
; 
32'd149629: dataIn1 = 32'd4545
; 
32'd149630: dataIn1 = 32'd4550
; 
32'd149631: dataIn1 = 32'd4551
; 
32'd149632: dataIn1 = 32'd4552
; 
32'd149633: dataIn1 = 32'd499
; 
32'd149634: dataIn1 = 32'd2467
; 
32'd149635: dataIn1 = 32'd4542
; 
32'd149636: dataIn1 = 32'd4550
; 
32'd149637: dataIn1 = 32'd4553
; 
32'd149638: dataIn1 = 32'd4554
; 
32'd149639: dataIn1 = 32'd4557
; 
32'd149640: dataIn1 = 32'd2467
; 
32'd149641: dataIn1 = 32'd2469
; 
32'd149642: dataIn1 = 32'd4553
; 
32'd149643: dataIn1 = 32'd4554
; 
32'd149644: dataIn1 = 32'd4555
; 
32'd149645: dataIn1 = 32'd4556
; 
32'd149646: dataIn1 = 32'd4557
; 
32'd149647: dataIn1 = 32'd2467
; 
32'd149648: dataIn1 = 32'd2468
; 
32'd149649: dataIn1 = 32'd4554
; 
32'd149650: dataIn1 = 32'd4555
; 
32'd149651: dataIn1 = 32'd4556
; 
32'd149652: dataIn1 = 32'd4558
; 
32'd149653: dataIn1 = 32'd4559
; 
32'd149654: dataIn1 = 32'd2468
; 
32'd149655: dataIn1 = 32'd2469
; 
32'd149656: dataIn1 = 32'd4554
; 
32'd149657: dataIn1 = 32'd4555
; 
32'd149658: dataIn1 = 32'd4556
; 
32'd149659: dataIn1 = 32'd4560
; 
32'd149660: dataIn1 = 32'd4561
; 
32'd149661: dataIn1 = 32'd499
; 
32'd149662: dataIn1 = 32'd2469
; 
32'd149663: dataIn1 = 32'd4553
; 
32'd149664: dataIn1 = 32'd4554
; 
32'd149665: dataIn1 = 32'd4557
; 
32'd149666: dataIn1 = 32'd5417
; 
32'd149667: dataIn1 = 32'd5419
; 
32'd149668: dataIn1 = 32'd191
; 
32'd149669: dataIn1 = 32'd2467
; 
32'd149670: dataIn1 = 32'd3382
; 
32'd149671: dataIn1 = 32'd4551
; 
32'd149672: dataIn1 = 32'd4555
; 
32'd149673: dataIn1 = 32'd4558
; 
32'd149674: dataIn1 = 32'd4559
; 
32'd149675: dataIn1 = 32'd191
; 
32'd149676: dataIn1 = 32'd2468
; 
32'd149677: dataIn1 = 32'd3374
; 
32'd149678: dataIn1 = 32'd4555
; 
32'd149679: dataIn1 = 32'd4558
; 
32'd149680: dataIn1 = 32'd4559
; 
32'd149681: dataIn1 = 32'd4572
; 
32'd149682: dataIn1 = 32'd500
; 
32'd149683: dataIn1 = 32'd2469
; 
32'd149684: dataIn1 = 32'd4556
; 
32'd149685: dataIn1 = 32'd4560
; 
32'd149686: dataIn1 = 32'd4561
; 
32'd149687: dataIn1 = 32'd5418
; 
32'd149688: dataIn1 = 32'd5419
; 
32'd149689: dataIn1 = 32'd500
; 
32'd149690: dataIn1 = 32'd2468
; 
32'd149691: dataIn1 = 32'd4556
; 
32'd149692: dataIn1 = 32'd4560
; 
32'd149693: dataIn1 = 32'd4561
; 
32'd149694: dataIn1 = 32'd4569
; 
32'd149695: dataIn1 = 32'd4573
; 
32'd149696: dataIn1 = 32'd2471
; 
32'd149697: dataIn1 = 32'd2472
; 
32'd149698: dataIn1 = 32'd4562
; 
32'd149699: dataIn1 = 32'd4563
; 
32'd149700: dataIn1 = 32'd4564
; 
32'd149701: dataIn1 = 32'd4565
; 
32'd149702: dataIn1 = 32'd4566
; 
32'd149703: dataIn1 = 32'd2470
; 
32'd149704: dataIn1 = 32'd2472
; 
32'd149705: dataIn1 = 32'd4562
; 
32'd149706: dataIn1 = 32'd4563
; 
32'd149707: dataIn1 = 32'd4564
; 
32'd149708: dataIn1 = 32'd4567
; 
32'd149709: dataIn1 = 32'd4568
; 
32'd149710: dataIn1 = 32'd2470
; 
32'd149711: dataIn1 = 32'd2471
; 
32'd149712: dataIn1 = 32'd4562
; 
32'd149713: dataIn1 = 32'd4563
; 
32'd149714: dataIn1 = 32'd4564
; 
32'd149715: dataIn1 = 32'd4569
; 
32'd149716: dataIn1 = 32'd4570
; 
32'd149717: dataIn1 = 32'd375
; 
32'd149718: dataIn1 = 32'd2472
; 
32'd149719: dataIn1 = 32'd3366
; 
32'd149720: dataIn1 = 32'd4562
; 
32'd149721: dataIn1 = 32'd4565
; 
32'd149722: dataIn1 = 32'd4566
; 
32'd149723: dataIn1 = 32'd4574
; 
32'd149724: dataIn1 = 32'd375
; 
32'd149725: dataIn1 = 32'd2471
; 
32'd149726: dataIn1 = 32'd3373
; 
32'd149727: dataIn1 = 32'd4562
; 
32'd149728: dataIn1 = 32'd4565
; 
32'd149729: dataIn1 = 32'd4566
; 
32'd149730: dataIn1 = 32'd4571
; 
32'd149731: dataIn1 = 32'd501
; 
32'd149732: dataIn1 = 32'd2472
; 
32'd149733: dataIn1 = 32'd4563
; 
32'd149734: dataIn1 = 32'd4567
; 
32'd149735: dataIn1 = 32'd4568
; 
32'd149736: dataIn1 = 32'd4575
; 
32'd149737: dataIn1 = 32'd4577
; 
32'd149738: dataIn1 = 32'd501
; 
32'd149739: dataIn1 = 32'd2470
; 
32'd149740: dataIn1 = 32'd4563
; 
32'd149741: dataIn1 = 32'd4567
; 
32'd149742: dataIn1 = 32'd4568
; 
32'd149743: dataIn1 = 32'd5420
; 
32'd149744: dataIn1 = 32'd5421
; 
32'd149745: dataIn1 = 32'd500
; 
32'd149746: dataIn1 = 32'd2471
; 
32'd149747: dataIn1 = 32'd4561
; 
32'd149748: dataIn1 = 32'd4564
; 
32'd149749: dataIn1 = 32'd4569
; 
32'd149750: dataIn1 = 32'd4570
; 
32'd149751: dataIn1 = 32'd4573
; 
32'd149752: dataIn1 = 32'd500
; 
32'd149753: dataIn1 = 32'd2470
; 
32'd149754: dataIn1 = 32'd4564
; 
32'd149755: dataIn1 = 32'd4569
; 
32'd149756: dataIn1 = 32'd4570
; 
32'd149757: dataIn1 = 32'd5418
; 
32'd149758: dataIn1 = 32'd5420
; 
32'd149759: dataIn1 = 32'd2024
; 
32'd149760: dataIn1 = 32'd2471
; 
32'd149761: dataIn1 = 32'd3373
; 
32'd149762: dataIn1 = 32'd4566
; 
32'd149763: dataIn1 = 32'd4571
; 
32'd149764: dataIn1 = 32'd4572
; 
32'd149765: dataIn1 = 32'd4573
; 
32'd149766: dataIn1 = 32'd2024
; 
32'd149767: dataIn1 = 32'd2468
; 
32'd149768: dataIn1 = 32'd3374
; 
32'd149769: dataIn1 = 32'd4559
; 
32'd149770: dataIn1 = 32'd4571
; 
32'd149771: dataIn1 = 32'd4572
; 
32'd149772: dataIn1 = 32'd4573
; 
32'd149773: dataIn1 = 32'd2468
; 
32'd149774: dataIn1 = 32'd2471
; 
32'd149775: dataIn1 = 32'd4561
; 
32'd149776: dataIn1 = 32'd4569
; 
32'd149777: dataIn1 = 32'd4571
; 
32'd149778: dataIn1 = 32'd4572
; 
32'd149779: dataIn1 = 32'd4573
; 
32'd149780: dataIn1 = 32'd2023
; 
32'd149781: dataIn1 = 32'd2472
; 
32'd149782: dataIn1 = 32'd3366
; 
32'd149783: dataIn1 = 32'd4565
; 
32'd149784: dataIn1 = 32'd4574
; 
32'd149785: dataIn1 = 32'd4575
; 
32'd149786: dataIn1 = 32'd4576
; 
32'd149787: dataIn1 = 32'd2472
; 
32'd149788: dataIn1 = 32'd2473
; 
32'd149789: dataIn1 = 32'd4567
; 
32'd149790: dataIn1 = 32'd4574
; 
32'd149791: dataIn1 = 32'd4575
; 
32'd149792: dataIn1 = 32'd4576
; 
32'd149793: dataIn1 = 32'd4577
; 
32'd149794: dataIn1 = 32'd2023
; 
32'd149795: dataIn1 = 32'd2473
; 
32'd149796: dataIn1 = 32'd3369
; 
32'd149797: dataIn1 = 32'd4574
; 
32'd149798: dataIn1 = 32'd4575
; 
32'd149799: dataIn1 = 32'd4576
; 
32'd149800: dataIn1 = 32'd4585
; 
32'd149801: dataIn1 = 32'd501
; 
32'd149802: dataIn1 = 32'd2473
; 
32'd149803: dataIn1 = 32'd4567
; 
32'd149804: dataIn1 = 32'd4575
; 
32'd149805: dataIn1 = 32'd4577
; 
32'd149806: dataIn1 = 32'd4579
; 
32'd149807: dataIn1 = 32'd4583
; 
32'd149808: dataIn1 = 32'd2474
; 
32'd149809: dataIn1 = 32'd2475
; 
32'd149810: dataIn1 = 32'd4578
; 
32'd149811: dataIn1 = 32'd4579
; 
32'd149812: dataIn1 = 32'd4580
; 
32'd149813: dataIn1 = 32'd4581
; 
32'd149814: dataIn1 = 32'd4582
; 
32'd149815: dataIn1 = 32'd2473
; 
32'd149816: dataIn1 = 32'd2475
; 
32'd149817: dataIn1 = 32'd4577
; 
32'd149818: dataIn1 = 32'd4578
; 
32'd149819: dataIn1 = 32'd4579
; 
32'd149820: dataIn1 = 32'd4580
; 
32'd149821: dataIn1 = 32'd4583
; 
32'd149822: dataIn1 = 32'd2473
; 
32'd149823: dataIn1 = 32'd2474
; 
32'd149824: dataIn1 = 32'd4578
; 
32'd149825: dataIn1 = 32'd4579
; 
32'd149826: dataIn1 = 32'd4580
; 
32'd149827: dataIn1 = 32'd4584
; 
32'd149828: dataIn1 = 32'd4585
; 
32'd149829: dataIn1 = 32'd502
; 
32'd149830: dataIn1 = 32'd2475
; 
32'd149831: dataIn1 = 32'd4578
; 
32'd149832: dataIn1 = 32'd4581
; 
32'd149833: dataIn1 = 32'd4582
; 
32'd149834: dataIn1 = 32'd5422
; 
32'd149835: dataIn1 = 32'd5423
; 
32'd149836: dataIn1 = 32'd502
; 
32'd149837: dataIn1 = 32'd2474
; 
32'd149838: dataIn1 = 32'd4578
; 
32'd149839: dataIn1 = 32'd4581
; 
32'd149840: dataIn1 = 32'd4582
; 
32'd149841: dataIn1 = 32'd4589
; 
32'd149842: dataIn1 = 32'd4599
; 
32'd149843: dataIn1 = 32'd501
; 
32'd149844: dataIn1 = 32'd2475
; 
32'd149845: dataIn1 = 32'd4577
; 
32'd149846: dataIn1 = 32'd4579
; 
32'd149847: dataIn1 = 32'd4583
; 
32'd149848: dataIn1 = 32'd5421
; 
32'd149849: dataIn1 = 32'd5422
; 
32'd149850: dataIn1 = 32'd192
; 
32'd149851: dataIn1 = 32'd2474
; 
32'd149852: dataIn1 = 32'd3397
; 
32'd149853: dataIn1 = 32'd4580
; 
32'd149854: dataIn1 = 32'd4584
; 
32'd149855: dataIn1 = 32'd4585
; 
32'd149856: dataIn1 = 32'd4601
; 
32'd149857: dataIn1 = 32'd192
; 
32'd149858: dataIn1 = 32'd2473
; 
32'd149859: dataIn1 = 32'd3369
; 
32'd149860: dataIn1 = 32'd4576
; 
32'd149861: dataIn1 = 32'd4580
; 
32'd149862: dataIn1 = 32'd4584
; 
32'd149863: dataIn1 = 32'd4585
; 
32'd149864: dataIn1 = 32'd2477
; 
32'd149865: dataIn1 = 32'd2478
; 
32'd149866: dataIn1 = 32'd4586
; 
32'd149867: dataIn1 = 32'd4587
; 
32'd149868: dataIn1 = 32'd4588
; 
32'd149869: dataIn1 = 32'd4589
; 
32'd149870: dataIn1 = 32'd4590
; 
32'd149871: dataIn1 = 32'd2476
; 
32'd149872: dataIn1 = 32'd2478
; 
32'd149873: dataIn1 = 32'd4586
; 
32'd149874: dataIn1 = 32'd4587
; 
32'd149875: dataIn1 = 32'd4588
; 
32'd149876: dataIn1 = 32'd4591
; 
32'd149877: dataIn1 = 32'd4592
; 
32'd149878: dataIn1 = 32'd2476
; 
32'd149879: dataIn1 = 32'd2477
; 
32'd149880: dataIn1 = 32'd4586
; 
32'd149881: dataIn1 = 32'd4587
; 
32'd149882: dataIn1 = 32'd4588
; 
32'd149883: dataIn1 = 32'd4593
; 
32'd149884: dataIn1 = 32'd4594
; 
32'd149885: dataIn1 = 32'd502
; 
32'd149886: dataIn1 = 32'd2478
; 
32'd149887: dataIn1 = 32'd4582
; 
32'd149888: dataIn1 = 32'd4586
; 
32'd149889: dataIn1 = 32'd4589
; 
32'd149890: dataIn1 = 32'd4590
; 
32'd149891: dataIn1 = 32'd4599
; 
32'd149892: dataIn1 = 32'd502
; 
32'd149893: dataIn1 = 32'd2477
; 
32'd149894: dataIn1 = 32'd4586
; 
32'd149895: dataIn1 = 32'd4589
; 
32'd149896: dataIn1 = 32'd4590
; 
32'd149897: dataIn1 = 32'd5423
; 
32'd149898: dataIn1 = 32'd5425
; 
32'd149899: dataIn1 = 32'd382
; 
32'd149900: dataIn1 = 32'd2478
; 
32'd149901: dataIn1 = 32'd3396
; 
32'd149902: dataIn1 = 32'd4587
; 
32'd149903: dataIn1 = 32'd4591
; 
32'd149904: dataIn1 = 32'd4592
; 
32'd149905: dataIn1 = 32'd4600
; 
32'd149906: dataIn1 = 32'd382
; 
32'd149907: dataIn1 = 32'd2476
; 
32'd149908: dataIn1 = 32'd3402
; 
32'd149909: dataIn1 = 32'd4587
; 
32'd149910: dataIn1 = 32'd4591
; 
32'd149911: dataIn1 = 32'd4592
; 
32'd149912: dataIn1 = 32'd4596
; 
32'd149913: dataIn1 = 32'd503
; 
32'd149914: dataIn1 = 32'd2477
; 
32'd149915: dataIn1 = 32'd4588
; 
32'd149916: dataIn1 = 32'd4593
; 
32'd149917: dataIn1 = 32'd4594
; 
32'd149918: dataIn1 = 32'd5424
; 
32'd149919: dataIn1 = 32'd5425
; 
32'd149920: dataIn1 = 32'd503
; 
32'd149921: dataIn1 = 32'd2476
; 
32'd149922: dataIn1 = 32'd4588
; 
32'd149923: dataIn1 = 32'd4593
; 
32'd149924: dataIn1 = 32'd4594
; 
32'd149925: dataIn1 = 32'd4597
; 
32'd149926: dataIn1 = 32'd4598
; 
32'd149927: dataIn1 = 32'd2028
; 
32'd149928: dataIn1 = 32'd2479
; 
32'd149929: dataIn1 = 32'd3401
; 
32'd149930: dataIn1 = 32'd4595
; 
32'd149931: dataIn1 = 32'd4596
; 
32'd149932: dataIn1 = 32'd4597
; 
32'd149933: dataIn1 = 32'd5305
; 
32'd149934: dataIn1 = 32'd2028
; 
32'd149935: dataIn1 = 32'd2476
; 
32'd149936: dataIn1 = 32'd3402
; 
32'd149937: dataIn1 = 32'd4592
; 
32'd149938: dataIn1 = 32'd4595
; 
32'd149939: dataIn1 = 32'd4596
; 
32'd149940: dataIn1 = 32'd4597
; 
32'd149941: dataIn1 = 32'd2476
; 
32'd149942: dataIn1 = 32'd2479
; 
32'd149943: dataIn1 = 32'd4594
; 
32'd149944: dataIn1 = 32'd4595
; 
32'd149945: dataIn1 = 32'd4596
; 
32'd149946: dataIn1 = 32'd4597
; 
32'd149947: dataIn1 = 32'd4598
; 
32'd149948: dataIn1 = 32'd503
; 
32'd149949: dataIn1 = 32'd2479
; 
32'd149950: dataIn1 = 32'd4594
; 
32'd149951: dataIn1 = 32'd4597
; 
32'd149952: dataIn1 = 32'd4598
; 
32'd149953: dataIn1 = 32'd2474
; 
32'd149954: dataIn1 = 32'd2478
; 
32'd149955: dataIn1 = 32'd4582
; 
32'd149956: dataIn1 = 32'd4589
; 
32'd149957: dataIn1 = 32'd4599
; 
32'd149958: dataIn1 = 32'd4600
; 
32'd149959: dataIn1 = 32'd4601
; 
32'd149960: dataIn1 = 32'd2027
; 
32'd149961: dataIn1 = 32'd2478
; 
32'd149962: dataIn1 = 32'd3396
; 
32'd149963: dataIn1 = 32'd4591
; 
32'd149964: dataIn1 = 32'd4599
; 
32'd149965: dataIn1 = 32'd4600
; 
32'd149966: dataIn1 = 32'd4601
; 
32'd149967: dataIn1 = 32'd2027
; 
32'd149968: dataIn1 = 32'd2474
; 
32'd149969: dataIn1 = 32'd3397
; 
32'd149970: dataIn1 = 32'd4584
; 
32'd149971: dataIn1 = 32'd4599
; 
32'd149972: dataIn1 = 32'd4600
; 
32'd149973: dataIn1 = 32'd4601
; 
32'd149974: dataIn1 = 32'd205
; 
32'd149975: dataIn1 = 32'd396
; 
32'd149976: dataIn1 = 32'd751
; 
32'd149977: dataIn1 = 32'd2489
; 
32'd149978: dataIn1 = 32'd3897
; 
32'd149979: dataIn1 = 32'd4602
; 
32'd149980: dataIn1 = 32'd5426
; 
32'd149981: dataIn1 = 32'd128
; 
32'd149982: dataIn1 = 32'd405
; 
32'd149983: dataIn1 = 32'd774
; 
32'd149984: dataIn1 = 32'd2490
; 
32'd149985: dataIn1 = 32'd3926
; 
32'd149986: dataIn1 = 32'd4603
; 
32'd149987: dataIn1 = 32'd5427
; 
32'd149988: dataIn1 = 32'd131
; 
32'd149989: dataIn1 = 32'd2532
; 
32'd149990: dataIn1 = 32'd4604
; 
32'd149991: dataIn1 = 32'd4605
; 
32'd149992: dataIn1 = 32'd4606
; 
32'd149993: dataIn1 = 32'd4619
; 
32'd149994: dataIn1 = 32'd4621
; 
32'd149995: dataIn1 = 32'd131
; 
32'd149996: dataIn1 = 32'd2531
; 
32'd149997: dataIn1 = 32'd4604
; 
32'd149998: dataIn1 = 32'd4605
; 
32'd149999: dataIn1 = 32'd4606
; 
32'd150000: dataIn1 = 32'd4632
; 
32'd150001: dataIn1 = 32'd4635
; 
32'd150002: dataIn1 = 32'd2051
; 
32'd150003: dataIn1 = 32'd2531
; 
32'd150004: dataIn1 = 32'd2532
; 
32'd150005: dataIn1 = 32'd4604
; 
32'd150006: dataIn1 = 32'd4605
; 
32'd150007: dataIn1 = 32'd4606
; 
32'd150008: dataIn1 = 32'd2287
; 
32'd150009: dataIn1 = 32'd2535
; 
32'd150010: dataIn1 = 32'd3864
; 
32'd150011: dataIn1 = 32'd4607
; 
32'd150012: dataIn1 = 32'd4608
; 
32'd150013: dataIn1 = 32'd4609
; 
32'd150014: dataIn1 = 32'd4610
; 
32'd150015: dataIn1 = 32'd2287
; 
32'd150016: dataIn1 = 32'd2533
; 
32'd150017: dataIn1 = 32'd4607
; 
32'd150018: dataIn1 = 32'd4608
; 
32'd150019: dataIn1 = 32'd4609
; 
32'd150020: dataIn1 = 32'd4611
; 
32'd150021: dataIn1 = 32'd4612
; 
32'd150022: dataIn1 = 32'd1039
; 
32'd150023: dataIn1 = 32'd2533
; 
32'd150024: dataIn1 = 32'd2535
; 
32'd150025: dataIn1 = 32'd4607
; 
32'd150026: dataIn1 = 32'd4608
; 
32'd150027: dataIn1 = 32'd4609
; 
32'd150028: dataIn1 = 32'd126
; 
32'd150029: dataIn1 = 32'd2535
; 
32'd150030: dataIn1 = 32'd3864
; 
32'd150031: dataIn1 = 32'd4607
; 
32'd150032: dataIn1 = 32'd4610
; 
32'd150033: dataIn1 = 32'd5952
; 
32'd150034: dataIn1 = 32'd6698
; 
32'd150035: dataIn1 = 32'd391
; 
32'd150036: dataIn1 = 32'd2287
; 
32'd150037: dataIn1 = 32'd4608
; 
32'd150038: dataIn1 = 32'd4611
; 
32'd150039: dataIn1 = 32'd4612
; 
32'd150040: dataIn1 = 32'd10257
; 
32'd150041: dataIn1 = 32'd10263
; 
32'd150042: dataIn1 = 32'd391
; 
32'd150043: dataIn1 = 32'd2533
; 
32'd150044: dataIn1 = 32'd3408
; 
32'd150045: dataIn1 = 32'd4608
; 
32'd150046: dataIn1 = 32'd4611
; 
32'd150047: dataIn1 = 32'd4612
; 
32'd150048: dataIn1 = 32'd5306
; 
32'd150049: dataIn1 = 32'd1041
; 
32'd150050: dataIn1 = 32'd2541
; 
32'd150051: dataIn1 = 32'd4613
; 
32'd150052: dataIn1 = 32'd4614
; 
32'd150053: dataIn1 = 32'd4615
; 
32'd150054: dataIn1 = 32'd4620
; 
32'd150055: dataIn1 = 32'd4622
; 
32'd150056: dataIn1 = 32'd1041
; 
32'd150057: dataIn1 = 32'd2540
; 
32'd150058: dataIn1 = 32'd4613
; 
32'd150059: dataIn1 = 32'd4614
; 
32'd150060: dataIn1 = 32'd4615
; 
32'd150061: dataIn1 = 32'd4616
; 
32'd150062: dataIn1 = 32'd4617
; 
32'd150063: dataIn1 = 32'd2047
; 
32'd150064: dataIn1 = 32'd2540
; 
32'd150065: dataIn1 = 32'd2541
; 
32'd150066: dataIn1 = 32'd4613
; 
32'd150067: dataIn1 = 32'd4614
; 
32'd150068: dataIn1 = 32'd4615
; 
32'd150069: dataIn1 = 32'd1041
; 
32'd150070: dataIn1 = 32'd2542
; 
32'd150071: dataIn1 = 32'd4614
; 
32'd150072: dataIn1 = 32'd4616
; 
32'd150073: dataIn1 = 32'd4617
; 
32'd150074: dataIn1 = 32'd5915
; 
32'd150075: dataIn1 = 32'd5919
; 
32'd150076: dataIn1 = 32'd2530
; 
32'd150077: dataIn1 = 32'd2540
; 
32'd150078: dataIn1 = 32'd2542
; 
32'd150079: dataIn1 = 32'd4614
; 
32'd150080: dataIn1 = 32'd4616
; 
32'd150081: dataIn1 = 32'd4617
; 
32'd150082: dataIn1 = 32'd982
; 
32'd150083: dataIn1 = 32'd2532
; 
32'd150084: dataIn1 = 32'd2541
; 
32'd150085: dataIn1 = 32'd4618
; 
32'd150086: dataIn1 = 32'd4619
; 
32'd150087: dataIn1 = 32'd4620
; 
32'd150088: dataIn1 = 32'd2532
; 
32'd150089: dataIn1 = 32'd2543
; 
32'd150090: dataIn1 = 32'd4604
; 
32'd150091: dataIn1 = 32'd4618
; 
32'd150092: dataIn1 = 32'd4619
; 
32'd150093: dataIn1 = 32'd4620
; 
32'd150094: dataIn1 = 32'd4621
; 
32'd150095: dataIn1 = 32'd2541
; 
32'd150096: dataIn1 = 32'd2543
; 
32'd150097: dataIn1 = 32'd4613
; 
32'd150098: dataIn1 = 32'd4618
; 
32'd150099: dataIn1 = 32'd4619
; 
32'd150100: dataIn1 = 32'd4620
; 
32'd150101: dataIn1 = 32'd4622
; 
32'd150102: dataIn1 = 32'd131
; 
32'd150103: dataIn1 = 32'd2543
; 
32'd150104: dataIn1 = 32'd4604
; 
32'd150105: dataIn1 = 32'd4619
; 
32'd150106: dataIn1 = 32'd4621
; 
32'd150107: dataIn1 = 32'd5922
; 
32'd150108: dataIn1 = 32'd5980
; 
32'd150109: dataIn1 = 32'd1041
; 
32'd150110: dataIn1 = 32'd2543
; 
32'd150111: dataIn1 = 32'd4613
; 
32'd150112: dataIn1 = 32'd4620
; 
32'd150113: dataIn1 = 32'd4622
; 
32'd150114: dataIn1 = 32'd5914
; 
32'd150115: dataIn1 = 32'd5923
; 
32'd150116: dataIn1 = 32'd2544
; 
32'd150117: dataIn1 = 32'd2545
; 
32'd150118: dataIn1 = 32'd4623
; 
32'd150119: dataIn1 = 32'd4624
; 
32'd150120: dataIn1 = 32'd4625
; 
32'd150121: dataIn1 = 32'd4626
; 
32'd150122: dataIn1 = 32'd4627
; 
32'd150123: dataIn1 = 32'd2048
; 
32'd150124: dataIn1 = 32'd2545
; 
32'd150125: dataIn1 = 32'd4623
; 
32'd150126: dataIn1 = 32'd4624
; 
32'd150127: dataIn1 = 32'd4625
; 
32'd150128: dataIn1 = 32'd4628
; 
32'd150129: dataIn1 = 32'd4629
; 
32'd150130: dataIn1 = 32'd2048
; 
32'd150131: dataIn1 = 32'd2544
; 
32'd150132: dataIn1 = 32'd3417
; 
32'd150133: dataIn1 = 32'd4623
; 
32'd150134: dataIn1 = 32'd4624
; 
32'd150135: dataIn1 = 32'd4625
; 
32'd150136: dataIn1 = 32'd5307
; 
32'd150137: dataIn1 = 32'd1042
; 
32'd150138: dataIn1 = 32'd2545
; 
32'd150139: dataIn1 = 32'd4623
; 
32'd150140: dataIn1 = 32'd4626
; 
32'd150141: dataIn1 = 32'd4627
; 
32'd150142: dataIn1 = 32'd4630
; 
32'd150143: dataIn1 = 32'd4633
; 
32'd150144: dataIn1 = 32'd1042
; 
32'd150145: dataIn1 = 32'd2544
; 
32'd150146: dataIn1 = 32'd4623
; 
32'd150147: dataIn1 = 32'd4626
; 
32'd150148: dataIn1 = 32'd4627
; 
32'd150149: dataIn1 = 32'd5429
; 
32'd150150: dataIn1 = 32'd983
; 
32'd150151: dataIn1 = 32'd2545
; 
32'd150152: dataIn1 = 32'd4624
; 
32'd150153: dataIn1 = 32'd4628
; 
32'd150154: dataIn1 = 32'd4629
; 
32'd150155: dataIn1 = 32'd4631
; 
32'd150156: dataIn1 = 32'd4634
; 
32'd150157: dataIn1 = 32'd983
; 
32'd150158: dataIn1 = 32'd2048
; 
32'd150159: dataIn1 = 32'd4624
; 
32'd150160: dataIn1 = 32'd4628
; 
32'd150161: dataIn1 = 32'd4629
; 
32'd150162: dataIn1 = 32'd10261
; 
32'd150163: dataIn1 = 32'd10273
; 
32'd150164: dataIn1 = 32'd2545
; 
32'd150165: dataIn1 = 32'd2546
; 
32'd150166: dataIn1 = 32'd4626
; 
32'd150167: dataIn1 = 32'd4630
; 
32'd150168: dataIn1 = 32'd4631
; 
32'd150169: dataIn1 = 32'd4632
; 
32'd150170: dataIn1 = 32'd4633
; 
32'd150171: dataIn1 = 32'd2531
; 
32'd150172: dataIn1 = 32'd2545
; 
32'd150173: dataIn1 = 32'd4628
; 
32'd150174: dataIn1 = 32'd4630
; 
32'd150175: dataIn1 = 32'd4631
; 
32'd150176: dataIn1 = 32'd4632
; 
32'd150177: dataIn1 = 32'd4634
; 
32'd150178: dataIn1 = 32'd2531
; 
32'd150179: dataIn1 = 32'd2546
; 
32'd150180: dataIn1 = 32'd4605
; 
32'd150181: dataIn1 = 32'd4630
; 
32'd150182: dataIn1 = 32'd4631
; 
32'd150183: dataIn1 = 32'd4632
; 
32'd150184: dataIn1 = 32'd4635
; 
32'd150185: dataIn1 = 32'd1042
; 
32'd150186: dataIn1 = 32'd2546
; 
32'd150187: dataIn1 = 32'd4626
; 
32'd150188: dataIn1 = 32'd4630
; 
32'd150189: dataIn1 = 32'd4633
; 
32'd150190: dataIn1 = 32'd4683
; 
32'd150191: dataIn1 = 32'd983
; 
32'd150192: dataIn1 = 32'd2051
; 
32'd150193: dataIn1 = 32'd2531
; 
32'd150194: dataIn1 = 32'd4628
; 
32'd150195: dataIn1 = 32'd4631
; 
32'd150196: dataIn1 = 32'd4634
; 
32'd150197: dataIn1 = 32'd131
; 
32'd150198: dataIn1 = 32'd2546
; 
32'd150199: dataIn1 = 32'd4605
; 
32'd150200: dataIn1 = 32'd4632
; 
32'd150201: dataIn1 = 32'd4635
; 
32'd150202: dataIn1 = 32'd5982
; 
32'd150203: dataIn1 = 32'd6699
; 
32'd150204: dataIn1 = 32'd3
; 
32'd150205: dataIn1 = 32'd2549
; 
32'd150206: dataIn1 = 32'd4636
; 
32'd150207: dataIn1 = 32'd4637
; 
32'd150208: dataIn1 = 32'd4638
; 
32'd150209: dataIn1 = 32'd1068
; 
32'd150210: dataIn1 = 32'd2547
; 
32'd150211: dataIn1 = 32'd2548
; 
32'd150212: dataIn1 = 32'd2549
; 
32'd150213: dataIn1 = 32'd4636
; 
32'd150214: dataIn1 = 32'd4637
; 
32'd150215: dataIn1 = 32'd4638
; 
32'd150216: dataIn1 = 32'd3
; 
32'd150217: dataIn1 = 32'd2547
; 
32'd150218: dataIn1 = 32'd4636
; 
32'd150219: dataIn1 = 32'd4637
; 
32'd150220: dataIn1 = 32'd4638
; 
32'd150221: dataIn1 = 32'd4801
; 
32'd150222: dataIn1 = 32'd4803
; 
32'd150223: dataIn1 = 32'd9689
; 
32'd150224: dataIn1 = 32'd2550
; 
32'd150225: dataIn1 = 32'd2551
; 
32'd150226: dataIn1 = 32'd2552
; 
32'd150227: dataIn1 = 32'd4639
; 
32'd150228: dataIn1 = 32'd4640
; 
32'd150229: dataIn1 = 32'd4641
; 
32'd150230: dataIn1 = 32'd124
; 
32'd150231: dataIn1 = 32'd2552
; 
32'd150232: dataIn1 = 32'd4639
; 
32'd150233: dataIn1 = 32'd4640
; 
32'd150234: dataIn1 = 32'd4641
; 
32'd150235: dataIn1 = 32'd4795
; 
32'd150236: dataIn1 = 32'd4798
; 
32'd150237: dataIn1 = 32'd9704
; 
32'd150238: dataIn1 = 32'd124
; 
32'd150239: dataIn1 = 32'd2551
; 
32'd150240: dataIn1 = 32'd4639
; 
32'd150241: dataIn1 = 32'd4640
; 
32'd150242: dataIn1 = 32'd4641
; 
32'd150243: dataIn1 = 32'd4808
; 
32'd150244: dataIn1 = 32'd4811
; 
32'd150245: dataIn1 = 32'd9724
; 
32'd150246: dataIn1 = 32'd1039
; 
32'd150247: dataIn1 = 32'd2535
; 
32'd150248: dataIn1 = 32'd2553
; 
32'd150249: dataIn1 = 32'd2554
; 
32'd150250: dataIn1 = 32'd4642
; 
32'd150251: dataIn1 = 32'd4643
; 
32'd150252: dataIn1 = 32'd6698
; 
32'd150253: dataIn1 = 32'd2554
; 
32'd150254: dataIn1 = 32'd4642
; 
32'd150255: dataIn1 = 32'd4643
; 
32'd150256: dataIn1 = 32'd5948
; 
32'd150257: dataIn1 = 32'd5949
; 
32'd150258: dataIn1 = 32'd5952
; 
32'd150259: dataIn1 = 32'd6698
; 
32'd150260: dataIn1 = 32'd4
; 
32'd150261: dataIn1 = 32'd2557
; 
32'd150262: dataIn1 = 32'd4644
; 
32'd150263: dataIn1 = 32'd4645
; 
32'd150264: dataIn1 = 32'd4646
; 
32'd150265: dataIn1 = 32'd4815
; 
32'd150266: dataIn1 = 32'd4817
; 
32'd150267: dataIn1 = 32'd2555
; 
32'd150268: dataIn1 = 32'd2556
; 
32'd150269: dataIn1 = 32'd2557
; 
32'd150270: dataIn1 = 32'd4644
; 
32'd150271: dataIn1 = 32'd4645
; 
32'd150272: dataIn1 = 32'd4646
; 
32'd150273: dataIn1 = 32'd4
; 
32'd150274: dataIn1 = 32'd2555
; 
32'd150275: dataIn1 = 32'd4644
; 
32'd150276: dataIn1 = 32'd4645
; 
32'd150277: dataIn1 = 32'd4646
; 
32'd150278: dataIn1 = 32'd4833
; 
32'd150279: dataIn1 = 32'd4836
; 
32'd150280: dataIn1 = 32'd2559
; 
32'd150281: dataIn1 = 32'd2560
; 
32'd150282: dataIn1 = 32'd4647
; 
32'd150283: dataIn1 = 32'd4648
; 
32'd150284: dataIn1 = 32'd4649
; 
32'd150285: dataIn1 = 32'd4650
; 
32'd150286: dataIn1 = 32'd4651
; 
32'd150287: dataIn1 = 32'd5889
; 
32'd150288: dataIn1 = 32'd2558
; 
32'd150289: dataIn1 = 32'd2560
; 
32'd150290: dataIn1 = 32'd4647
; 
32'd150291: dataIn1 = 32'd4648
; 
32'd150292: dataIn1 = 32'd4649
; 
32'd150293: dataIn1 = 32'd4652
; 
32'd150294: dataIn1 = 32'd4653
; 
32'd150295: dataIn1 = 32'd2558
; 
32'd150296: dataIn1 = 32'd2559
; 
32'd150297: dataIn1 = 32'd4647
; 
32'd150298: dataIn1 = 32'd4648
; 
32'd150299: dataIn1 = 32'd4649
; 
32'd150300: dataIn1 = 32'd4654
; 
32'd150301: dataIn1 = 32'd4655
; 
32'd150302: dataIn1 = 32'd2560
; 
32'd150303: dataIn1 = 32'd4647
; 
32'd150304: dataIn1 = 32'd4650
; 
32'd150305: dataIn1 = 32'd5889
; 
32'd150306: dataIn1 = 32'd5891
; 
32'd150307: dataIn1 = 32'd5927
; 
32'd150308: dataIn1 = 32'd5929
; 
32'd150309: dataIn1 = 32'd2559
; 
32'd150310: dataIn1 = 32'd4647
; 
32'd150311: dataIn1 = 32'd4651
; 
32'd150312: dataIn1 = 32'd5889
; 
32'd150313: dataIn1 = 32'd5890
; 
32'd150314: dataIn1 = 32'd5917
; 
32'd150315: dataIn1 = 32'd5918
; 
32'd150316: dataIn1 = 32'd1074
; 
32'd150317: dataIn1 = 32'd2560
; 
32'd150318: dataIn1 = 32'd4648
; 
32'd150319: dataIn1 = 32'd4652
; 
32'd150320: dataIn1 = 32'd4653
; 
32'd150321: dataIn1 = 32'd4669
; 
32'd150322: dataIn1 = 32'd4671
; 
32'd150323: dataIn1 = 32'd5909
; 
32'd150324: dataIn1 = 32'd2558
; 
32'd150325: dataIn1 = 32'd4648
; 
32'd150326: dataIn1 = 32'd4652
; 
32'd150327: dataIn1 = 32'd4653
; 
32'd150328: dataIn1 = 32'd5906
; 
32'd150329: dataIn1 = 32'd5907
; 
32'd150330: dataIn1 = 32'd5909
; 
32'd150331: dataIn1 = 32'd1075
; 
32'd150332: dataIn1 = 32'd2559
; 
32'd150333: dataIn1 = 32'd4649
; 
32'd150334: dataIn1 = 32'd4654
; 
32'd150335: dataIn1 = 32'd4655
; 
32'd150336: dataIn1 = 32'd4665
; 
32'd150337: dataIn1 = 32'd4667
; 
32'd150338: dataIn1 = 32'd1075
; 
32'd150339: dataIn1 = 32'd2558
; 
32'd150340: dataIn1 = 32'd4649
; 
32'd150341: dataIn1 = 32'd4654
; 
32'd150342: dataIn1 = 32'd4655
; 
32'd150343: dataIn1 = 32'd4658
; 
32'd150344: dataIn1 = 32'd4662
; 
32'd150345: dataIn1 = 32'd5912
; 
32'd150346: dataIn1 = 32'd4656
; 
32'd150347: dataIn1 = 32'd5893
; 
32'd150348: dataIn1 = 32'd5894
; 
32'd150349: dataIn1 = 32'd5896
; 
32'd150350: dataIn1 = 32'd5898
; 
32'd150351: dataIn1 = 32'd5900
; 
32'd150352: dataIn1 = 32'd5901
; 
32'd150353: dataIn1 = 32'd2558
; 
32'd150354: dataIn1 = 32'd4657
; 
32'd150355: dataIn1 = 32'd5892
; 
32'd150356: dataIn1 = 32'd5894
; 
32'd150357: dataIn1 = 32'd5897
; 
32'd150358: dataIn1 = 32'd5906
; 
32'd150359: dataIn1 = 32'd5908
; 
32'd150360: dataIn1 = 32'd2558
; 
32'd150361: dataIn1 = 32'd4655
; 
32'd150362: dataIn1 = 32'd4658
; 
32'd150363: dataIn1 = 32'd5892
; 
32'd150364: dataIn1 = 32'd5893
; 
32'd150365: dataIn1 = 32'd5895
; 
32'd150366: dataIn1 = 32'd5912
; 
32'd150367: dataIn1 = 32'd4659
; 
32'd150368: dataIn1 = 32'd5899
; 
32'd150369: dataIn1 = 32'd5901
; 
32'd150370: dataIn1 = 32'd5903
; 
32'd150371: dataIn1 = 32'd5905
; 
32'd150372: dataIn1 = 32'd6030
; 
32'd150373: dataIn1 = 32'd6032
; 
32'd150374: dataIn1 = 32'd4660
; 
32'd150375: dataIn1 = 32'd5899
; 
32'd150376: dataIn1 = 32'd5900
; 
32'd150377: dataIn1 = 32'd5902
; 
32'd150378: dataIn1 = 32'd5904
; 
32'd150379: dataIn1 = 32'd5969
; 
32'd150380: dataIn1 = 32'd5970
; 
32'd150381: dataIn1 = 32'd4661
; 
32'd150382: dataIn1 = 32'd5907
; 
32'd150383: dataIn1 = 32'd5908
; 
32'd150384: dataIn1 = 32'd5910
; 
32'd150385: dataIn1 = 32'd5911
; 
32'd150386: dataIn1 = 32'd6036
; 
32'd150387: dataIn1 = 32'd6037
; 
32'd150388: dataIn1 = 32'd1075
; 
32'd150389: dataIn1 = 32'd4655
; 
32'd150390: dataIn1 = 32'd4662
; 
32'd150391: dataIn1 = 32'd4847
; 
32'd150392: dataIn1 = 32'd5912
; 
32'd150393: dataIn1 = 32'd5913
; 
32'd150394: dataIn1 = 32'd5979
; 
32'd150395: dataIn1 = 32'd2559
; 
32'd150396: dataIn1 = 32'd4663
; 
32'd150397: dataIn1 = 32'd4665
; 
32'd150398: dataIn1 = 32'd5915
; 
32'd150399: dataIn1 = 32'd5916
; 
32'd150400: dataIn1 = 32'd5918
; 
32'd150401: dataIn1 = 32'd5919
; 
32'd150402: dataIn1 = 32'd2563
; 
32'd150403: dataIn1 = 32'd4664
; 
32'd150404: dataIn1 = 32'd4665
; 
32'd150405: dataIn1 = 32'd5914
; 
32'd150406: dataIn1 = 32'd5916
; 
32'd150407: dataIn1 = 32'd5921
; 
32'd150408: dataIn1 = 32'd5923
; 
32'd150409: dataIn1 = 32'd2559
; 
32'd150410: dataIn1 = 32'd2563
; 
32'd150411: dataIn1 = 32'd4654
; 
32'd150412: dataIn1 = 32'd4663
; 
32'd150413: dataIn1 = 32'd4664
; 
32'd150414: dataIn1 = 32'd4665
; 
32'd150415: dataIn1 = 32'd4667
; 
32'd150416: dataIn1 = 32'd5916
; 
32'd150417: dataIn1 = 32'd2563
; 
32'd150418: dataIn1 = 32'd4666
; 
32'd150419: dataIn1 = 32'd4854
; 
32'd150420: dataIn1 = 32'd5921
; 
32'd150421: dataIn1 = 32'd5922
; 
32'd150422: dataIn1 = 32'd5980
; 
32'd150423: dataIn1 = 32'd5981
; 
32'd150424: dataIn1 = 32'd1075
; 
32'd150425: dataIn1 = 32'd2563
; 
32'd150426: dataIn1 = 32'd4654
; 
32'd150427: dataIn1 = 32'd4665
; 
32'd150428: dataIn1 = 32'd4667
; 
32'd150429: dataIn1 = 32'd4846
; 
32'd150430: dataIn1 = 32'd4855
; 
32'd150431: dataIn1 = 32'd2560
; 
32'd150432: dataIn1 = 32'd4668
; 
32'd150433: dataIn1 = 32'd4669
; 
32'd150434: dataIn1 = 32'd5925
; 
32'd150435: dataIn1 = 32'd5926
; 
32'd150436: dataIn1 = 32'd5928
; 
32'd150437: dataIn1 = 32'd5929
; 
32'd150438: dataIn1 = 32'd2560
; 
32'd150439: dataIn1 = 32'd2564
; 
32'd150440: dataIn1 = 32'd4652
; 
32'd150441: dataIn1 = 32'd4668
; 
32'd150442: dataIn1 = 32'd4669
; 
32'd150443: dataIn1 = 32'd4670
; 
32'd150444: dataIn1 = 32'd4671
; 
32'd150445: dataIn1 = 32'd5925
; 
32'd150446: dataIn1 = 32'd2564
; 
32'd150447: dataIn1 = 32'd4669
; 
32'd150448: dataIn1 = 32'd4670
; 
32'd150449: dataIn1 = 32'd5924
; 
32'd150450: dataIn1 = 32'd5925
; 
32'd150451: dataIn1 = 32'd5932
; 
32'd150452: dataIn1 = 32'd5933
; 
32'd150453: dataIn1 = 32'd1074
; 
32'd150454: dataIn1 = 32'd2564
; 
32'd150455: dataIn1 = 32'd4652
; 
32'd150456: dataIn1 = 32'd4669
; 
32'd150457: dataIn1 = 32'd4671
; 
32'd150458: dataIn1 = 32'd4867
; 
32'd150459: dataIn1 = 32'd4882
; 
32'd150460: dataIn1 = 32'd6702
; 
32'd150461: dataIn1 = 32'd2564
; 
32'd150462: dataIn1 = 32'd4672
; 
32'd150463: dataIn1 = 32'd5932
; 
32'd150464: dataIn1 = 32'd5934
; 
32'd150465: dataIn1 = 32'd5936
; 
32'd150466: dataIn1 = 32'd6061
; 
32'd150467: dataIn1 = 32'd6063
; 
32'd150468: dataIn1 = 32'd2566
; 
32'd150469: dataIn1 = 32'd2569
; 
32'd150470: dataIn1 = 32'd4673
; 
32'd150471: dataIn1 = 32'd4674
; 
32'd150472: dataIn1 = 32'd4675
; 
32'd150473: dataIn1 = 32'd4676
; 
32'd150474: dataIn1 = 32'd4677
; 
32'd150475: dataIn1 = 32'd2568
; 
32'd150476: dataIn1 = 32'd2569
; 
32'd150477: dataIn1 = 32'd4673
; 
32'd150478: dataIn1 = 32'd4674
; 
32'd150479: dataIn1 = 32'd4675
; 
32'd150480: dataIn1 = 32'd4678
; 
32'd150481: dataIn1 = 32'd4679
; 
32'd150482: dataIn1 = 32'd5939
; 
32'd150483: dataIn1 = 32'd2566
; 
32'd150484: dataIn1 = 32'd2568
; 
32'd150485: dataIn1 = 32'd4673
; 
32'd150486: dataIn1 = 32'd4674
; 
32'd150487: dataIn1 = 32'd4675
; 
32'd150488: dataIn1 = 32'd4680
; 
32'd150489: dataIn1 = 32'd4681
; 
32'd150490: dataIn1 = 32'd1076
; 
32'd150491: dataIn1 = 32'd2569
; 
32'd150492: dataIn1 = 32'd4673
; 
32'd150493: dataIn1 = 32'd4676
; 
32'd150494: dataIn1 = 32'd4677
; 
32'd150495: dataIn1 = 32'd4842
; 
32'd150496: dataIn1 = 32'd4857
; 
32'd150497: dataIn1 = 32'd1076
; 
32'd150498: dataIn1 = 32'd2566
; 
32'd150499: dataIn1 = 32'd4673
; 
32'd150500: dataIn1 = 32'd4676
; 
32'd150501: dataIn1 = 32'd4677
; 
32'd150502: dataIn1 = 32'd10268
; 
32'd150503: dataIn1 = 32'd10274
; 
32'd150504: dataIn1 = 32'd2569
; 
32'd150505: dataIn1 = 32'd4674
; 
32'd150506: dataIn1 = 32'd4678
; 
32'd150507: dataIn1 = 32'd5939
; 
32'd150508: dataIn1 = 32'd5940
; 
32'd150509: dataIn1 = 32'd5992
; 
32'd150510: dataIn1 = 32'd5993
; 
32'd150511: dataIn1 = 32'd2568
; 
32'd150512: dataIn1 = 32'd4674
; 
32'd150513: dataIn1 = 32'd4679
; 
32'd150514: dataIn1 = 32'd4899
; 
32'd150515: dataIn1 = 32'd5938
; 
32'd150516: dataIn1 = 32'd5939
; 
32'd150517: dataIn1 = 32'd6066
; 
32'd150518: dataIn1 = 32'd1077
; 
32'd150519: dataIn1 = 32'd2565
; 
32'd150520: dataIn1 = 32'd2566
; 
32'd150521: dataIn1 = 32'd4675
; 
32'd150522: dataIn1 = 32'd4680
; 
32'd150523: dataIn1 = 32'd4681
; 
32'd150524: dataIn1 = 32'd1077
; 
32'd150525: dataIn1 = 32'd2568
; 
32'd150526: dataIn1 = 32'd4675
; 
32'd150527: dataIn1 = 32'd4680
; 
32'd150528: dataIn1 = 32'd4681
; 
32'd150529: dataIn1 = 32'd4888
; 
32'd150530: dataIn1 = 32'd4898
; 
32'd150531: dataIn1 = 32'd2570
; 
32'd150532: dataIn1 = 32'd4682
; 
32'd150533: dataIn1 = 32'd4683
; 
32'd150534: dataIn1 = 32'd4854
; 
32'd150535: dataIn1 = 32'd5981
; 
32'd150536: dataIn1 = 32'd5982
; 
32'd150537: dataIn1 = 32'd6699
; 
32'd150538: dataIn1 = 32'd1042
; 
32'd150539: dataIn1 = 32'd2546
; 
32'd150540: dataIn1 = 32'd2570
; 
32'd150541: dataIn1 = 32'd4633
; 
32'd150542: dataIn1 = 32'd4682
; 
32'd150543: dataIn1 = 32'd4683
; 
32'd150544: dataIn1 = 32'd6699
; 
32'd150545: dataIn1 = 32'd10266
; 
32'd150546: dataIn1 = 32'd10267
; 
32'd150547: dataIn1 = 32'd2572
; 
32'd150548: dataIn1 = 32'd2573
; 
32'd150549: dataIn1 = 32'd4684
; 
32'd150550: dataIn1 = 32'd4685
; 
32'd150551: dataIn1 = 32'd4686
; 
32'd150552: dataIn1 = 32'd4687
; 
32'd150553: dataIn1 = 32'd4688
; 
32'd150554: dataIn1 = 32'd9602
; 
32'd150555: dataIn1 = 32'd2571
; 
32'd150556: dataIn1 = 32'd2573
; 
32'd150557: dataIn1 = 32'd4684
; 
32'd150558: dataIn1 = 32'd4685
; 
32'd150559: dataIn1 = 32'd4686
; 
32'd150560: dataIn1 = 32'd4689
; 
32'd150561: dataIn1 = 32'd4690
; 
32'd150562: dataIn1 = 32'd2571
; 
32'd150563: dataIn1 = 32'd2572
; 
32'd150564: dataIn1 = 32'd4684
; 
32'd150565: dataIn1 = 32'd4685
; 
32'd150566: dataIn1 = 32'd4686
; 
32'd150567: dataIn1 = 32'd4691
; 
32'd150568: dataIn1 = 32'd4692
; 
32'd150569: dataIn1 = 32'd2573
; 
32'd150570: dataIn1 = 32'd4684
; 
32'd150571: dataIn1 = 32'd4687
; 
32'd150572: dataIn1 = 32'd9602
; 
32'd150573: dataIn1 = 32'd9604
; 
32'd150574: dataIn1 = 32'd9617
; 
32'd150575: dataIn1 = 32'd9619
; 
32'd150576: dataIn1 = 32'd2572
; 
32'd150577: dataIn1 = 32'd4684
; 
32'd150578: dataIn1 = 32'd4688
; 
32'd150579: dataIn1 = 32'd9602
; 
32'd150580: dataIn1 = 32'd9603
; 
32'd150581: dataIn1 = 32'd9629
; 
32'd150582: dataIn1 = 32'd9630
; 
32'd150583: dataIn1 = 32'd1078
; 
32'd150584: dataIn1 = 32'd2573
; 
32'd150585: dataIn1 = 32'd4685
; 
32'd150586: dataIn1 = 32'd4689
; 
32'd150587: dataIn1 = 32'd4690
; 
32'd150588: dataIn1 = 32'd4890
; 
32'd150589: dataIn1 = 32'd4894
; 
32'd150590: dataIn1 = 32'd1078
; 
32'd150591: dataIn1 = 32'd2571
; 
32'd150592: dataIn1 = 32'd3456
; 
32'd150593: dataIn1 = 32'd4685
; 
32'd150594: dataIn1 = 32'd4689
; 
32'd150595: dataIn1 = 32'd4690
; 
32'd150596: dataIn1 = 32'd1079
; 
32'd150597: dataIn1 = 32'd2572
; 
32'd150598: dataIn1 = 32'd4686
; 
32'd150599: dataIn1 = 32'd4691
; 
32'd150600: dataIn1 = 32'd4692
; 
32'd150601: dataIn1 = 32'd4911
; 
32'd150602: dataIn1 = 32'd4914
; 
32'd150603: dataIn1 = 32'd1079
; 
32'd150604: dataIn1 = 32'd2571
; 
32'd150605: dataIn1 = 32'd3466
; 
32'd150606: dataIn1 = 32'd4686
; 
32'd150607: dataIn1 = 32'd4691
; 
32'd150608: dataIn1 = 32'd4692
; 
32'd150609: dataIn1 = 32'd2575
; 
32'd150610: dataIn1 = 32'd2576
; 
32'd150611: dataIn1 = 32'd4693
; 
32'd150612: dataIn1 = 32'd4694
; 
32'd150613: dataIn1 = 32'd4695
; 
32'd150614: dataIn1 = 32'd4696
; 
32'd150615: dataIn1 = 32'd4697
; 
32'd150616: dataIn1 = 32'd2574
; 
32'd150617: dataIn1 = 32'd2576
; 
32'd150618: dataIn1 = 32'd4693
; 
32'd150619: dataIn1 = 32'd4694
; 
32'd150620: dataIn1 = 32'd4695
; 
32'd150621: dataIn1 = 32'd4698
; 
32'd150622: dataIn1 = 32'd4699
; 
32'd150623: dataIn1 = 32'd9606
; 
32'd150624: dataIn1 = 32'd2574
; 
32'd150625: dataIn1 = 32'd2575
; 
32'd150626: dataIn1 = 32'd4693
; 
32'd150627: dataIn1 = 32'd4694
; 
32'd150628: dataIn1 = 32'd4695
; 
32'd150629: dataIn1 = 32'd4700
; 
32'd150630: dataIn1 = 32'd4701
; 
32'd150631: dataIn1 = 32'd1080
; 
32'd150632: dataIn1 = 32'd2576
; 
32'd150633: dataIn1 = 32'd4693
; 
32'd150634: dataIn1 = 32'd4696
; 
32'd150635: dataIn1 = 32'd4697
; 
32'd150636: dataIn1 = 32'd4906
; 
32'd150637: dataIn1 = 32'd4917
; 
32'd150638: dataIn1 = 32'd1080
; 
32'd150639: dataIn1 = 32'd2575
; 
32'd150640: dataIn1 = 32'd3481
; 
32'd150641: dataIn1 = 32'd4693
; 
32'd150642: dataIn1 = 32'd4696
; 
32'd150643: dataIn1 = 32'd4697
; 
32'd150644: dataIn1 = 32'd2576
; 
32'd150645: dataIn1 = 32'd4694
; 
32'd150646: dataIn1 = 32'd4698
; 
32'd150647: dataIn1 = 32'd9606
; 
32'd150648: dataIn1 = 32'd9607
; 
32'd150649: dataIn1 = 32'd9642
; 
32'd150650: dataIn1 = 32'd9643
; 
32'd150651: dataIn1 = 32'd2574
; 
32'd150652: dataIn1 = 32'd4694
; 
32'd150653: dataIn1 = 32'd4699
; 
32'd150654: dataIn1 = 32'd9605
; 
32'd150655: dataIn1 = 32'd9606
; 
32'd150656: dataIn1 = 32'd9660
; 
32'd150657: dataIn1 = 32'd9661
; 
32'd150658: dataIn1 = 32'd1081
; 
32'd150659: dataIn1 = 32'd2575
; 
32'd150660: dataIn1 = 32'd3485
; 
32'd150661: dataIn1 = 32'd4695
; 
32'd150662: dataIn1 = 32'd4700
; 
32'd150663: dataIn1 = 32'd4701
; 
32'd150664: dataIn1 = 32'd1081
; 
32'd150665: dataIn1 = 32'd2574
; 
32'd150666: dataIn1 = 32'd4695
; 
32'd150667: dataIn1 = 32'd4700
; 
32'd150668: dataIn1 = 32'd4701
; 
32'd150669: dataIn1 = 32'd4926
; 
32'd150670: dataIn1 = 32'd4936
; 
32'd150671: dataIn1 = 32'd2578
; 
32'd150672: dataIn1 = 32'd2579
; 
32'd150673: dataIn1 = 32'd4702
; 
32'd150674: dataIn1 = 32'd4703
; 
32'd150675: dataIn1 = 32'd4704
; 
32'd150676: dataIn1 = 32'd4705
; 
32'd150677: dataIn1 = 32'd4706
; 
32'd150678: dataIn1 = 32'd9608
; 
32'd150679: dataIn1 = 32'd2577
; 
32'd150680: dataIn1 = 32'd2579
; 
32'd150681: dataIn1 = 32'd4702
; 
32'd150682: dataIn1 = 32'd4703
; 
32'd150683: dataIn1 = 32'd4704
; 
32'd150684: dataIn1 = 32'd4707
; 
32'd150685: dataIn1 = 32'd4708
; 
32'd150686: dataIn1 = 32'd2577
; 
32'd150687: dataIn1 = 32'd2578
; 
32'd150688: dataIn1 = 32'd4702
; 
32'd150689: dataIn1 = 32'd4703
; 
32'd150690: dataIn1 = 32'd4704
; 
32'd150691: dataIn1 = 32'd4709
; 
32'd150692: dataIn1 = 32'd4710
; 
32'd150693: dataIn1 = 32'd2579
; 
32'd150694: dataIn1 = 32'd4702
; 
32'd150695: dataIn1 = 32'd4705
; 
32'd150696: dataIn1 = 32'd9608
; 
32'd150697: dataIn1 = 32'd9610
; 
32'd150698: dataIn1 = 32'd9650
; 
32'd150699: dataIn1 = 32'd9652
; 
32'd150700: dataIn1 = 32'd2578
; 
32'd150701: dataIn1 = 32'd4702
; 
32'd150702: dataIn1 = 32'd4706
; 
32'd150703: dataIn1 = 32'd9608
; 
32'd150704: dataIn1 = 32'd9609
; 
32'd150705: dataIn1 = 32'd9665
; 
32'd150706: dataIn1 = 32'd9666
; 
32'd150707: dataIn1 = 32'd1082
; 
32'd150708: dataIn1 = 32'd2579
; 
32'd150709: dataIn1 = 32'd4703
; 
32'd150710: dataIn1 = 32'd4707
; 
32'd150711: dataIn1 = 32'd4708
; 
32'd150712: dataIn1 = 32'd4928
; 
32'd150713: dataIn1 = 32'd4932
; 
32'd150714: dataIn1 = 32'd1082
; 
32'd150715: dataIn1 = 32'd2577
; 
32'd150716: dataIn1 = 32'd3497
; 
32'd150717: dataIn1 = 32'd4703
; 
32'd150718: dataIn1 = 32'd4707
; 
32'd150719: dataIn1 = 32'd4708
; 
32'd150720: dataIn1 = 32'd1083
; 
32'd150721: dataIn1 = 32'd2578
; 
32'd150722: dataIn1 = 32'd4704
; 
32'd150723: dataIn1 = 32'd4709
; 
32'd150724: dataIn1 = 32'd4710
; 
32'd150725: dataIn1 = 32'd4949
; 
32'd150726: dataIn1 = 32'd4952
; 
32'd150727: dataIn1 = 32'd1083
; 
32'd150728: dataIn1 = 32'd2577
; 
32'd150729: dataIn1 = 32'd3500
; 
32'd150730: dataIn1 = 32'd4704
; 
32'd150731: dataIn1 = 32'd4709
; 
32'd150732: dataIn1 = 32'd4710
; 
32'd150733: dataIn1 = 32'd2581
; 
32'd150734: dataIn1 = 32'd2582
; 
32'd150735: dataIn1 = 32'd4711
; 
32'd150736: dataIn1 = 32'd4712
; 
32'd150737: dataIn1 = 32'd4713
; 
32'd150738: dataIn1 = 32'd4714
; 
32'd150739: dataIn1 = 32'd4715
; 
32'd150740: dataIn1 = 32'd2580
; 
32'd150741: dataIn1 = 32'd2582
; 
32'd150742: dataIn1 = 32'd4711
; 
32'd150743: dataIn1 = 32'd4712
; 
32'd150744: dataIn1 = 32'd4713
; 
32'd150745: dataIn1 = 32'd4716
; 
32'd150746: dataIn1 = 32'd4717
; 
32'd150747: dataIn1 = 32'd2580
; 
32'd150748: dataIn1 = 32'd2581
; 
32'd150749: dataIn1 = 32'd4711
; 
32'd150750: dataIn1 = 32'd4712
; 
32'd150751: dataIn1 = 32'd4713
; 
32'd150752: dataIn1 = 32'd4718
; 
32'd150753: dataIn1 = 32'd4719
; 
32'd150754: dataIn1 = 32'd1084
; 
32'd150755: dataIn1 = 32'd2582
; 
32'd150756: dataIn1 = 32'd4711
; 
32'd150757: dataIn1 = 32'd4714
; 
32'd150758: dataIn1 = 32'd4715
; 
32'd150759: dataIn1 = 32'd4944
; 
32'd150760: dataIn1 = 32'd4955
; 
32'd150761: dataIn1 = 32'd1084
; 
32'd150762: dataIn1 = 32'd2581
; 
32'd150763: dataIn1 = 32'd3507
; 
32'd150764: dataIn1 = 32'd4711
; 
32'd150765: dataIn1 = 32'd4714
; 
32'd150766: dataIn1 = 32'd4715
; 
32'd150767: dataIn1 = 32'd8
; 
32'd150768: dataIn1 = 32'd2582
; 
32'd150769: dataIn1 = 32'd4712
; 
32'd150770: dataIn1 = 32'd4716
; 
32'd150771: dataIn1 = 32'd4717
; 
32'd150772: dataIn1 = 32'd4957
; 
32'd150773: dataIn1 = 32'd4959
; 
32'd150774: dataIn1 = 32'd7859
; 
32'd150775: dataIn1 = 32'd8
; 
32'd150776: dataIn1 = 32'd2580
; 
32'd150777: dataIn1 = 32'd4712
; 
32'd150778: dataIn1 = 32'd4716
; 
32'd150779: dataIn1 = 32'd4717
; 
32'd150780: dataIn1 = 32'd4975
; 
32'd150781: dataIn1 = 32'd4977
; 
32'd150782: dataIn1 = 32'd7965
; 
32'd150783: dataIn1 = 32'd1085
; 
32'd150784: dataIn1 = 32'd2581
; 
32'd150785: dataIn1 = 32'd3509
; 
32'd150786: dataIn1 = 32'd4713
; 
32'd150787: dataIn1 = 32'd4718
; 
32'd150788: dataIn1 = 32'd4719
; 
32'd150789: dataIn1 = 32'd1085
; 
32'd150790: dataIn1 = 32'd2580
; 
32'd150791: dataIn1 = 32'd4713
; 
32'd150792: dataIn1 = 32'd4718
; 
32'd150793: dataIn1 = 32'd4719
; 
32'd150794: dataIn1 = 32'd4964
; 
32'd150795: dataIn1 = 32'd4974
; 
32'd150796: dataIn1 = 32'd2584
; 
32'd150797: dataIn1 = 32'd2585
; 
32'd150798: dataIn1 = 32'd4720
; 
32'd150799: dataIn1 = 32'd4721
; 
32'd150800: dataIn1 = 32'd4722
; 
32'd150801: dataIn1 = 32'd4723
; 
32'd150802: dataIn1 = 32'd4724
; 
32'd150803: dataIn1 = 32'd2583
; 
32'd150804: dataIn1 = 32'd2585
; 
32'd150805: dataIn1 = 32'd4720
; 
32'd150806: dataIn1 = 32'd4721
; 
32'd150807: dataIn1 = 32'd4722
; 
32'd150808: dataIn1 = 32'd4725
; 
32'd150809: dataIn1 = 32'd4726
; 
32'd150810: dataIn1 = 32'd2583
; 
32'd150811: dataIn1 = 32'd2584
; 
32'd150812: dataIn1 = 32'd4720
; 
32'd150813: dataIn1 = 32'd4721
; 
32'd150814: dataIn1 = 32'd4722
; 
32'd150815: dataIn1 = 32'd4727
; 
32'd150816: dataIn1 = 32'd4728
; 
32'd150817: dataIn1 = 32'd139
; 
32'd150818: dataIn1 = 32'd2585
; 
32'd150819: dataIn1 = 32'd4720
; 
32'd150820: dataIn1 = 32'd4723
; 
32'd150821: dataIn1 = 32'd4724
; 
32'd150822: dataIn1 = 32'd4969
; 
32'd150823: dataIn1 = 32'd4972
; 
32'd150824: dataIn1 = 32'd7995
; 
32'd150825: dataIn1 = 32'd139
; 
32'd150826: dataIn1 = 32'd2584
; 
32'd150827: dataIn1 = 32'd4720
; 
32'd150828: dataIn1 = 32'd4723
; 
32'd150829: dataIn1 = 32'd4724
; 
32'd150830: dataIn1 = 32'd4988
; 
32'd150831: dataIn1 = 32'd4991
; 
32'd150832: dataIn1 = 32'd8082
; 
32'd150833: dataIn1 = 32'd1086
; 
32'd150834: dataIn1 = 32'd2585
; 
32'd150835: dataIn1 = 32'd4721
; 
32'd150836: dataIn1 = 32'd4725
; 
32'd150837: dataIn1 = 32'd4726
; 
32'd150838: dataIn1 = 32'd4966
; 
32'd150839: dataIn1 = 32'd4970
; 
32'd150840: dataIn1 = 32'd1086
; 
32'd150841: dataIn1 = 32'd2583
; 
32'd150842: dataIn1 = 32'd3515
; 
32'd150843: dataIn1 = 32'd4721
; 
32'd150844: dataIn1 = 32'd4725
; 
32'd150845: dataIn1 = 32'd4726
; 
32'd150846: dataIn1 = 32'd1087
; 
32'd150847: dataIn1 = 32'd2584
; 
32'd150848: dataIn1 = 32'd4722
; 
32'd150849: dataIn1 = 32'd4727
; 
32'd150850: dataIn1 = 32'd4728
; 
32'd150851: dataIn1 = 32'd4987
; 
32'd150852: dataIn1 = 32'd4990
; 
32'd150853: dataIn1 = 32'd1087
; 
32'd150854: dataIn1 = 32'd2583
; 
32'd150855: dataIn1 = 32'd3517
; 
32'd150856: dataIn1 = 32'd4722
; 
32'd150857: dataIn1 = 32'd4727
; 
32'd150858: dataIn1 = 32'd4728
; 
32'd150859: dataIn1 = 32'd2587
; 
32'd150860: dataIn1 = 32'd2588
; 
32'd150861: dataIn1 = 32'd4729
; 
32'd150862: dataIn1 = 32'd4730
; 
32'd150863: dataIn1 = 32'd4731
; 
32'd150864: dataIn1 = 32'd4732
; 
32'd150865: dataIn1 = 32'd4733
; 
32'd150866: dataIn1 = 32'd2586
; 
32'd150867: dataIn1 = 32'd2588
; 
32'd150868: dataIn1 = 32'd4729
; 
32'd150869: dataIn1 = 32'd4730
; 
32'd150870: dataIn1 = 32'd4731
; 
32'd150871: dataIn1 = 32'd4734
; 
32'd150872: dataIn1 = 32'd4735
; 
32'd150873: dataIn1 = 32'd2586
; 
32'd150874: dataIn1 = 32'd2587
; 
32'd150875: dataIn1 = 32'd4729
; 
32'd150876: dataIn1 = 32'd4730
; 
32'd150877: dataIn1 = 32'd4731
; 
32'd150878: dataIn1 = 32'd4736
; 
32'd150879: dataIn1 = 32'd4737
; 
32'd150880: dataIn1 = 32'd1088
; 
32'd150881: dataIn1 = 32'd2588
; 
32'd150882: dataIn1 = 32'd4729
; 
32'd150883: dataIn1 = 32'd4732
; 
32'd150884: dataIn1 = 32'd4733
; 
32'd150885: dataIn1 = 32'd4982
; 
32'd150886: dataIn1 = 32'd4993
; 
32'd150887: dataIn1 = 32'd1088
; 
32'd150888: dataIn1 = 32'd2587
; 
32'd150889: dataIn1 = 32'd3523
; 
32'd150890: dataIn1 = 32'd4729
; 
32'd150891: dataIn1 = 32'd4732
; 
32'd150892: dataIn1 = 32'd4733
; 
32'd150893: dataIn1 = 32'd9
; 
32'd150894: dataIn1 = 32'd2588
; 
32'd150895: dataIn1 = 32'd4730
; 
32'd150896: dataIn1 = 32'd4734
; 
32'd150897: dataIn1 = 32'd4735
; 
32'd150898: dataIn1 = 32'd4995
; 
32'd150899: dataIn1 = 32'd4997
; 
32'd150900: dataIn1 = 32'd8112
; 
32'd150901: dataIn1 = 32'd9
; 
32'd150902: dataIn1 = 32'd2586
; 
32'd150903: dataIn1 = 32'd4730
; 
32'd150904: dataIn1 = 32'd4734
; 
32'd150905: dataIn1 = 32'd4735
; 
32'd150906: dataIn1 = 32'd5013
; 
32'd150907: dataIn1 = 32'd5015
; 
32'd150908: dataIn1 = 32'd8218
; 
32'd150909: dataIn1 = 32'd1089
; 
32'd150910: dataIn1 = 32'd2587
; 
32'd150911: dataIn1 = 32'd3525
; 
32'd150912: dataIn1 = 32'd4731
; 
32'd150913: dataIn1 = 32'd4736
; 
32'd150914: dataIn1 = 32'd4737
; 
32'd150915: dataIn1 = 32'd1089
; 
32'd150916: dataIn1 = 32'd2586
; 
32'd150917: dataIn1 = 32'd4731
; 
32'd150918: dataIn1 = 32'd4736
; 
32'd150919: dataIn1 = 32'd4737
; 
32'd150920: dataIn1 = 32'd5002
; 
32'd150921: dataIn1 = 32'd5012
; 
32'd150922: dataIn1 = 32'd2590
; 
32'd150923: dataIn1 = 32'd2591
; 
32'd150924: dataIn1 = 32'd4738
; 
32'd150925: dataIn1 = 32'd4739
; 
32'd150926: dataIn1 = 32'd4740
; 
32'd150927: dataIn1 = 32'd4741
; 
32'd150928: dataIn1 = 32'd4742
; 
32'd150929: dataIn1 = 32'd2589
; 
32'd150930: dataIn1 = 32'd2591
; 
32'd150931: dataIn1 = 32'd4738
; 
32'd150932: dataIn1 = 32'd4739
; 
32'd150933: dataIn1 = 32'd4740
; 
32'd150934: dataIn1 = 32'd4743
; 
32'd150935: dataIn1 = 32'd4744
; 
32'd150936: dataIn1 = 32'd2589
; 
32'd150937: dataIn1 = 32'd2590
; 
32'd150938: dataIn1 = 32'd4738
; 
32'd150939: dataIn1 = 32'd4739
; 
32'd150940: dataIn1 = 32'd4740
; 
32'd150941: dataIn1 = 32'd4745
; 
32'd150942: dataIn1 = 32'd4746
; 
32'd150943: dataIn1 = 32'd142
; 
32'd150944: dataIn1 = 32'd2591
; 
32'd150945: dataIn1 = 32'd4738
; 
32'd150946: dataIn1 = 32'd4741
; 
32'd150947: dataIn1 = 32'd4742
; 
32'd150948: dataIn1 = 32'd5007
; 
32'd150949: dataIn1 = 32'd5010
; 
32'd150950: dataIn1 = 32'd8248
; 
32'd150951: dataIn1 = 32'd142
; 
32'd150952: dataIn1 = 32'd2590
; 
32'd150953: dataIn1 = 32'd4738
; 
32'd150954: dataIn1 = 32'd4741
; 
32'd150955: dataIn1 = 32'd4742
; 
32'd150956: dataIn1 = 32'd5026
; 
32'd150957: dataIn1 = 32'd5029
; 
32'd150958: dataIn1 = 32'd8334
; 
32'd150959: dataIn1 = 32'd1090
; 
32'd150960: dataIn1 = 32'd2591
; 
32'd150961: dataIn1 = 32'd4739
; 
32'd150962: dataIn1 = 32'd4743
; 
32'd150963: dataIn1 = 32'd4744
; 
32'd150964: dataIn1 = 32'd5004
; 
32'd150965: dataIn1 = 32'd5008
; 
32'd150966: dataIn1 = 32'd1090
; 
32'd150967: dataIn1 = 32'd2589
; 
32'd150968: dataIn1 = 32'd3531
; 
32'd150969: dataIn1 = 32'd4739
; 
32'd150970: dataIn1 = 32'd4743
; 
32'd150971: dataIn1 = 32'd4744
; 
32'd150972: dataIn1 = 32'd1091
; 
32'd150973: dataIn1 = 32'd2590
; 
32'd150974: dataIn1 = 32'd4740
; 
32'd150975: dataIn1 = 32'd4745
; 
32'd150976: dataIn1 = 32'd4746
; 
32'd150977: dataIn1 = 32'd5025
; 
32'd150978: dataIn1 = 32'd5028
; 
32'd150979: dataIn1 = 32'd1091
; 
32'd150980: dataIn1 = 32'd2589
; 
32'd150981: dataIn1 = 32'd3533
; 
32'd150982: dataIn1 = 32'd4740
; 
32'd150983: dataIn1 = 32'd4745
; 
32'd150984: dataIn1 = 32'd4746
; 
32'd150985: dataIn1 = 32'd2593
; 
32'd150986: dataIn1 = 32'd2594
; 
32'd150987: dataIn1 = 32'd4747
; 
32'd150988: dataIn1 = 32'd4748
; 
32'd150989: dataIn1 = 32'd4749
; 
32'd150990: dataIn1 = 32'd4750
; 
32'd150991: dataIn1 = 32'd4751
; 
32'd150992: dataIn1 = 32'd2592
; 
32'd150993: dataIn1 = 32'd2594
; 
32'd150994: dataIn1 = 32'd4747
; 
32'd150995: dataIn1 = 32'd4748
; 
32'd150996: dataIn1 = 32'd4749
; 
32'd150997: dataIn1 = 32'd4752
; 
32'd150998: dataIn1 = 32'd4753
; 
32'd150999: dataIn1 = 32'd2592
; 
32'd151000: dataIn1 = 32'd2593
; 
32'd151001: dataIn1 = 32'd4747
; 
32'd151002: dataIn1 = 32'd4748
; 
32'd151003: dataIn1 = 32'd4749
; 
32'd151004: dataIn1 = 32'd4754
; 
32'd151005: dataIn1 = 32'd4755
; 
32'd151006: dataIn1 = 32'd1092
; 
32'd151007: dataIn1 = 32'd2594
; 
32'd151008: dataIn1 = 32'd4747
; 
32'd151009: dataIn1 = 32'd4750
; 
32'd151010: dataIn1 = 32'd4751
; 
32'd151011: dataIn1 = 32'd5020
; 
32'd151012: dataIn1 = 32'd5031
; 
32'd151013: dataIn1 = 32'd1092
; 
32'd151014: dataIn1 = 32'd2593
; 
32'd151015: dataIn1 = 32'd3539
; 
32'd151016: dataIn1 = 32'd4747
; 
32'd151017: dataIn1 = 32'd4750
; 
32'd151018: dataIn1 = 32'd4751
; 
32'd151019: dataIn1 = 32'd10
; 
32'd151020: dataIn1 = 32'd2594
; 
32'd151021: dataIn1 = 32'd4748
; 
32'd151022: dataIn1 = 32'd4752
; 
32'd151023: dataIn1 = 32'd4753
; 
32'd151024: dataIn1 = 32'd5033
; 
32'd151025: dataIn1 = 32'd5035
; 
32'd151026: dataIn1 = 32'd8364
; 
32'd151027: dataIn1 = 32'd10
; 
32'd151028: dataIn1 = 32'd2592
; 
32'd151029: dataIn1 = 32'd4748
; 
32'd151030: dataIn1 = 32'd4752
; 
32'd151031: dataIn1 = 32'd4753
; 
32'd151032: dataIn1 = 32'd5051
; 
32'd151033: dataIn1 = 32'd5053
; 
32'd151034: dataIn1 = 32'd8470
; 
32'd151035: dataIn1 = 32'd1093
; 
32'd151036: dataIn1 = 32'd2593
; 
32'd151037: dataIn1 = 32'd3541
; 
32'd151038: dataIn1 = 32'd4749
; 
32'd151039: dataIn1 = 32'd4754
; 
32'd151040: dataIn1 = 32'd4755
; 
32'd151041: dataIn1 = 32'd1093
; 
32'd151042: dataIn1 = 32'd2592
; 
32'd151043: dataIn1 = 32'd4749
; 
32'd151044: dataIn1 = 32'd4754
; 
32'd151045: dataIn1 = 32'd4755
; 
32'd151046: dataIn1 = 32'd5040
; 
32'd151047: dataIn1 = 32'd5050
; 
32'd151048: dataIn1 = 32'd2596
; 
32'd151049: dataIn1 = 32'd2597
; 
32'd151050: dataIn1 = 32'd4756
; 
32'd151051: dataIn1 = 32'd4757
; 
32'd151052: dataIn1 = 32'd4758
; 
32'd151053: dataIn1 = 32'd4759
; 
32'd151054: dataIn1 = 32'd4760
; 
32'd151055: dataIn1 = 32'd2595
; 
32'd151056: dataIn1 = 32'd2597
; 
32'd151057: dataIn1 = 32'd4756
; 
32'd151058: dataIn1 = 32'd4757
; 
32'd151059: dataIn1 = 32'd4758
; 
32'd151060: dataIn1 = 32'd4761
; 
32'd151061: dataIn1 = 32'd4762
; 
32'd151062: dataIn1 = 32'd2595
; 
32'd151063: dataIn1 = 32'd2596
; 
32'd151064: dataIn1 = 32'd4756
; 
32'd151065: dataIn1 = 32'd4757
; 
32'd151066: dataIn1 = 32'd4758
; 
32'd151067: dataIn1 = 32'd4763
; 
32'd151068: dataIn1 = 32'd4764
; 
32'd151069: dataIn1 = 32'd145
; 
32'd151070: dataIn1 = 32'd2597
; 
32'd151071: dataIn1 = 32'd4756
; 
32'd151072: dataIn1 = 32'd4759
; 
32'd151073: dataIn1 = 32'd4760
; 
32'd151074: dataIn1 = 32'd5045
; 
32'd151075: dataIn1 = 32'd5048
; 
32'd151076: dataIn1 = 32'd8500
; 
32'd151077: dataIn1 = 32'd145
; 
32'd151078: dataIn1 = 32'd2596
; 
32'd151079: dataIn1 = 32'd4756
; 
32'd151080: dataIn1 = 32'd4759
; 
32'd151081: dataIn1 = 32'd4760
; 
32'd151082: dataIn1 = 32'd5064
; 
32'd151083: dataIn1 = 32'd5067
; 
32'd151084: dataIn1 = 32'd8587
; 
32'd151085: dataIn1 = 32'd1094
; 
32'd151086: dataIn1 = 32'd2597
; 
32'd151087: dataIn1 = 32'd4757
; 
32'd151088: dataIn1 = 32'd4761
; 
32'd151089: dataIn1 = 32'd4762
; 
32'd151090: dataIn1 = 32'd5042
; 
32'd151091: dataIn1 = 32'd5046
; 
32'd151092: dataIn1 = 32'd1094
; 
32'd151093: dataIn1 = 32'd2595
; 
32'd151094: dataIn1 = 32'd3547
; 
32'd151095: dataIn1 = 32'd4757
; 
32'd151096: dataIn1 = 32'd4761
; 
32'd151097: dataIn1 = 32'd4762
; 
32'd151098: dataIn1 = 32'd1095
; 
32'd151099: dataIn1 = 32'd2596
; 
32'd151100: dataIn1 = 32'd4758
; 
32'd151101: dataIn1 = 32'd4763
; 
32'd151102: dataIn1 = 32'd4764
; 
32'd151103: dataIn1 = 32'd5063
; 
32'd151104: dataIn1 = 32'd5066
; 
32'd151105: dataIn1 = 32'd1095
; 
32'd151106: dataIn1 = 32'd2595
; 
32'd151107: dataIn1 = 32'd3549
; 
32'd151108: dataIn1 = 32'd4758
; 
32'd151109: dataIn1 = 32'd4763
; 
32'd151110: dataIn1 = 32'd4764
; 
32'd151111: dataIn1 = 32'd2599
; 
32'd151112: dataIn1 = 32'd2600
; 
32'd151113: dataIn1 = 32'd4765
; 
32'd151114: dataIn1 = 32'd4766
; 
32'd151115: dataIn1 = 32'd4767
; 
32'd151116: dataIn1 = 32'd4768
; 
32'd151117: dataIn1 = 32'd4769
; 
32'd151118: dataIn1 = 32'd2598
; 
32'd151119: dataIn1 = 32'd2600
; 
32'd151120: dataIn1 = 32'd4765
; 
32'd151121: dataIn1 = 32'd4766
; 
32'd151122: dataIn1 = 32'd4767
; 
32'd151123: dataIn1 = 32'd4770
; 
32'd151124: dataIn1 = 32'd4771
; 
32'd151125: dataIn1 = 32'd2598
; 
32'd151126: dataIn1 = 32'd2599
; 
32'd151127: dataIn1 = 32'd4765
; 
32'd151128: dataIn1 = 32'd4766
; 
32'd151129: dataIn1 = 32'd4767
; 
32'd151130: dataIn1 = 32'd4772
; 
32'd151131: dataIn1 = 32'd4773
; 
32'd151132: dataIn1 = 32'd1096
; 
32'd151133: dataIn1 = 32'd2600
; 
32'd151134: dataIn1 = 32'd4765
; 
32'd151135: dataIn1 = 32'd4768
; 
32'd151136: dataIn1 = 32'd4769
; 
32'd151137: dataIn1 = 32'd5058
; 
32'd151138: dataIn1 = 32'd5069
; 
32'd151139: dataIn1 = 32'd1096
; 
32'd151140: dataIn1 = 32'd2599
; 
32'd151141: dataIn1 = 32'd3555
; 
32'd151142: dataIn1 = 32'd4765
; 
32'd151143: dataIn1 = 32'd4768
; 
32'd151144: dataIn1 = 32'd4769
; 
32'd151145: dataIn1 = 32'd11
; 
32'd151146: dataIn1 = 32'd2600
; 
32'd151147: dataIn1 = 32'd4766
; 
32'd151148: dataIn1 = 32'd4770
; 
32'd151149: dataIn1 = 32'd4771
; 
32'd151150: dataIn1 = 32'd5071
; 
32'd151151: dataIn1 = 32'd5073
; 
32'd151152: dataIn1 = 32'd8617
; 
32'd151153: dataIn1 = 32'd11
; 
32'd151154: dataIn1 = 32'd2598
; 
32'd151155: dataIn1 = 32'd4766
; 
32'd151156: dataIn1 = 32'd4770
; 
32'd151157: dataIn1 = 32'd4771
; 
32'd151158: dataIn1 = 32'd5089
; 
32'd151159: dataIn1 = 32'd5091
; 
32'd151160: dataIn1 = 32'd8723
; 
32'd151161: dataIn1 = 32'd1097
; 
32'd151162: dataIn1 = 32'd2599
; 
32'd151163: dataIn1 = 32'd3557
; 
32'd151164: dataIn1 = 32'd4767
; 
32'd151165: dataIn1 = 32'd4772
; 
32'd151166: dataIn1 = 32'd4773
; 
32'd151167: dataIn1 = 32'd1097
; 
32'd151168: dataIn1 = 32'd2598
; 
32'd151169: dataIn1 = 32'd4767
; 
32'd151170: dataIn1 = 32'd4772
; 
32'd151171: dataIn1 = 32'd4773
; 
32'd151172: dataIn1 = 32'd5078
; 
32'd151173: dataIn1 = 32'd5088
; 
32'd151174: dataIn1 = 32'd2602
; 
32'd151175: dataIn1 = 32'd2603
; 
32'd151176: dataIn1 = 32'd4774
; 
32'd151177: dataIn1 = 32'd4775
; 
32'd151178: dataIn1 = 32'd4776
; 
32'd151179: dataIn1 = 32'd4777
; 
32'd151180: dataIn1 = 32'd4778
; 
32'd151181: dataIn1 = 32'd2601
; 
32'd151182: dataIn1 = 32'd2603
; 
32'd151183: dataIn1 = 32'd4774
; 
32'd151184: dataIn1 = 32'd4775
; 
32'd151185: dataIn1 = 32'd4776
; 
32'd151186: dataIn1 = 32'd4779
; 
32'd151187: dataIn1 = 32'd4780
; 
32'd151188: dataIn1 = 32'd2601
; 
32'd151189: dataIn1 = 32'd2602
; 
32'd151190: dataIn1 = 32'd4774
; 
32'd151191: dataIn1 = 32'd4775
; 
32'd151192: dataIn1 = 32'd4776
; 
32'd151193: dataIn1 = 32'd4781
; 
32'd151194: dataIn1 = 32'd4782
; 
32'd151195: dataIn1 = 32'd148
; 
32'd151196: dataIn1 = 32'd2603
; 
32'd151197: dataIn1 = 32'd4774
; 
32'd151198: dataIn1 = 32'd4777
; 
32'd151199: dataIn1 = 32'd4778
; 
32'd151200: dataIn1 = 32'd5083
; 
32'd151201: dataIn1 = 32'd5086
; 
32'd151202: dataIn1 = 32'd8753
; 
32'd151203: dataIn1 = 32'd148
; 
32'd151204: dataIn1 = 32'd2602
; 
32'd151205: dataIn1 = 32'd4774
; 
32'd151206: dataIn1 = 32'd4777
; 
32'd151207: dataIn1 = 32'd4778
; 
32'd151208: dataIn1 = 32'd5102
; 
32'd151209: dataIn1 = 32'd5105
; 
32'd151210: dataIn1 = 32'd8839
; 
32'd151211: dataIn1 = 32'd1098
; 
32'd151212: dataIn1 = 32'd2603
; 
32'd151213: dataIn1 = 32'd4775
; 
32'd151214: dataIn1 = 32'd4779
; 
32'd151215: dataIn1 = 32'd4780
; 
32'd151216: dataIn1 = 32'd5080
; 
32'd151217: dataIn1 = 32'd5084
; 
32'd151218: dataIn1 = 32'd1098
; 
32'd151219: dataIn1 = 32'd2601
; 
32'd151220: dataIn1 = 32'd3563
; 
32'd151221: dataIn1 = 32'd4775
; 
32'd151222: dataIn1 = 32'd4779
; 
32'd151223: dataIn1 = 32'd4780
; 
32'd151224: dataIn1 = 32'd1099
; 
32'd151225: dataIn1 = 32'd2602
; 
32'd151226: dataIn1 = 32'd4776
; 
32'd151227: dataIn1 = 32'd4781
; 
32'd151228: dataIn1 = 32'd4782
; 
32'd151229: dataIn1 = 32'd5101
; 
32'd151230: dataIn1 = 32'd5104
; 
32'd151231: dataIn1 = 32'd1099
; 
32'd151232: dataIn1 = 32'd2601
; 
32'd151233: dataIn1 = 32'd3565
; 
32'd151234: dataIn1 = 32'd4776
; 
32'd151235: dataIn1 = 32'd4781
; 
32'd151236: dataIn1 = 32'd4782
; 
32'd151237: dataIn1 = 32'd2605
; 
32'd151238: dataIn1 = 32'd2606
; 
32'd151239: dataIn1 = 32'd4783
; 
32'd151240: dataIn1 = 32'd4784
; 
32'd151241: dataIn1 = 32'd4785
; 
32'd151242: dataIn1 = 32'd4786
; 
32'd151243: dataIn1 = 32'd4787
; 
32'd151244: dataIn1 = 32'd2604
; 
32'd151245: dataIn1 = 32'd2606
; 
32'd151246: dataIn1 = 32'd4783
; 
32'd151247: dataIn1 = 32'd4784
; 
32'd151248: dataIn1 = 32'd4785
; 
32'd151249: dataIn1 = 32'd4788
; 
32'd151250: dataIn1 = 32'd4789
; 
32'd151251: dataIn1 = 32'd2604
; 
32'd151252: dataIn1 = 32'd2605
; 
32'd151253: dataIn1 = 32'd4783
; 
32'd151254: dataIn1 = 32'd4784
; 
32'd151255: dataIn1 = 32'd4785
; 
32'd151256: dataIn1 = 32'd4790
; 
32'd151257: dataIn1 = 32'd4791
; 
32'd151258: dataIn1 = 32'd1100
; 
32'd151259: dataIn1 = 32'd2606
; 
32'd151260: dataIn1 = 32'd4783
; 
32'd151261: dataIn1 = 32'd4786
; 
32'd151262: dataIn1 = 32'd4787
; 
32'd151263: dataIn1 = 32'd5096
; 
32'd151264: dataIn1 = 32'd5107
; 
32'd151265: dataIn1 = 32'd1100
; 
32'd151266: dataIn1 = 32'd2605
; 
32'd151267: dataIn1 = 32'd3571
; 
32'd151268: dataIn1 = 32'd3573
; 
32'd151269: dataIn1 = 32'd4783
; 
32'd151270: dataIn1 = 32'd4786
; 
32'd151271: dataIn1 = 32'd4787
; 
32'd151272: dataIn1 = 32'd12
; 
32'd151273: dataIn1 = 32'd2606
; 
32'd151274: dataIn1 = 32'd4784
; 
32'd151275: dataIn1 = 32'd4788
; 
32'd151276: dataIn1 = 32'd4789
; 
32'd151277: dataIn1 = 32'd5109
; 
32'd151278: dataIn1 = 32'd5111
; 
32'd151279: dataIn1 = 32'd8869
; 
32'd151280: dataIn1 = 32'd12
; 
32'd151281: dataIn1 = 32'd2604
; 
32'd151282: dataIn1 = 32'd4784
; 
32'd151283: dataIn1 = 32'd4788
; 
32'd151284: dataIn1 = 32'd4789
; 
32'd151285: dataIn1 = 32'd1101
; 
32'd151286: dataIn1 = 32'd2605
; 
32'd151287: dataIn1 = 32'd3573
; 
32'd151288: dataIn1 = 32'd3575
; 
32'd151289: dataIn1 = 32'd4785
; 
32'd151290: dataIn1 = 32'd4790
; 
32'd151291: dataIn1 = 32'd4791
; 
32'd151292: dataIn1 = 32'd1101
; 
32'd151293: dataIn1 = 32'd2604
; 
32'd151294: dataIn1 = 32'd4785
; 
32'd151295: dataIn1 = 32'd4790
; 
32'd151296: dataIn1 = 32'd4791
; 
32'd151297: dataIn1 = 32'd1102
; 
32'd151298: dataIn1 = 32'd2608
; 
32'd151299: dataIn1 = 32'd4792
; 
32'd151300: dataIn1 = 32'd4793
; 
32'd151301: dataIn1 = 32'd4794
; 
32'd151302: dataIn1 = 32'd4802
; 
32'd151303: dataIn1 = 32'd4804
; 
32'd151304: dataIn1 = 32'd9696
; 
32'd151305: dataIn1 = 32'd1102
; 
32'd151306: dataIn1 = 32'd2607
; 
32'd151307: dataIn1 = 32'd4792
; 
32'd151308: dataIn1 = 32'd4793
; 
32'd151309: dataIn1 = 32'd4794
; 
32'd151310: dataIn1 = 32'd4797
; 
32'd151311: dataIn1 = 32'd4799
; 
32'd151312: dataIn1 = 32'd9709
; 
32'd151313: dataIn1 = 32'd2607
; 
32'd151314: dataIn1 = 32'd2608
; 
32'd151315: dataIn1 = 32'd2609
; 
32'd151316: dataIn1 = 32'd4792
; 
32'd151317: dataIn1 = 32'd4793
; 
32'd151318: dataIn1 = 32'd4794
; 
32'd151319: dataIn1 = 32'd2552
; 
32'd151320: dataIn1 = 32'd2610
; 
32'd151321: dataIn1 = 32'd4640
; 
32'd151322: dataIn1 = 32'd4795
; 
32'd151323: dataIn1 = 32'd4796
; 
32'd151324: dataIn1 = 32'd4797
; 
32'd151325: dataIn1 = 32'd4798
; 
32'd151326: dataIn1 = 32'd9703
; 
32'd151327: dataIn1 = 32'd1070
; 
32'd151328: dataIn1 = 32'd2552
; 
32'd151329: dataIn1 = 32'd2607
; 
32'd151330: dataIn1 = 32'd4795
; 
32'd151331: dataIn1 = 32'd4796
; 
32'd151332: dataIn1 = 32'd4797
; 
32'd151333: dataIn1 = 32'd2607
; 
32'd151334: dataIn1 = 32'd2610
; 
32'd151335: dataIn1 = 32'd4793
; 
32'd151336: dataIn1 = 32'd4795
; 
32'd151337: dataIn1 = 32'd4796
; 
32'd151338: dataIn1 = 32'd4797
; 
32'd151339: dataIn1 = 32'd4799
; 
32'd151340: dataIn1 = 32'd9708
; 
32'd151341: dataIn1 = 32'd4640
; 
32'd151342: dataIn1 = 32'd4795
; 
32'd151343: dataIn1 = 32'd4798
; 
32'd151344: dataIn1 = 32'd9700
; 
32'd151345: dataIn1 = 32'd9701
; 
32'd151346: dataIn1 = 32'd9703
; 
32'd151347: dataIn1 = 32'd9704
; 
32'd151348: dataIn1 = 32'd4793
; 
32'd151349: dataIn1 = 32'd4797
; 
32'd151350: dataIn1 = 32'd4799
; 
32'd151351: dataIn1 = 32'd9705
; 
32'd151352: dataIn1 = 32'd9707
; 
32'd151353: dataIn1 = 32'd9708
; 
32'd151354: dataIn1 = 32'd9709
; 
32'd151355: dataIn1 = 32'd1069
; 
32'd151356: dataIn1 = 32'd2547
; 
32'd151357: dataIn1 = 32'd2608
; 
32'd151358: dataIn1 = 32'd4800
; 
32'd151359: dataIn1 = 32'd4801
; 
32'd151360: dataIn1 = 32'd4802
; 
32'd151361: dataIn1 = 32'd2547
; 
32'd151362: dataIn1 = 32'd2611
; 
32'd151363: dataIn1 = 32'd4638
; 
32'd151364: dataIn1 = 32'd4800
; 
32'd151365: dataIn1 = 32'd4801
; 
32'd151366: dataIn1 = 32'd4802
; 
32'd151367: dataIn1 = 32'd4803
; 
32'd151368: dataIn1 = 32'd9691
; 
32'd151369: dataIn1 = 32'd2608
; 
32'd151370: dataIn1 = 32'd2611
; 
32'd151371: dataIn1 = 32'd4792
; 
32'd151372: dataIn1 = 32'd4800
; 
32'd151373: dataIn1 = 32'd4801
; 
32'd151374: dataIn1 = 32'd4802
; 
32'd151375: dataIn1 = 32'd4804
; 
32'd151376: dataIn1 = 32'd9695
; 
32'd151377: dataIn1 = 32'd4638
; 
32'd151378: dataIn1 = 32'd4801
; 
32'd151379: dataIn1 = 32'd4803
; 
32'd151380: dataIn1 = 32'd9686
; 
32'd151381: dataIn1 = 32'd9687
; 
32'd151382: dataIn1 = 32'd9689
; 
32'd151383: dataIn1 = 32'd9691
; 
32'd151384: dataIn1 = 32'd4792
; 
32'd151385: dataIn1 = 32'd4802
; 
32'd151386: dataIn1 = 32'd4804
; 
32'd151387: dataIn1 = 32'd9693
; 
32'd151388: dataIn1 = 32'd9694
; 
32'd151389: dataIn1 = 32'd9695
; 
32'd151390: dataIn1 = 32'd9696
; 
32'd151391: dataIn1 = 32'd1103
; 
32'd151392: dataIn1 = 32'd2614
; 
32'd151393: dataIn1 = 32'd4805
; 
32'd151394: dataIn1 = 32'd4806
; 
32'd151395: dataIn1 = 32'd4807
; 
32'd151396: dataIn1 = 32'd4814
; 
32'd151397: dataIn1 = 32'd4816
; 
32'd151398: dataIn1 = 32'd9729
; 
32'd151399: dataIn1 = 32'd2612
; 
32'd151400: dataIn1 = 32'd2613
; 
32'd151401: dataIn1 = 32'd2614
; 
32'd151402: dataIn1 = 32'd4805
; 
32'd151403: dataIn1 = 32'd4806
; 
32'd151404: dataIn1 = 32'd4807
; 
32'd151405: dataIn1 = 32'd1103
; 
32'd151406: dataIn1 = 32'd2612
; 
32'd151407: dataIn1 = 32'd4805
; 
32'd151408: dataIn1 = 32'd4806
; 
32'd151409: dataIn1 = 32'd4807
; 
32'd151410: dataIn1 = 32'd4809
; 
32'd151411: dataIn1 = 32'd4812
; 
32'd151412: dataIn1 = 32'd9719
; 
32'd151413: dataIn1 = 32'd2551
; 
32'd151414: dataIn1 = 32'd2615
; 
32'd151415: dataIn1 = 32'd4641
; 
32'd151416: dataIn1 = 32'd4808
; 
32'd151417: dataIn1 = 32'd4809
; 
32'd151418: dataIn1 = 32'd4810
; 
32'd151419: dataIn1 = 32'd4811
; 
32'd151420: dataIn1 = 32'd9725
; 
32'd151421: dataIn1 = 32'd2612
; 
32'd151422: dataIn1 = 32'd2615
; 
32'd151423: dataIn1 = 32'd4807
; 
32'd151424: dataIn1 = 32'd4808
; 
32'd151425: dataIn1 = 32'd4809
; 
32'd151426: dataIn1 = 32'd4810
; 
32'd151427: dataIn1 = 32'd4812
; 
32'd151428: dataIn1 = 32'd9720
; 
32'd151429: dataIn1 = 32'd1071
; 
32'd151430: dataIn1 = 32'd2551
; 
32'd151431: dataIn1 = 32'd2612
; 
32'd151432: dataIn1 = 32'd4808
; 
32'd151433: dataIn1 = 32'd4809
; 
32'd151434: dataIn1 = 32'd4810
; 
32'd151435: dataIn1 = 32'd4641
; 
32'd151436: dataIn1 = 32'd4808
; 
32'd151437: dataIn1 = 32'd4811
; 
32'd151438: dataIn1 = 32'd9722
; 
32'd151439: dataIn1 = 32'd9723
; 
32'd151440: dataIn1 = 32'd9724
; 
32'd151441: dataIn1 = 32'd9725
; 
32'd151442: dataIn1 = 32'd4807
; 
32'd151443: dataIn1 = 32'd4809
; 
32'd151444: dataIn1 = 32'd4812
; 
32'd151445: dataIn1 = 32'd9716
; 
32'd151446: dataIn1 = 32'd9718
; 
32'd151447: dataIn1 = 32'd9719
; 
32'd151448: dataIn1 = 32'd9720
; 
32'd151449: dataIn1 = 32'd1072
; 
32'd151450: dataIn1 = 32'd2557
; 
32'd151451: dataIn1 = 32'd2614
; 
32'd151452: dataIn1 = 32'd4813
; 
32'd151453: dataIn1 = 32'd4814
; 
32'd151454: dataIn1 = 32'd4815
; 
32'd151455: dataIn1 = 32'd2614
; 
32'd151456: dataIn1 = 32'd2616
; 
32'd151457: dataIn1 = 32'd4805
; 
32'd151458: dataIn1 = 32'd4813
; 
32'd151459: dataIn1 = 32'd4814
; 
32'd151460: dataIn1 = 32'd4815
; 
32'd151461: dataIn1 = 32'd4816
; 
32'd151462: dataIn1 = 32'd9730
; 
32'd151463: dataIn1 = 32'd2557
; 
32'd151464: dataIn1 = 32'd2616
; 
32'd151465: dataIn1 = 32'd4644
; 
32'd151466: dataIn1 = 32'd4813
; 
32'd151467: dataIn1 = 32'd4814
; 
32'd151468: dataIn1 = 32'd4815
; 
32'd151469: dataIn1 = 32'd4817
; 
32'd151470: dataIn1 = 32'd4805
; 
32'd151471: dataIn1 = 32'd4814
; 
32'd151472: dataIn1 = 32'd4816
; 
32'd151473: dataIn1 = 32'd9726
; 
32'd151474: dataIn1 = 32'd9727
; 
32'd151475: dataIn1 = 32'd9729
; 
32'd151476: dataIn1 = 32'd9730
; 
32'd151477: dataIn1 = 32'd4
; 
32'd151478: dataIn1 = 32'd2616
; 
32'd151479: dataIn1 = 32'd4644
; 
32'd151480: dataIn1 = 32'd4815
; 
32'd151481: dataIn1 = 32'd4817
; 
32'd151482: dataIn1 = 32'd6138
; 
32'd151483: dataIn1 = 32'd6140
; 
32'd151484: dataIn1 = 32'd7220
; 
32'd151485: dataIn1 = 32'd9758
; 
32'd151486: dataIn1 = 32'd2618
; 
32'd151487: dataIn1 = 32'd2619
; 
32'd151488: dataIn1 = 32'd4818
; 
32'd151489: dataIn1 = 32'd4819
; 
32'd151490: dataIn1 = 32'd4820
; 
32'd151491: dataIn1 = 32'd4821
; 
32'd151492: dataIn1 = 32'd4822
; 
32'd151493: dataIn1 = 32'd2617
; 
32'd151494: dataIn1 = 32'd2619
; 
32'd151495: dataIn1 = 32'd4818
; 
32'd151496: dataIn1 = 32'd4819
; 
32'd151497: dataIn1 = 32'd4820
; 
32'd151498: dataIn1 = 32'd4823
; 
32'd151499: dataIn1 = 32'd4824
; 
32'd151500: dataIn1 = 32'd2617
; 
32'd151501: dataIn1 = 32'd2618
; 
32'd151502: dataIn1 = 32'd4818
; 
32'd151503: dataIn1 = 32'd4819
; 
32'd151504: dataIn1 = 32'd4820
; 
32'd151505: dataIn1 = 32'd4825
; 
32'd151506: dataIn1 = 32'd4826
; 
32'd151507: dataIn1 = 32'd1073
; 
32'd151508: dataIn1 = 32'd2619
; 
32'd151509: dataIn1 = 32'd4818
; 
32'd151510: dataIn1 = 32'd4821
; 
32'd151511: dataIn1 = 32'd4822
; 
32'd151512: dataIn1 = 32'd5430
; 
32'd151513: dataIn1 = 32'd5512
; 
32'd151514: dataIn1 = 32'd1073
; 
32'd151515: dataIn1 = 32'd2618
; 
32'd151516: dataIn1 = 32'd4818
; 
32'd151517: dataIn1 = 32'd4821
; 
32'd151518: dataIn1 = 32'd4822
; 
32'd151519: dataIn1 = 32'd4832
; 
32'd151520: dataIn1 = 32'd4835
; 
32'd151521: dataIn1 = 32'd444
; 
32'd151522: dataIn1 = 32'd2619
; 
32'd151523: dataIn1 = 32'd3898
; 
32'd151524: dataIn1 = 32'd4819
; 
32'd151525: dataIn1 = 32'd4823
; 
32'd151526: dataIn1 = 32'd4824
; 
32'd151527: dataIn1 = 32'd5318
; 
32'd151528: dataIn1 = 32'd444
; 
32'd151529: dataIn1 = 32'd2617
; 
32'd151530: dataIn1 = 32'd3885
; 
32'd151531: dataIn1 = 32'd4819
; 
32'd151532: dataIn1 = 32'd4823
; 
32'd151533: dataIn1 = 32'd4824
; 
32'd151534: dataIn1 = 32'd4828
; 
32'd151535: dataIn1 = 32'd1104
; 
32'd151536: dataIn1 = 32'd2618
; 
32'd151537: dataIn1 = 32'd4820
; 
32'd151538: dataIn1 = 32'd4825
; 
32'd151539: dataIn1 = 32'd4826
; 
32'd151540: dataIn1 = 32'd4834
; 
32'd151541: dataIn1 = 32'd4837
; 
32'd151542: dataIn1 = 32'd1104
; 
32'd151543: dataIn1 = 32'd2617
; 
32'd151544: dataIn1 = 32'd4820
; 
32'd151545: dataIn1 = 32'd4825
; 
32'd151546: dataIn1 = 32'd4826
; 
32'd151547: dataIn1 = 32'd4829
; 
32'd151548: dataIn1 = 32'd4831
; 
32'd151549: dataIn1 = 32'd6971
; 
32'd151550: dataIn1 = 32'd2300
; 
32'd151551: dataIn1 = 32'd4827
; 
32'd151552: dataIn1 = 32'd4828
; 
32'd151553: dataIn1 = 32'd4829
; 
32'd151554: dataIn1 = 32'd5942
; 
32'd151555: dataIn1 = 32'd5943
; 
32'd151556: dataIn1 = 32'd5946
; 
32'd151557: dataIn1 = 32'd2300
; 
32'd151558: dataIn1 = 32'd2617
; 
32'd151559: dataIn1 = 32'd3885
; 
32'd151560: dataIn1 = 32'd4824
; 
32'd151561: dataIn1 = 32'd4827
; 
32'd151562: dataIn1 = 32'd4828
; 
32'd151563: dataIn1 = 32'd4829
; 
32'd151564: dataIn1 = 32'd2617
; 
32'd151565: dataIn1 = 32'd2620
; 
32'd151566: dataIn1 = 32'd4826
; 
32'd151567: dataIn1 = 32'd4827
; 
32'd151568: dataIn1 = 32'd4828
; 
32'd151569: dataIn1 = 32'd4829
; 
32'd151570: dataIn1 = 32'd4831
; 
32'd151571: dataIn1 = 32'd5946
; 
32'd151572: dataIn1 = 32'd6970
; 
32'd151573: dataIn1 = 32'd4830
; 
32'd151574: dataIn1 = 32'd5941
; 
32'd151575: dataIn1 = 32'd5942
; 
32'd151576: dataIn1 = 32'd5944
; 
32'd151577: dataIn1 = 32'd5945
; 
32'd151578: dataIn1 = 32'd6964
; 
32'd151579: dataIn1 = 32'd6965
; 
32'd151580: dataIn1 = 32'd4826
; 
32'd151581: dataIn1 = 32'd4829
; 
32'd151582: dataIn1 = 32'd4831
; 
32'd151583: dataIn1 = 32'd6967
; 
32'd151584: dataIn1 = 32'd6969
; 
32'd151585: dataIn1 = 32'd6970
; 
32'd151586: dataIn1 = 32'd6971
; 
32'd151587: dataIn1 = 32'd2555
; 
32'd151588: dataIn1 = 32'd2618
; 
32'd151589: dataIn1 = 32'd4822
; 
32'd151590: dataIn1 = 32'd4832
; 
32'd151591: dataIn1 = 32'd4833
; 
32'd151592: dataIn1 = 32'd4834
; 
32'd151593: dataIn1 = 32'd4835
; 
32'd151594: dataIn1 = 32'd2555
; 
32'd151595: dataIn1 = 32'd2621
; 
32'd151596: dataIn1 = 32'd4646
; 
32'd151597: dataIn1 = 32'd4832
; 
32'd151598: dataIn1 = 32'd4833
; 
32'd151599: dataIn1 = 32'd4834
; 
32'd151600: dataIn1 = 32'd4836
; 
32'd151601: dataIn1 = 32'd2618
; 
32'd151602: dataIn1 = 32'd2621
; 
32'd151603: dataIn1 = 32'd4825
; 
32'd151604: dataIn1 = 32'd4832
; 
32'd151605: dataIn1 = 32'd4833
; 
32'd151606: dataIn1 = 32'd4834
; 
32'd151607: dataIn1 = 32'd4837
; 
32'd151608: dataIn1 = 32'd1073
; 
32'd151609: dataIn1 = 32'd2555
; 
32'd151610: dataIn1 = 32'd2556
; 
32'd151611: dataIn1 = 32'd4822
; 
32'd151612: dataIn1 = 32'd4832
; 
32'd151613: dataIn1 = 32'd4835
; 
32'd151614: dataIn1 = 32'd4
; 
32'd151615: dataIn1 = 32'd2621
; 
32'd151616: dataIn1 = 32'd4646
; 
32'd151617: dataIn1 = 32'd4833
; 
32'd151618: dataIn1 = 32'd4836
; 
32'd151619: dataIn1 = 32'd5858
; 
32'd151620: dataIn1 = 32'd5861
; 
32'd151621: dataIn1 = 32'd6945
; 
32'd151622: dataIn1 = 32'd1104
; 
32'd151623: dataIn1 = 32'd2621
; 
32'd151624: dataIn1 = 32'd4825
; 
32'd151625: dataIn1 = 32'd4834
; 
32'd151626: dataIn1 = 32'd4837
; 
32'd151627: dataIn1 = 32'd5857
; 
32'd151628: dataIn1 = 32'd5860
; 
32'd151629: dataIn1 = 32'd6935
; 
32'd151630: dataIn1 = 32'd6951
; 
32'd151631: dataIn1 = 32'd2554
; 
32'd151632: dataIn1 = 32'd4838
; 
32'd151633: dataIn1 = 32'd5318
; 
32'd151634: dataIn1 = 32'd5430
; 
32'd151635: dataIn1 = 32'd5947
; 
32'd151636: dataIn1 = 32'd5948
; 
32'd151637: dataIn1 = 32'd5950
; 
32'd151638: dataIn1 = 32'd2623
; 
32'd151639: dataIn1 = 32'd2624
; 
32'd151640: dataIn1 = 32'd4839
; 
32'd151641: dataIn1 = 32'd4840
; 
32'd151642: dataIn1 = 32'd4841
; 
32'd151643: dataIn1 = 32'd4842
; 
32'd151644: dataIn1 = 32'd4843
; 
32'd151645: dataIn1 = 32'd2624
; 
32'd151646: dataIn1 = 32'd4839
; 
32'd151647: dataIn1 = 32'd4840
; 
32'd151648: dataIn1 = 32'd4841
; 
32'd151649: dataIn1 = 32'd5953
; 
32'd151650: dataIn1 = 32'd5955
; 
32'd151651: dataIn1 = 32'd5957
; 
32'd151652: dataIn1 = 32'd2622
; 
32'd151653: dataIn1 = 32'd2623
; 
32'd151654: dataIn1 = 32'd4839
; 
32'd151655: dataIn1 = 32'd4840
; 
32'd151656: dataIn1 = 32'd4841
; 
32'd151657: dataIn1 = 32'd4846
; 
32'd151658: dataIn1 = 32'd4847
; 
32'd151659: dataIn1 = 32'd5957
; 
32'd151660: dataIn1 = 32'd1076
; 
32'd151661: dataIn1 = 32'd2624
; 
32'd151662: dataIn1 = 32'd4676
; 
32'd151663: dataIn1 = 32'd4839
; 
32'd151664: dataIn1 = 32'd4842
; 
32'd151665: dataIn1 = 32'd4843
; 
32'd151666: dataIn1 = 32'd4857
; 
32'd151667: dataIn1 = 32'd1076
; 
32'd151668: dataIn1 = 32'd2623
; 
32'd151669: dataIn1 = 32'd4839
; 
32'd151670: dataIn1 = 32'd4842
; 
32'd151671: dataIn1 = 32'd4843
; 
32'd151672: dataIn1 = 32'd4853
; 
32'd151673: dataIn1 = 32'd4856
; 
32'd151674: dataIn1 = 32'd2624
; 
32'd151675: dataIn1 = 32'd4844
; 
32'd151676: dataIn1 = 32'd5954
; 
32'd151677: dataIn1 = 32'd5955
; 
32'd151678: dataIn1 = 32'd5959
; 
32'd151679: dataIn1 = 32'd5987
; 
32'd151680: dataIn1 = 32'd5988
; 
32'd151681: dataIn1 = 32'd4845
; 
32'd151682: dataIn1 = 32'd5953
; 
32'd151683: dataIn1 = 32'd5954
; 
32'd151684: dataIn1 = 32'd5956
; 
32'd151685: dataIn1 = 32'd5958
; 
32'd151686: dataIn1 = 32'd5974
; 
32'd151687: dataIn1 = 32'd5975
; 
32'd151688: dataIn1 = 32'd1075
; 
32'd151689: dataIn1 = 32'd2623
; 
32'd151690: dataIn1 = 32'd4667
; 
32'd151691: dataIn1 = 32'd4841
; 
32'd151692: dataIn1 = 32'd4846
; 
32'd151693: dataIn1 = 32'd4847
; 
32'd151694: dataIn1 = 32'd4855
; 
32'd151695: dataIn1 = 32'd1075
; 
32'd151696: dataIn1 = 32'd2622
; 
32'd151697: dataIn1 = 32'd4662
; 
32'd151698: dataIn1 = 32'd4841
; 
32'd151699: dataIn1 = 32'd4846
; 
32'd151700: dataIn1 = 32'd4847
; 
32'd151701: dataIn1 = 32'd4850
; 
32'd151702: dataIn1 = 32'd5963
; 
32'd151703: dataIn1 = 32'd5979
; 
32'd151704: dataIn1 = 32'd4848
; 
32'd151705: dataIn1 = 32'd5961
; 
32'd151706: dataIn1 = 32'd5962
; 
32'd151707: dataIn1 = 32'd5966
; 
32'd151708: dataIn1 = 32'd5968
; 
32'd151709: dataIn1 = 32'd5970
; 
32'd151710: dataIn1 = 32'd5971
; 
32'd151711: dataIn1 = 32'd4849
; 
32'd151712: dataIn1 = 32'd5960
; 
32'd151713: dataIn1 = 32'd5962
; 
32'd151714: dataIn1 = 32'd5964
; 
32'd151715: dataIn1 = 32'd5967
; 
32'd151716: dataIn1 = 32'd5974
; 
32'd151717: dataIn1 = 32'd5976
; 
32'd151718: dataIn1 = 32'd4847
; 
32'd151719: dataIn1 = 32'd4850
; 
32'd151720: dataIn1 = 32'd5960
; 
32'd151721: dataIn1 = 32'd5961
; 
32'd151722: dataIn1 = 32'd5963
; 
32'd151723: dataIn1 = 32'd5965
; 
32'd151724: dataIn1 = 32'd5979
; 
32'd151725: dataIn1 = 32'd4851
; 
32'd151726: dataIn1 = 32'd5969
; 
32'd151727: dataIn1 = 32'd5971
; 
32'd151728: dataIn1 = 32'd5972
; 
32'd151729: dataIn1 = 32'd5973
; 
32'd151730: dataIn1 = 32'd7330
; 
32'd151731: dataIn1 = 32'd7331
; 
32'd151732: dataIn1 = 32'd4852
; 
32'd151733: dataIn1 = 32'd5975
; 
32'd151734: dataIn1 = 32'd5976
; 
32'd151735: dataIn1 = 32'd5977
; 
32'd151736: dataIn1 = 32'd5978
; 
32'd151737: dataIn1 = 32'd7326
; 
32'd151738: dataIn1 = 32'd7328
; 
32'd151739: dataIn1 = 32'd2570
; 
32'd151740: dataIn1 = 32'd2623
; 
32'd151741: dataIn1 = 32'd4843
; 
32'd151742: dataIn1 = 32'd4853
; 
32'd151743: dataIn1 = 32'd4854
; 
32'd151744: dataIn1 = 32'd4855
; 
32'd151745: dataIn1 = 32'd4856
; 
32'd151746: dataIn1 = 32'd2563
; 
32'd151747: dataIn1 = 32'd2570
; 
32'd151748: dataIn1 = 32'd4666
; 
32'd151749: dataIn1 = 32'd4682
; 
32'd151750: dataIn1 = 32'd4853
; 
32'd151751: dataIn1 = 32'd4854
; 
32'd151752: dataIn1 = 32'd4855
; 
32'd151753: dataIn1 = 32'd5981
; 
32'd151754: dataIn1 = 32'd2563
; 
32'd151755: dataIn1 = 32'd2623
; 
32'd151756: dataIn1 = 32'd4667
; 
32'd151757: dataIn1 = 32'd4846
; 
32'd151758: dataIn1 = 32'd4853
; 
32'd151759: dataIn1 = 32'd4854
; 
32'd151760: dataIn1 = 32'd4855
; 
32'd151761: dataIn1 = 32'd1076
; 
32'd151762: dataIn1 = 32'd2570
; 
32'd151763: dataIn1 = 32'd4843
; 
32'd151764: dataIn1 = 32'd4853
; 
32'd151765: dataIn1 = 32'd4856
; 
32'd151766: dataIn1 = 32'd10266
; 
32'd151767: dataIn1 = 32'd10268
; 
32'd151768: dataIn1 = 32'd2569
; 
32'd151769: dataIn1 = 32'd2624
; 
32'd151770: dataIn1 = 32'd4676
; 
32'd151771: dataIn1 = 32'd4842
; 
32'd151772: dataIn1 = 32'd4857
; 
32'd151773: dataIn1 = 32'd4858
; 
32'd151774: dataIn1 = 32'd4859
; 
32'd151775: dataIn1 = 32'd5983
; 
32'd151776: dataIn1 = 32'd2624
; 
32'd151777: dataIn1 = 32'd4857
; 
32'd151778: dataIn1 = 32'd4858
; 
32'd151779: dataIn1 = 32'd5983
; 
32'd151780: dataIn1 = 32'd5985
; 
32'd151781: dataIn1 = 32'd5986
; 
32'd151782: dataIn1 = 32'd5988
; 
32'd151783: dataIn1 = 32'd2569
; 
32'd151784: dataIn1 = 32'd4857
; 
32'd151785: dataIn1 = 32'd4859
; 
32'd151786: dataIn1 = 32'd5983
; 
32'd151787: dataIn1 = 32'd5984
; 
32'd151788: dataIn1 = 32'd5991
; 
32'd151789: dataIn1 = 32'd5992
; 
32'd151790: dataIn1 = 32'd4860
; 
32'd151791: dataIn1 = 32'd5986
; 
32'd151792: dataIn1 = 32'd5987
; 
32'd151793: dataIn1 = 32'd5989
; 
32'd151794: dataIn1 = 32'd5990
; 
32'd151795: dataIn1 = 32'd7344
; 
32'd151796: dataIn1 = 32'd7345
; 
32'd151797: dataIn1 = 32'd4861
; 
32'd151798: dataIn1 = 32'd5991
; 
32'd151799: dataIn1 = 32'd5993
; 
32'd151800: dataIn1 = 32'd5994
; 
32'd151801: dataIn1 = 32'd5995
; 
32'd151802: dataIn1 = 32'd7353
; 
32'd151803: dataIn1 = 32'd7354
; 
32'd151804: dataIn1 = 32'd4862
; 
32'd151805: dataIn1 = 32'd5997
; 
32'd151806: dataIn1 = 32'd5998
; 
32'd151807: dataIn1 = 32'd6002
; 
32'd151808: dataIn1 = 32'd6004
; 
32'd151809: dataIn1 = 32'd6006
; 
32'd151810: dataIn1 = 32'd6008
; 
32'd151811: dataIn1 = 32'd4863
; 
32'd151812: dataIn1 = 32'd5996
; 
32'd151813: dataIn1 = 32'd5998
; 
32'd151814: dataIn1 = 32'd6000
; 
32'd151815: dataIn1 = 32'd6003
; 
32'd151816: dataIn1 = 32'd6009
; 
32'd151817: dataIn1 = 32'd6011
; 
32'd151818: dataIn1 = 32'd4864
; 
32'd151819: dataIn1 = 32'd5996
; 
32'd151820: dataIn1 = 32'd5997
; 
32'd151821: dataIn1 = 32'd5999
; 
32'd151822: dataIn1 = 32'd6001
; 
32'd151823: dataIn1 = 32'd6014
; 
32'd151824: dataIn1 = 32'd6015
; 
32'd151825: dataIn1 = 32'd447
; 
32'd151826: dataIn1 = 32'd3913
; 
32'd151827: dataIn1 = 32'd4865
; 
32'd151828: dataIn1 = 32'd4881
; 
32'd151829: dataIn1 = 32'd6007
; 
32'd151830: dataIn1 = 32'd6008
; 
32'd151831: dataIn1 = 32'd6700
; 
32'd151832: dataIn1 = 32'd447
; 
32'd151833: dataIn1 = 32'd4866
; 
32'd151834: dataIn1 = 32'd6005
; 
32'd151835: dataIn1 = 32'd6006
; 
32'd151836: dataIn1 = 32'd6700
; 
32'd151837: dataIn1 = 32'd6701
; 
32'd151838: dataIn1 = 32'd6732
; 
32'd151839: dataIn1 = 32'd4671
; 
32'd151840: dataIn1 = 32'd4867
; 
32'd151841: dataIn1 = 32'd4882
; 
32'd151842: dataIn1 = 32'd6010
; 
32'd151843: dataIn1 = 32'd6011
; 
32'd151844: dataIn1 = 32'd6013
; 
32'd151845: dataIn1 = 32'd6702
; 
32'd151846: dataIn1 = 32'd4868
; 
32'd151847: dataIn1 = 32'd6009
; 
32'd151848: dataIn1 = 32'd6010
; 
32'd151849: dataIn1 = 32'd6012
; 
32'd151850: dataIn1 = 32'd6035
; 
32'd151851: dataIn1 = 32'd6036
; 
32'd151852: dataIn1 = 32'd6697
; 
32'd151853: dataIn1 = 32'd4869
; 
32'd151854: dataIn1 = 32'd6015
; 
32'd151855: dataIn1 = 32'd6016
; 
32'd151856: dataIn1 = 32'd6018
; 
32'd151857: dataIn1 = 32'd6020
; 
32'd151858: dataIn1 = 32'd6057
; 
32'd151859: dataIn1 = 32'd6058
; 
32'd151860: dataIn1 = 32'd4870
; 
32'd151861: dataIn1 = 32'd6014
; 
32'd151862: dataIn1 = 32'd6016
; 
32'd151863: dataIn1 = 32'd6017
; 
32'd151864: dataIn1 = 32'd6019
; 
32'd151865: dataIn1 = 32'd6038
; 
32'd151866: dataIn1 = 32'd6040
; 
32'd151867: dataIn1 = 32'd4871
; 
32'd151868: dataIn1 = 32'd6022
; 
32'd151869: dataIn1 = 32'd6023
; 
32'd151870: dataIn1 = 32'd6027
; 
32'd151871: dataIn1 = 32'd6029
; 
32'd151872: dataIn1 = 32'd6031
; 
32'd151873: dataIn1 = 32'd6032
; 
32'd151874: dataIn1 = 32'd4872
; 
32'd151875: dataIn1 = 32'd6021
; 
32'd151876: dataIn1 = 32'd6023
; 
32'd151877: dataIn1 = 32'd6025
; 
32'd151878: dataIn1 = 32'd6028
; 
32'd151879: dataIn1 = 32'd6035
; 
32'd151880: dataIn1 = 32'd6037
; 
32'd151881: dataIn1 = 32'd4873
; 
32'd151882: dataIn1 = 32'd6021
; 
32'd151883: dataIn1 = 32'd6022
; 
32'd151884: dataIn1 = 32'd6024
; 
32'd151885: dataIn1 = 32'd6026
; 
32'd151886: dataIn1 = 32'd6038
; 
32'd151887: dataIn1 = 32'd6039
; 
32'd151888: dataIn1 = 32'd4874
; 
32'd151889: dataIn1 = 32'd6030
; 
32'd151890: dataIn1 = 32'd6031
; 
32'd151891: dataIn1 = 32'd6033
; 
32'd151892: dataIn1 = 32'd6034
; 
32'd151893: dataIn1 = 32'd7276
; 
32'd151894: dataIn1 = 32'd7277
; 
32'd151895: dataIn1 = 32'd4875
; 
32'd151896: dataIn1 = 32'd6039
; 
32'd151897: dataIn1 = 32'd6040
; 
32'd151898: dataIn1 = 32'd6041
; 
32'd151899: dataIn1 = 32'd6042
; 
32'd151900: dataIn1 = 32'd7279
; 
32'd151901: dataIn1 = 32'd7281
; 
32'd151902: dataIn1 = 32'd4876
; 
32'd151903: dataIn1 = 32'd6047
; 
32'd151904: dataIn1 = 32'd6048
; 
32'd151905: dataIn1 = 32'd6050
; 
32'd151906: dataIn1 = 32'd6051
; 
32'd151907: dataIn1 = 32'd6696
; 
32'd151908: dataIn1 = 32'd6701
; 
32'd151909: dataIn1 = 32'd4877
; 
32'd151910: dataIn1 = 32'd6043
; 
32'd151911: dataIn1 = 32'd6045
; 
32'd151912: dataIn1 = 32'd6049
; 
32'd151913: dataIn1 = 32'd6051
; 
32'd151914: dataIn1 = 32'd6052
; 
32'd151915: dataIn1 = 32'd6054
; 
32'd151916: dataIn1 = 32'd4878
; 
32'd151917: dataIn1 = 32'd6043
; 
32'd151918: dataIn1 = 32'd6044
; 
32'd151919: dataIn1 = 32'd6046
; 
32'd151920: dataIn1 = 32'd6047
; 
32'd151921: dataIn1 = 32'd6056
; 
32'd151922: dataIn1 = 32'd6057
; 
32'd151923: dataIn1 = 32'd4879
; 
32'd151924: dataIn1 = 32'd6052
; 
32'd151925: dataIn1 = 32'd6053
; 
32'd151926: dataIn1 = 32'd6055
; 
32'd151927: dataIn1 = 32'd6703
; 
32'd151928: dataIn1 = 32'd7256
; 
32'd151929: dataIn1 = 32'd7257
; 
32'd151930: dataIn1 = 32'd4880
; 
32'd151931: dataIn1 = 32'd6056
; 
32'd151932: dataIn1 = 32'd6058
; 
32'd151933: dataIn1 = 32'd6059
; 
32'd151934: dataIn1 = 32'd6060
; 
32'd151935: dataIn1 = 32'd7260
; 
32'd151936: dataIn1 = 32'd7261
; 
32'd151937: dataIn1 = 32'd2306
; 
32'd151938: dataIn1 = 32'd2629
; 
32'd151939: dataIn1 = 32'd3913
; 
32'd151940: dataIn1 = 32'd4865
; 
32'd151941: dataIn1 = 32'd4881
; 
32'd151942: dataIn1 = 32'd4882
; 
32'd151943: dataIn1 = 32'd4883
; 
32'd151944: dataIn1 = 32'd6007
; 
32'd151945: dataIn1 = 32'd6064
; 
32'd151946: dataIn1 = 32'd2564
; 
32'd151947: dataIn1 = 32'd2629
; 
32'd151948: dataIn1 = 32'd4671
; 
32'd151949: dataIn1 = 32'd4867
; 
32'd151950: dataIn1 = 32'd4881
; 
32'd151951: dataIn1 = 32'd4882
; 
32'd151952: dataIn1 = 32'd4883
; 
32'd151953: dataIn1 = 32'd6013
; 
32'd151954: dataIn1 = 32'd2564
; 
32'd151955: dataIn1 = 32'd4881
; 
32'd151956: dataIn1 = 32'd4882
; 
32'd151957: dataIn1 = 32'd4883
; 
32'd151958: dataIn1 = 32'd6061
; 
32'd151959: dataIn1 = 32'd6062
; 
32'd151960: dataIn1 = 32'd6064
; 
32'd151961: dataIn1 = 32'd2633
; 
32'd151962: dataIn1 = 32'd2634
; 
32'd151963: dataIn1 = 32'd4884
; 
32'd151964: dataIn1 = 32'd4885
; 
32'd151965: dataIn1 = 32'd4886
; 
32'd151966: dataIn1 = 32'd4887
; 
32'd151967: dataIn1 = 32'd4888
; 
32'd151968: dataIn1 = 32'd2632
; 
32'd151969: dataIn1 = 32'd2634
; 
32'd151970: dataIn1 = 32'd4884
; 
32'd151971: dataIn1 = 32'd4885
; 
32'd151972: dataIn1 = 32'd4886
; 
32'd151973: dataIn1 = 32'd4889
; 
32'd151974: dataIn1 = 32'd4890
; 
32'd151975: dataIn1 = 32'd2632
; 
32'd151976: dataIn1 = 32'd2633
; 
32'd151977: dataIn1 = 32'd4884
; 
32'd151978: dataIn1 = 32'd4885
; 
32'd151979: dataIn1 = 32'd4886
; 
32'd151980: dataIn1 = 32'd4891
; 
32'd151981: dataIn1 = 32'd4892
; 
32'd151982: dataIn1 = 32'd9613
; 
32'd151983: dataIn1 = 32'd1077
; 
32'd151984: dataIn1 = 32'd2634
; 
32'd151985: dataIn1 = 32'd3431
; 
32'd151986: dataIn1 = 32'd4884
; 
32'd151987: dataIn1 = 32'd4887
; 
32'd151988: dataIn1 = 32'd4888
; 
32'd151989: dataIn1 = 32'd1077
; 
32'd151990: dataIn1 = 32'd2633
; 
32'd151991: dataIn1 = 32'd4681
; 
32'd151992: dataIn1 = 32'd4884
; 
32'd151993: dataIn1 = 32'd4887
; 
32'd151994: dataIn1 = 32'd4888
; 
32'd151995: dataIn1 = 32'd4898
; 
32'd151996: dataIn1 = 32'd1078
; 
32'd151997: dataIn1 = 32'd2634
; 
32'd151998: dataIn1 = 32'd3432
; 
32'd151999: dataIn1 = 32'd4885
; 
32'd152000: dataIn1 = 32'd4889
; 
32'd152001: dataIn1 = 32'd4890
; 
32'd152002: dataIn1 = 32'd1078
; 
32'd152003: dataIn1 = 32'd2632
; 
32'd152004: dataIn1 = 32'd4689
; 
32'd152005: dataIn1 = 32'd4885
; 
32'd152006: dataIn1 = 32'd4889
; 
32'd152007: dataIn1 = 32'd4890
; 
32'd152008: dataIn1 = 32'd4894
; 
32'd152009: dataIn1 = 32'd2633
; 
32'd152010: dataIn1 = 32'd4886
; 
32'd152011: dataIn1 = 32'd4891
; 
32'd152012: dataIn1 = 32'd4900
; 
32'd152013: dataIn1 = 32'd9612
; 
32'd152014: dataIn1 = 32'd9613
; 
32'd152015: dataIn1 = 32'd9763
; 
32'd152016: dataIn1 = 32'd2632
; 
32'd152017: dataIn1 = 32'd4886
; 
32'd152018: dataIn1 = 32'd4892
; 
32'd152019: dataIn1 = 32'd9611
; 
32'd152020: dataIn1 = 32'd9613
; 
32'd152021: dataIn1 = 32'd9620
; 
32'd152022: dataIn1 = 32'd9622
; 
32'd152023: dataIn1 = 32'd2573
; 
32'd152024: dataIn1 = 32'd4893
; 
32'd152025: dataIn1 = 32'd4894
; 
32'd152026: dataIn1 = 32'd9615
; 
32'd152027: dataIn1 = 32'd9616
; 
32'd152028: dataIn1 = 32'd9618
; 
32'd152029: dataIn1 = 32'd9619
; 
32'd152030: dataIn1 = 32'd2573
; 
32'd152031: dataIn1 = 32'd2632
; 
32'd152032: dataIn1 = 32'd4689
; 
32'd152033: dataIn1 = 32'd4890
; 
32'd152034: dataIn1 = 32'd4893
; 
32'd152035: dataIn1 = 32'd4894
; 
32'd152036: dataIn1 = 32'd4895
; 
32'd152037: dataIn1 = 32'd9615
; 
32'd152038: dataIn1 = 32'd2632
; 
32'd152039: dataIn1 = 32'd4894
; 
32'd152040: dataIn1 = 32'd4895
; 
32'd152041: dataIn1 = 32'd9614
; 
32'd152042: dataIn1 = 32'd9615
; 
32'd152043: dataIn1 = 32'd9620
; 
32'd152044: dataIn1 = 32'd9621
; 
32'd152045: dataIn1 = 32'd4896
; 
32'd152046: dataIn1 = 32'd7485
; 
32'd152047: dataIn1 = 32'd7486
; 
32'd152048: dataIn1 = 32'd7488
; 
32'd152049: dataIn1 = 32'd7489
; 
32'd152050: dataIn1 = 32'd9617
; 
32'd152051: dataIn1 = 32'd9618
; 
32'd152052: dataIn1 = 32'd4897
; 
32'd152053: dataIn1 = 32'd7490
; 
32'd152054: dataIn1 = 32'd7492
; 
32'd152055: dataIn1 = 32'd7493
; 
32'd152056: dataIn1 = 32'd7494
; 
32'd152057: dataIn1 = 32'd9621
; 
32'd152058: dataIn1 = 32'd9622
; 
32'd152059: dataIn1 = 32'd2568
; 
32'd152060: dataIn1 = 32'd2633
; 
32'd152061: dataIn1 = 32'd4681
; 
32'd152062: dataIn1 = 32'd4888
; 
32'd152063: dataIn1 = 32'd4898
; 
32'd152064: dataIn1 = 32'd4899
; 
32'd152065: dataIn1 = 32'd4900
; 
32'd152066: dataIn1 = 32'd2568
; 
32'd152067: dataIn1 = 32'd2636
; 
32'd152068: dataIn1 = 32'd4679
; 
32'd152069: dataIn1 = 32'd4898
; 
32'd152070: dataIn1 = 32'd4899
; 
32'd152071: dataIn1 = 32'd4900
; 
32'd152072: dataIn1 = 32'd4901
; 
32'd152073: dataIn1 = 32'd6066
; 
32'd152074: dataIn1 = 32'd7461
; 
32'd152075: dataIn1 = 32'd2633
; 
32'd152076: dataIn1 = 32'd2636
; 
32'd152077: dataIn1 = 32'd4891
; 
32'd152078: dataIn1 = 32'd4898
; 
32'd152079: dataIn1 = 32'd4899
; 
32'd152080: dataIn1 = 32'd4900
; 
32'd152081: dataIn1 = 32'd4902
; 
32'd152082: dataIn1 = 32'd7471
; 
32'd152083: dataIn1 = 32'd9763
; 
32'd152084: dataIn1 = 32'd4899
; 
32'd152085: dataIn1 = 32'd4901
; 
32'd152086: dataIn1 = 32'd6065
; 
32'd152087: dataIn1 = 32'd6066
; 
32'd152088: dataIn1 = 32'd7458
; 
32'd152089: dataIn1 = 32'd7459
; 
32'd152090: dataIn1 = 32'd7461
; 
32'd152091: dataIn1 = 32'd4900
; 
32'd152092: dataIn1 = 32'd4902
; 
32'd152093: dataIn1 = 32'd7469
; 
32'd152094: dataIn1 = 32'd7470
; 
32'd152095: dataIn1 = 32'd7471
; 
32'd152096: dataIn1 = 32'd7472
; 
32'd152097: dataIn1 = 32'd9763
; 
32'd152098: dataIn1 = 32'd2638
; 
32'd152099: dataIn1 = 32'd2639
; 
32'd152100: dataIn1 = 32'd4903
; 
32'd152101: dataIn1 = 32'd4904
; 
32'd152102: dataIn1 = 32'd4905
; 
32'd152103: dataIn1 = 32'd4906
; 
32'd152104: dataIn1 = 32'd4907
; 
32'd152105: dataIn1 = 32'd2637
; 
32'd152106: dataIn1 = 32'd2639
; 
32'd152107: dataIn1 = 32'd4903
; 
32'd152108: dataIn1 = 32'd4904
; 
32'd152109: dataIn1 = 32'd4905
; 
32'd152110: dataIn1 = 32'd4908
; 
32'd152111: dataIn1 = 32'd4909
; 
32'd152112: dataIn1 = 32'd9624
; 
32'd152113: dataIn1 = 32'd2637
; 
32'd152114: dataIn1 = 32'd2638
; 
32'd152115: dataIn1 = 32'd4903
; 
32'd152116: dataIn1 = 32'd4904
; 
32'd152117: dataIn1 = 32'd4905
; 
32'd152118: dataIn1 = 32'd4910
; 
32'd152119: dataIn1 = 32'd4911
; 
32'd152120: dataIn1 = 32'd1080
; 
32'd152121: dataIn1 = 32'd2639
; 
32'd152122: dataIn1 = 32'd4696
; 
32'd152123: dataIn1 = 32'd4903
; 
32'd152124: dataIn1 = 32'd4906
; 
32'd152125: dataIn1 = 32'd4907
; 
32'd152126: dataIn1 = 32'd4917
; 
32'd152127: dataIn1 = 32'd1080
; 
32'd152128: dataIn1 = 32'd2638
; 
32'd152129: dataIn1 = 32'd3477
; 
32'd152130: dataIn1 = 32'd4903
; 
32'd152131: dataIn1 = 32'd4906
; 
32'd152132: dataIn1 = 32'd4907
; 
32'd152133: dataIn1 = 32'd2639
; 
32'd152134: dataIn1 = 32'd4904
; 
32'd152135: dataIn1 = 32'd4908
; 
32'd152136: dataIn1 = 32'd9624
; 
32'd152137: dataIn1 = 32'd9625
; 
32'd152138: dataIn1 = 32'd9639
; 
32'd152139: dataIn1 = 32'd9640
; 
32'd152140: dataIn1 = 32'd2637
; 
32'd152141: dataIn1 = 32'd4904
; 
32'd152142: dataIn1 = 32'd4909
; 
32'd152143: dataIn1 = 32'd9623
; 
32'd152144: dataIn1 = 32'd9624
; 
32'd152145: dataIn1 = 32'd9632
; 
32'd152146: dataIn1 = 32'd9633
; 
32'd152147: dataIn1 = 32'd1079
; 
32'd152148: dataIn1 = 32'd2638
; 
32'd152149: dataIn1 = 32'd3473
; 
32'd152150: dataIn1 = 32'd4905
; 
32'd152151: dataIn1 = 32'd4910
; 
32'd152152: dataIn1 = 32'd4911
; 
32'd152153: dataIn1 = 32'd1079
; 
32'd152154: dataIn1 = 32'd2637
; 
32'd152155: dataIn1 = 32'd4691
; 
32'd152156: dataIn1 = 32'd4905
; 
32'd152157: dataIn1 = 32'd4910
; 
32'd152158: dataIn1 = 32'd4911
; 
32'd152159: dataIn1 = 32'd4914
; 
32'd152160: dataIn1 = 32'd2572
; 
32'd152161: dataIn1 = 32'd4912
; 
32'd152162: dataIn1 = 32'd4914
; 
32'd152163: dataIn1 = 32'd9627
; 
32'd152164: dataIn1 = 32'd9628
; 
32'd152165: dataIn1 = 32'd9630
; 
32'd152166: dataIn1 = 32'd9631
; 
32'd152167: dataIn1 = 32'd2637
; 
32'd152168: dataIn1 = 32'd4913
; 
32'd152169: dataIn1 = 32'd4914
; 
32'd152170: dataIn1 = 32'd9626
; 
32'd152171: dataIn1 = 32'd9628
; 
32'd152172: dataIn1 = 32'd9632
; 
32'd152173: dataIn1 = 32'd9634
; 
32'd152174: dataIn1 = 32'd2572
; 
32'd152175: dataIn1 = 32'd2637
; 
32'd152176: dataIn1 = 32'd4691
; 
32'd152177: dataIn1 = 32'd4911
; 
32'd152178: dataIn1 = 32'd4912
; 
32'd152179: dataIn1 = 32'd4913
; 
32'd152180: dataIn1 = 32'd4914
; 
32'd152181: dataIn1 = 32'd9628
; 
32'd152182: dataIn1 = 32'd4915
; 
32'd152183: dataIn1 = 32'd7574
; 
32'd152184: dataIn1 = 32'd7575
; 
32'd152185: dataIn1 = 32'd7576
; 
32'd152186: dataIn1 = 32'd7577
; 
32'd152187: dataIn1 = 32'd9629
; 
32'd152188: dataIn1 = 32'd9631
; 
32'd152189: dataIn1 = 32'd4916
; 
32'd152190: dataIn1 = 32'd7568
; 
32'd152191: dataIn1 = 32'd7570
; 
32'd152192: dataIn1 = 32'd7571
; 
32'd152193: dataIn1 = 32'd7572
; 
32'd152194: dataIn1 = 32'd9633
; 
32'd152195: dataIn1 = 32'd9634
; 
32'd152196: dataIn1 = 32'd2576
; 
32'd152197: dataIn1 = 32'd2639
; 
32'd152198: dataIn1 = 32'd4696
; 
32'd152199: dataIn1 = 32'd4906
; 
32'd152200: dataIn1 = 32'd4917
; 
32'd152201: dataIn1 = 32'd4918
; 
32'd152202: dataIn1 = 32'd4919
; 
32'd152203: dataIn1 = 32'd9635
; 
32'd152204: dataIn1 = 32'd2639
; 
32'd152205: dataIn1 = 32'd4917
; 
32'd152206: dataIn1 = 32'd4918
; 
32'd152207: dataIn1 = 32'd9635
; 
32'd152208: dataIn1 = 32'd9637
; 
32'd152209: dataIn1 = 32'd9638
; 
32'd152210: dataIn1 = 32'd9640
; 
32'd152211: dataIn1 = 32'd2576
; 
32'd152212: dataIn1 = 32'd4917
; 
32'd152213: dataIn1 = 32'd4919
; 
32'd152214: dataIn1 = 32'd9635
; 
32'd152215: dataIn1 = 32'd9636
; 
32'd152216: dataIn1 = 32'd9641
; 
32'd152217: dataIn1 = 32'd9642
; 
32'd152218: dataIn1 = 32'd4920
; 
32'd152219: dataIn1 = 32'd7590
; 
32'd152220: dataIn1 = 32'd7591
; 
32'd152221: dataIn1 = 32'd7593
; 
32'd152222: dataIn1 = 32'd7594
; 
32'd152223: dataIn1 = 32'd9638
; 
32'd152224: dataIn1 = 32'd9639
; 
32'd152225: dataIn1 = 32'd4921
; 
32'd152226: dataIn1 = 32'd7601
; 
32'd152227: dataIn1 = 32'd7602
; 
32'd152228: dataIn1 = 32'd7604
; 
32'd152229: dataIn1 = 32'd7606
; 
32'd152230: dataIn1 = 32'd9641
; 
32'd152231: dataIn1 = 32'd9643
; 
32'd152232: dataIn1 = 32'd2643
; 
32'd152233: dataIn1 = 32'd2644
; 
32'd152234: dataIn1 = 32'd4922
; 
32'd152235: dataIn1 = 32'd4923
; 
32'd152236: dataIn1 = 32'd4924
; 
32'd152237: dataIn1 = 32'd4925
; 
32'd152238: dataIn1 = 32'd4926
; 
32'd152239: dataIn1 = 32'd2642
; 
32'd152240: dataIn1 = 32'd2644
; 
32'd152241: dataIn1 = 32'd4922
; 
32'd152242: dataIn1 = 32'd4923
; 
32'd152243: dataIn1 = 32'd4924
; 
32'd152244: dataIn1 = 32'd4927
; 
32'd152245: dataIn1 = 32'd4928
; 
32'd152246: dataIn1 = 32'd2642
; 
32'd152247: dataIn1 = 32'd2643
; 
32'd152248: dataIn1 = 32'd4922
; 
32'd152249: dataIn1 = 32'd4923
; 
32'd152250: dataIn1 = 32'd4924
; 
32'd152251: dataIn1 = 32'd4929
; 
32'd152252: dataIn1 = 32'd4930
; 
32'd152253: dataIn1 = 32'd9646
; 
32'd152254: dataIn1 = 32'd1081
; 
32'd152255: dataIn1 = 32'd2644
; 
32'd152256: dataIn1 = 32'd3489
; 
32'd152257: dataIn1 = 32'd4922
; 
32'd152258: dataIn1 = 32'd4925
; 
32'd152259: dataIn1 = 32'd4926
; 
32'd152260: dataIn1 = 32'd1081
; 
32'd152261: dataIn1 = 32'd2643
; 
32'd152262: dataIn1 = 32'd4701
; 
32'd152263: dataIn1 = 32'd4922
; 
32'd152264: dataIn1 = 32'd4925
; 
32'd152265: dataIn1 = 32'd4926
; 
32'd152266: dataIn1 = 32'd4936
; 
32'd152267: dataIn1 = 32'd1082
; 
32'd152268: dataIn1 = 32'd2644
; 
32'd152269: dataIn1 = 32'd3493
; 
32'd152270: dataIn1 = 32'd4923
; 
32'd152271: dataIn1 = 32'd4927
; 
32'd152272: dataIn1 = 32'd4928
; 
32'd152273: dataIn1 = 32'd1082
; 
32'd152274: dataIn1 = 32'd2642
; 
32'd152275: dataIn1 = 32'd4707
; 
32'd152276: dataIn1 = 32'd4923
; 
32'd152277: dataIn1 = 32'd4927
; 
32'd152278: dataIn1 = 32'd4928
; 
32'd152279: dataIn1 = 32'd4932
; 
32'd152280: dataIn1 = 32'd2643
; 
32'd152281: dataIn1 = 32'd4924
; 
32'd152282: dataIn1 = 32'd4929
; 
32'd152283: dataIn1 = 32'd9645
; 
32'd152284: dataIn1 = 32'd9646
; 
32'd152285: dataIn1 = 32'd9663
; 
32'd152286: dataIn1 = 32'd9664
; 
32'd152287: dataIn1 = 32'd2642
; 
32'd152288: dataIn1 = 32'd4924
; 
32'd152289: dataIn1 = 32'd4930
; 
32'd152290: dataIn1 = 32'd9644
; 
32'd152291: dataIn1 = 32'd9646
; 
32'd152292: dataIn1 = 32'd9653
; 
32'd152293: dataIn1 = 32'd9655
; 
32'd152294: dataIn1 = 32'd2579
; 
32'd152295: dataIn1 = 32'd4931
; 
32'd152296: dataIn1 = 32'd4932
; 
32'd152297: dataIn1 = 32'd9648
; 
32'd152298: dataIn1 = 32'd9649
; 
32'd152299: dataIn1 = 32'd9651
; 
32'd152300: dataIn1 = 32'd9652
; 
32'd152301: dataIn1 = 32'd2579
; 
32'd152302: dataIn1 = 32'd2642
; 
32'd152303: dataIn1 = 32'd4707
; 
32'd152304: dataIn1 = 32'd4928
; 
32'd152305: dataIn1 = 32'd4931
; 
32'd152306: dataIn1 = 32'd4932
; 
32'd152307: dataIn1 = 32'd4933
; 
32'd152308: dataIn1 = 32'd9648
; 
32'd152309: dataIn1 = 32'd2642
; 
32'd152310: dataIn1 = 32'd4932
; 
32'd152311: dataIn1 = 32'd4933
; 
32'd152312: dataIn1 = 32'd9647
; 
32'd152313: dataIn1 = 32'd9648
; 
32'd152314: dataIn1 = 32'd9653
; 
32'd152315: dataIn1 = 32'd9654
; 
32'd152316: dataIn1 = 32'd4934
; 
32'd152317: dataIn1 = 32'd7738
; 
32'd152318: dataIn1 = 32'd7739
; 
32'd152319: dataIn1 = 32'd7741
; 
32'd152320: dataIn1 = 32'd7742
; 
32'd152321: dataIn1 = 32'd9650
; 
32'd152322: dataIn1 = 32'd9651
; 
32'd152323: dataIn1 = 32'd4935
; 
32'd152324: dataIn1 = 32'd7743
; 
32'd152325: dataIn1 = 32'd7745
; 
32'd152326: dataIn1 = 32'd7746
; 
32'd152327: dataIn1 = 32'd7747
; 
32'd152328: dataIn1 = 32'd9654
; 
32'd152329: dataIn1 = 32'd9655
; 
32'd152330: dataIn1 = 32'd2574
; 
32'd152331: dataIn1 = 32'd2643
; 
32'd152332: dataIn1 = 32'd4701
; 
32'd152333: dataIn1 = 32'd4926
; 
32'd152334: dataIn1 = 32'd4936
; 
32'd152335: dataIn1 = 32'd4937
; 
32'd152336: dataIn1 = 32'd4938
; 
32'd152337: dataIn1 = 32'd9656
; 
32'd152338: dataIn1 = 32'd2574
; 
32'd152339: dataIn1 = 32'd4936
; 
32'd152340: dataIn1 = 32'd4937
; 
32'd152341: dataIn1 = 32'd9656
; 
32'd152342: dataIn1 = 32'd9658
; 
32'd152343: dataIn1 = 32'd9659
; 
32'd152344: dataIn1 = 32'd9661
; 
32'd152345: dataIn1 = 32'd2643
; 
32'd152346: dataIn1 = 32'd4936
; 
32'd152347: dataIn1 = 32'd4938
; 
32'd152348: dataIn1 = 32'd9656
; 
32'd152349: dataIn1 = 32'd9657
; 
32'd152350: dataIn1 = 32'd9662
; 
32'd152351: dataIn1 = 32'd9663
; 
32'd152352: dataIn1 = 32'd4939
; 
32'd152353: dataIn1 = 32'd7709
; 
32'd152354: dataIn1 = 32'd7710
; 
32'd152355: dataIn1 = 32'd7712
; 
32'd152356: dataIn1 = 32'd7714
; 
32'd152357: dataIn1 = 32'd9659
; 
32'd152358: dataIn1 = 32'd9660
; 
32'd152359: dataIn1 = 32'd4940
; 
32'd152360: dataIn1 = 32'd7722
; 
32'd152361: dataIn1 = 32'd7723
; 
32'd152362: dataIn1 = 32'd7724
; 
32'd152363: dataIn1 = 32'd7725
; 
32'd152364: dataIn1 = 32'd9662
; 
32'd152365: dataIn1 = 32'd9664
; 
32'd152366: dataIn1 = 32'd2648
; 
32'd152367: dataIn1 = 32'd2649
; 
32'd152368: dataIn1 = 32'd4941
; 
32'd152369: dataIn1 = 32'd4942
; 
32'd152370: dataIn1 = 32'd4943
; 
32'd152371: dataIn1 = 32'd4944
; 
32'd152372: dataIn1 = 32'd4945
; 
32'd152373: dataIn1 = 32'd2647
; 
32'd152374: dataIn1 = 32'd2649
; 
32'd152375: dataIn1 = 32'd4941
; 
32'd152376: dataIn1 = 32'd4942
; 
32'd152377: dataIn1 = 32'd4943
; 
32'd152378: dataIn1 = 32'd4946
; 
32'd152379: dataIn1 = 32'd4947
; 
32'd152380: dataIn1 = 32'd2647
; 
32'd152381: dataIn1 = 32'd2648
; 
32'd152382: dataIn1 = 32'd4941
; 
32'd152383: dataIn1 = 32'd4942
; 
32'd152384: dataIn1 = 32'd4943
; 
32'd152385: dataIn1 = 32'd4948
; 
32'd152386: dataIn1 = 32'd4949
; 
32'd152387: dataIn1 = 32'd1084
; 
32'd152388: dataIn1 = 32'd2649
; 
32'd152389: dataIn1 = 32'd4714
; 
32'd152390: dataIn1 = 32'd4941
; 
32'd152391: dataIn1 = 32'd4944
; 
32'd152392: dataIn1 = 32'd4945
; 
32'd152393: dataIn1 = 32'd4955
; 
32'd152394: dataIn1 = 32'd1084
; 
32'd152395: dataIn1 = 32'd2648
; 
32'd152396: dataIn1 = 32'd3505
; 
32'd152397: dataIn1 = 32'd4941
; 
32'd152398: dataIn1 = 32'd4944
; 
32'd152399: dataIn1 = 32'd4945
; 
32'd152400: dataIn1 = 32'd1110
; 
32'd152401: dataIn1 = 32'd2649
; 
32'd152402: dataIn1 = 32'd4942
; 
32'd152403: dataIn1 = 32'd4946
; 
32'd152404: dataIn1 = 32'd4947
; 
32'd152405: dataIn1 = 32'd4956
; 
32'd152406: dataIn1 = 32'd4958
; 
32'd152407: dataIn1 = 32'd7846
; 
32'd152408: dataIn1 = 32'd1110
; 
32'd152409: dataIn1 = 32'd2647
; 
32'd152410: dataIn1 = 32'd4942
; 
32'd152411: dataIn1 = 32'd4946
; 
32'd152412: dataIn1 = 32'd4947
; 
32'd152413: dataIn1 = 32'd4951
; 
32'd152414: dataIn1 = 32'd4954
; 
32'd152415: dataIn1 = 32'd7824
; 
32'd152416: dataIn1 = 32'd1083
; 
32'd152417: dataIn1 = 32'd2648
; 
32'd152418: dataIn1 = 32'd3503
; 
32'd152419: dataIn1 = 32'd4943
; 
32'd152420: dataIn1 = 32'd4948
; 
32'd152421: dataIn1 = 32'd4949
; 
32'd152422: dataIn1 = 32'd1083
; 
32'd152423: dataIn1 = 32'd2647
; 
32'd152424: dataIn1 = 32'd4709
; 
32'd152425: dataIn1 = 32'd4943
; 
32'd152426: dataIn1 = 32'd4948
; 
32'd152427: dataIn1 = 32'd4949
; 
32'd152428: dataIn1 = 32'd4952
; 
32'd152429: dataIn1 = 32'd2578
; 
32'd152430: dataIn1 = 32'd4950
; 
32'd152431: dataIn1 = 32'd4951
; 
32'd152432: dataIn1 = 32'd4952
; 
32'd152433: dataIn1 = 32'd9666
; 
32'd152434: dataIn1 = 32'd9667
; 
32'd152435: dataIn1 = 32'd9764
; 
32'd152436: dataIn1 = 32'd2647
; 
32'd152437: dataIn1 = 32'd2650
; 
32'd152438: dataIn1 = 32'd4947
; 
32'd152439: dataIn1 = 32'd4950
; 
32'd152440: dataIn1 = 32'd4951
; 
32'd152441: dataIn1 = 32'd4952
; 
32'd152442: dataIn1 = 32'd4954
; 
32'd152443: dataIn1 = 32'd7825
; 
32'd152444: dataIn1 = 32'd9764
; 
32'd152445: dataIn1 = 32'd2578
; 
32'd152446: dataIn1 = 32'd2647
; 
32'd152447: dataIn1 = 32'd4709
; 
32'd152448: dataIn1 = 32'd4949
; 
32'd152449: dataIn1 = 32'd4950
; 
32'd152450: dataIn1 = 32'd4951
; 
32'd152451: dataIn1 = 32'd4952
; 
32'd152452: dataIn1 = 32'd4953
; 
32'd152453: dataIn1 = 32'd7827
; 
32'd152454: dataIn1 = 32'd7828
; 
32'd152455: dataIn1 = 32'd7829
; 
32'd152456: dataIn1 = 32'd7830
; 
32'd152457: dataIn1 = 32'd9665
; 
32'd152458: dataIn1 = 32'd9667
; 
32'd152459: dataIn1 = 32'd4947
; 
32'd152460: dataIn1 = 32'd4951
; 
32'd152461: dataIn1 = 32'd4954
; 
32'd152462: dataIn1 = 32'd7821
; 
32'd152463: dataIn1 = 32'd7823
; 
32'd152464: dataIn1 = 32'd7824
; 
32'd152465: dataIn1 = 32'd7825
; 
32'd152466: dataIn1 = 32'd2582
; 
32'd152467: dataIn1 = 32'd2649
; 
32'd152468: dataIn1 = 32'd4714
; 
32'd152469: dataIn1 = 32'd4944
; 
32'd152470: dataIn1 = 32'd4955
; 
32'd152471: dataIn1 = 32'd4956
; 
32'd152472: dataIn1 = 32'd4957
; 
32'd152473: dataIn1 = 32'd2649
; 
32'd152474: dataIn1 = 32'd2651
; 
32'd152475: dataIn1 = 32'd4946
; 
32'd152476: dataIn1 = 32'd4955
; 
32'd152477: dataIn1 = 32'd4956
; 
32'd152478: dataIn1 = 32'd4957
; 
32'd152479: dataIn1 = 32'd4958
; 
32'd152480: dataIn1 = 32'd7847
; 
32'd152481: dataIn1 = 32'd2582
; 
32'd152482: dataIn1 = 32'd2651
; 
32'd152483: dataIn1 = 32'd4716
; 
32'd152484: dataIn1 = 32'd4955
; 
32'd152485: dataIn1 = 32'd4956
; 
32'd152486: dataIn1 = 32'd4957
; 
32'd152487: dataIn1 = 32'd4959
; 
32'd152488: dataIn1 = 32'd7857
; 
32'd152489: dataIn1 = 32'd4946
; 
32'd152490: dataIn1 = 32'd4956
; 
32'd152491: dataIn1 = 32'd4958
; 
32'd152492: dataIn1 = 32'd7843
; 
32'd152493: dataIn1 = 32'd7844
; 
32'd152494: dataIn1 = 32'd7846
; 
32'd152495: dataIn1 = 32'd7847
; 
32'd152496: dataIn1 = 32'd4716
; 
32'd152497: dataIn1 = 32'd4957
; 
32'd152498: dataIn1 = 32'd4959
; 
32'd152499: dataIn1 = 32'd7854
; 
32'd152500: dataIn1 = 32'd7855
; 
32'd152501: dataIn1 = 32'd7857
; 
32'd152502: dataIn1 = 32'd7859
; 
32'd152503: dataIn1 = 32'd2653
; 
32'd152504: dataIn1 = 32'd2654
; 
32'd152505: dataIn1 = 32'd4960
; 
32'd152506: dataIn1 = 32'd4961
; 
32'd152507: dataIn1 = 32'd4962
; 
32'd152508: dataIn1 = 32'd4963
; 
32'd152509: dataIn1 = 32'd4964
; 
32'd152510: dataIn1 = 32'd2652
; 
32'd152511: dataIn1 = 32'd2654
; 
32'd152512: dataIn1 = 32'd4960
; 
32'd152513: dataIn1 = 32'd4961
; 
32'd152514: dataIn1 = 32'd4962
; 
32'd152515: dataIn1 = 32'd4965
; 
32'd152516: dataIn1 = 32'd4966
; 
32'd152517: dataIn1 = 32'd2652
; 
32'd152518: dataIn1 = 32'd2653
; 
32'd152519: dataIn1 = 32'd4960
; 
32'd152520: dataIn1 = 32'd4961
; 
32'd152521: dataIn1 = 32'd4962
; 
32'd152522: dataIn1 = 32'd4967
; 
32'd152523: dataIn1 = 32'd4968
; 
32'd152524: dataIn1 = 32'd1085
; 
32'd152525: dataIn1 = 32'd2654
; 
32'd152526: dataIn1 = 32'd3511
; 
32'd152527: dataIn1 = 32'd4960
; 
32'd152528: dataIn1 = 32'd4963
; 
32'd152529: dataIn1 = 32'd4964
; 
32'd152530: dataIn1 = 32'd1085
; 
32'd152531: dataIn1 = 32'd2653
; 
32'd152532: dataIn1 = 32'd4719
; 
32'd152533: dataIn1 = 32'd4960
; 
32'd152534: dataIn1 = 32'd4963
; 
32'd152535: dataIn1 = 32'd4964
; 
32'd152536: dataIn1 = 32'd4974
; 
32'd152537: dataIn1 = 32'd1086
; 
32'd152538: dataIn1 = 32'd2654
; 
32'd152539: dataIn1 = 32'd3513
; 
32'd152540: dataIn1 = 32'd4961
; 
32'd152541: dataIn1 = 32'd4965
; 
32'd152542: dataIn1 = 32'd4966
; 
32'd152543: dataIn1 = 32'd1086
; 
32'd152544: dataIn1 = 32'd2652
; 
32'd152545: dataIn1 = 32'd4725
; 
32'd152546: dataIn1 = 32'd4961
; 
32'd152547: dataIn1 = 32'd4965
; 
32'd152548: dataIn1 = 32'd4966
; 
32'd152549: dataIn1 = 32'd4970
; 
32'd152550: dataIn1 = 32'd1111
; 
32'd152551: dataIn1 = 32'd2653
; 
32'd152552: dataIn1 = 32'd4962
; 
32'd152553: dataIn1 = 32'd4967
; 
32'd152554: dataIn1 = 32'd4968
; 
32'd152555: dataIn1 = 32'd4976
; 
32'd152556: dataIn1 = 32'd4978
; 
32'd152557: dataIn1 = 32'd7978
; 
32'd152558: dataIn1 = 32'd1111
; 
32'd152559: dataIn1 = 32'd2652
; 
32'd152560: dataIn1 = 32'd4962
; 
32'd152561: dataIn1 = 32'd4967
; 
32'd152562: dataIn1 = 32'd4968
; 
32'd152563: dataIn1 = 32'd4971
; 
32'd152564: dataIn1 = 32'd4973
; 
32'd152565: dataIn1 = 32'd8000
; 
32'd152566: dataIn1 = 32'd2585
; 
32'd152567: dataIn1 = 32'd2655
; 
32'd152568: dataIn1 = 32'd4723
; 
32'd152569: dataIn1 = 32'd4969
; 
32'd152570: dataIn1 = 32'd4970
; 
32'd152571: dataIn1 = 32'd4971
; 
32'd152572: dataIn1 = 32'd4972
; 
32'd152573: dataIn1 = 32'd7994
; 
32'd152574: dataIn1 = 32'd2585
; 
32'd152575: dataIn1 = 32'd2652
; 
32'd152576: dataIn1 = 32'd4725
; 
32'd152577: dataIn1 = 32'd4966
; 
32'd152578: dataIn1 = 32'd4969
; 
32'd152579: dataIn1 = 32'd4970
; 
32'd152580: dataIn1 = 32'd4971
; 
32'd152581: dataIn1 = 32'd2652
; 
32'd152582: dataIn1 = 32'd2655
; 
32'd152583: dataIn1 = 32'd4968
; 
32'd152584: dataIn1 = 32'd4969
; 
32'd152585: dataIn1 = 32'd4970
; 
32'd152586: dataIn1 = 32'd4971
; 
32'd152587: dataIn1 = 32'd4973
; 
32'd152588: dataIn1 = 32'd7999
; 
32'd152589: dataIn1 = 32'd4723
; 
32'd152590: dataIn1 = 32'd4969
; 
32'd152591: dataIn1 = 32'd4972
; 
32'd152592: dataIn1 = 32'd7991
; 
32'd152593: dataIn1 = 32'd7992
; 
32'd152594: dataIn1 = 32'd7994
; 
32'd152595: dataIn1 = 32'd7995
; 
32'd152596: dataIn1 = 32'd4968
; 
32'd152597: dataIn1 = 32'd4971
; 
32'd152598: dataIn1 = 32'd4973
; 
32'd152599: dataIn1 = 32'd7996
; 
32'd152600: dataIn1 = 32'd7998
; 
32'd152601: dataIn1 = 32'd7999
; 
32'd152602: dataIn1 = 32'd8000
; 
32'd152603: dataIn1 = 32'd2580
; 
32'd152604: dataIn1 = 32'd2653
; 
32'd152605: dataIn1 = 32'd4719
; 
32'd152606: dataIn1 = 32'd4964
; 
32'd152607: dataIn1 = 32'd4974
; 
32'd152608: dataIn1 = 32'd4975
; 
32'd152609: dataIn1 = 32'd4976
; 
32'd152610: dataIn1 = 32'd2580
; 
32'd152611: dataIn1 = 32'd2656
; 
32'd152612: dataIn1 = 32'd4717
; 
32'd152613: dataIn1 = 32'd4974
; 
32'd152614: dataIn1 = 32'd4975
; 
32'd152615: dataIn1 = 32'd4976
; 
32'd152616: dataIn1 = 32'd4977
; 
32'd152617: dataIn1 = 32'd7967
; 
32'd152618: dataIn1 = 32'd2653
; 
32'd152619: dataIn1 = 32'd2656
; 
32'd152620: dataIn1 = 32'd4967
; 
32'd152621: dataIn1 = 32'd4974
; 
32'd152622: dataIn1 = 32'd4975
; 
32'd152623: dataIn1 = 32'd4976
; 
32'd152624: dataIn1 = 32'd4978
; 
32'd152625: dataIn1 = 32'd7977
; 
32'd152626: dataIn1 = 32'd4717
; 
32'd152627: dataIn1 = 32'd4975
; 
32'd152628: dataIn1 = 32'd4977
; 
32'd152629: dataIn1 = 32'd7962
; 
32'd152630: dataIn1 = 32'd7963
; 
32'd152631: dataIn1 = 32'd7965
; 
32'd152632: dataIn1 = 32'd7967
; 
32'd152633: dataIn1 = 32'd4967
; 
32'd152634: dataIn1 = 32'd4976
; 
32'd152635: dataIn1 = 32'd4978
; 
32'd152636: dataIn1 = 32'd7975
; 
32'd152637: dataIn1 = 32'd7976
; 
32'd152638: dataIn1 = 32'd7977
; 
32'd152639: dataIn1 = 32'd7978
; 
32'd152640: dataIn1 = 32'd2658
; 
32'd152641: dataIn1 = 32'd2659
; 
32'd152642: dataIn1 = 32'd4979
; 
32'd152643: dataIn1 = 32'd4980
; 
32'd152644: dataIn1 = 32'd4981
; 
32'd152645: dataIn1 = 32'd4982
; 
32'd152646: dataIn1 = 32'd4983
; 
32'd152647: dataIn1 = 32'd2657
; 
32'd152648: dataIn1 = 32'd2659
; 
32'd152649: dataIn1 = 32'd4979
; 
32'd152650: dataIn1 = 32'd4980
; 
32'd152651: dataIn1 = 32'd4981
; 
32'd152652: dataIn1 = 32'd4984
; 
32'd152653: dataIn1 = 32'd4985
; 
32'd152654: dataIn1 = 32'd2657
; 
32'd152655: dataIn1 = 32'd2658
; 
32'd152656: dataIn1 = 32'd4979
; 
32'd152657: dataIn1 = 32'd4980
; 
32'd152658: dataIn1 = 32'd4981
; 
32'd152659: dataIn1 = 32'd4986
; 
32'd152660: dataIn1 = 32'd4987
; 
32'd152661: dataIn1 = 32'd1088
; 
32'd152662: dataIn1 = 32'd2659
; 
32'd152663: dataIn1 = 32'd4732
; 
32'd152664: dataIn1 = 32'd4979
; 
32'd152665: dataIn1 = 32'd4982
; 
32'd152666: dataIn1 = 32'd4983
; 
32'd152667: dataIn1 = 32'd4993
; 
32'd152668: dataIn1 = 32'd1088
; 
32'd152669: dataIn1 = 32'd2658
; 
32'd152670: dataIn1 = 32'd3521
; 
32'd152671: dataIn1 = 32'd4979
; 
32'd152672: dataIn1 = 32'd4982
; 
32'd152673: dataIn1 = 32'd4983
; 
32'd152674: dataIn1 = 32'd1112
; 
32'd152675: dataIn1 = 32'd2659
; 
32'd152676: dataIn1 = 32'd4980
; 
32'd152677: dataIn1 = 32'd4984
; 
32'd152678: dataIn1 = 32'd4985
; 
32'd152679: dataIn1 = 32'd4994
; 
32'd152680: dataIn1 = 32'd4996
; 
32'd152681: dataIn1 = 32'd8099
; 
32'd152682: dataIn1 = 32'd1112
; 
32'd152683: dataIn1 = 32'd2657
; 
32'd152684: dataIn1 = 32'd4980
; 
32'd152685: dataIn1 = 32'd4984
; 
32'd152686: dataIn1 = 32'd4985
; 
32'd152687: dataIn1 = 32'd4989
; 
32'd152688: dataIn1 = 32'd4992
; 
32'd152689: dataIn1 = 32'd8077
; 
32'd152690: dataIn1 = 32'd1087
; 
32'd152691: dataIn1 = 32'd2658
; 
32'd152692: dataIn1 = 32'd3519
; 
32'd152693: dataIn1 = 32'd4981
; 
32'd152694: dataIn1 = 32'd4986
; 
32'd152695: dataIn1 = 32'd4987
; 
32'd152696: dataIn1 = 32'd1087
; 
32'd152697: dataIn1 = 32'd2657
; 
32'd152698: dataIn1 = 32'd4727
; 
32'd152699: dataIn1 = 32'd4981
; 
32'd152700: dataIn1 = 32'd4986
; 
32'd152701: dataIn1 = 32'd4987
; 
32'd152702: dataIn1 = 32'd4990
; 
32'd152703: dataIn1 = 32'd2584
; 
32'd152704: dataIn1 = 32'd2660
; 
32'd152705: dataIn1 = 32'd4724
; 
32'd152706: dataIn1 = 32'd4988
; 
32'd152707: dataIn1 = 32'd4989
; 
32'd152708: dataIn1 = 32'd4990
; 
32'd152709: dataIn1 = 32'd4991
; 
32'd152710: dataIn1 = 32'd8083
; 
32'd152711: dataIn1 = 32'd2657
; 
32'd152712: dataIn1 = 32'd2660
; 
32'd152713: dataIn1 = 32'd4985
; 
32'd152714: dataIn1 = 32'd4988
; 
32'd152715: dataIn1 = 32'd4989
; 
32'd152716: dataIn1 = 32'd4990
; 
32'd152717: dataIn1 = 32'd4992
; 
32'd152718: dataIn1 = 32'd8078
; 
32'd152719: dataIn1 = 32'd2584
; 
32'd152720: dataIn1 = 32'd2657
; 
32'd152721: dataIn1 = 32'd4727
; 
32'd152722: dataIn1 = 32'd4987
; 
32'd152723: dataIn1 = 32'd4988
; 
32'd152724: dataIn1 = 32'd4989
; 
32'd152725: dataIn1 = 32'd4990
; 
32'd152726: dataIn1 = 32'd4724
; 
32'd152727: dataIn1 = 32'd4988
; 
32'd152728: dataIn1 = 32'd4991
; 
32'd152729: dataIn1 = 32'd8080
; 
32'd152730: dataIn1 = 32'd8081
; 
32'd152731: dataIn1 = 32'd8082
; 
32'd152732: dataIn1 = 32'd8083
; 
32'd152733: dataIn1 = 32'd4985
; 
32'd152734: dataIn1 = 32'd4989
; 
32'd152735: dataIn1 = 32'd4992
; 
32'd152736: dataIn1 = 32'd8074
; 
32'd152737: dataIn1 = 32'd8076
; 
32'd152738: dataIn1 = 32'd8077
; 
32'd152739: dataIn1 = 32'd8078
; 
32'd152740: dataIn1 = 32'd2588
; 
32'd152741: dataIn1 = 32'd2659
; 
32'd152742: dataIn1 = 32'd4732
; 
32'd152743: dataIn1 = 32'd4982
; 
32'd152744: dataIn1 = 32'd4993
; 
32'd152745: dataIn1 = 32'd4994
; 
32'd152746: dataIn1 = 32'd4995
; 
32'd152747: dataIn1 = 32'd2659
; 
32'd152748: dataIn1 = 32'd2661
; 
32'd152749: dataIn1 = 32'd4984
; 
32'd152750: dataIn1 = 32'd4993
; 
32'd152751: dataIn1 = 32'd4994
; 
32'd152752: dataIn1 = 32'd4995
; 
32'd152753: dataIn1 = 32'd4996
; 
32'd152754: dataIn1 = 32'd8100
; 
32'd152755: dataIn1 = 32'd2588
; 
32'd152756: dataIn1 = 32'd2661
; 
32'd152757: dataIn1 = 32'd4734
; 
32'd152758: dataIn1 = 32'd4993
; 
32'd152759: dataIn1 = 32'd4994
; 
32'd152760: dataIn1 = 32'd4995
; 
32'd152761: dataIn1 = 32'd4997
; 
32'd152762: dataIn1 = 32'd8110
; 
32'd152763: dataIn1 = 32'd4984
; 
32'd152764: dataIn1 = 32'd4994
; 
32'd152765: dataIn1 = 32'd4996
; 
32'd152766: dataIn1 = 32'd8096
; 
32'd152767: dataIn1 = 32'd8097
; 
32'd152768: dataIn1 = 32'd8099
; 
32'd152769: dataIn1 = 32'd8100
; 
32'd152770: dataIn1 = 32'd4734
; 
32'd152771: dataIn1 = 32'd4995
; 
32'd152772: dataIn1 = 32'd4997
; 
32'd152773: dataIn1 = 32'd8107
; 
32'd152774: dataIn1 = 32'd8108
; 
32'd152775: dataIn1 = 32'd8110
; 
32'd152776: dataIn1 = 32'd8112
; 
32'd152777: dataIn1 = 32'd2663
; 
32'd152778: dataIn1 = 32'd2664
; 
32'd152779: dataIn1 = 32'd4998
; 
32'd152780: dataIn1 = 32'd4999
; 
32'd152781: dataIn1 = 32'd5000
; 
32'd152782: dataIn1 = 32'd5001
; 
32'd152783: dataIn1 = 32'd5002
; 
32'd152784: dataIn1 = 32'd2662
; 
32'd152785: dataIn1 = 32'd2664
; 
32'd152786: dataIn1 = 32'd4998
; 
32'd152787: dataIn1 = 32'd4999
; 
32'd152788: dataIn1 = 32'd5000
; 
32'd152789: dataIn1 = 32'd5003
; 
32'd152790: dataIn1 = 32'd5004
; 
32'd152791: dataIn1 = 32'd2662
; 
32'd152792: dataIn1 = 32'd2663
; 
32'd152793: dataIn1 = 32'd4998
; 
32'd152794: dataIn1 = 32'd4999
; 
32'd152795: dataIn1 = 32'd5000
; 
32'd152796: dataIn1 = 32'd5005
; 
32'd152797: dataIn1 = 32'd5006
; 
32'd152798: dataIn1 = 32'd1089
; 
32'd152799: dataIn1 = 32'd2664
; 
32'd152800: dataIn1 = 32'd3527
; 
32'd152801: dataIn1 = 32'd4998
; 
32'd152802: dataIn1 = 32'd5001
; 
32'd152803: dataIn1 = 32'd5002
; 
32'd152804: dataIn1 = 32'd1089
; 
32'd152805: dataIn1 = 32'd2663
; 
32'd152806: dataIn1 = 32'd4737
; 
32'd152807: dataIn1 = 32'd4998
; 
32'd152808: dataIn1 = 32'd5001
; 
32'd152809: dataIn1 = 32'd5002
; 
32'd152810: dataIn1 = 32'd5012
; 
32'd152811: dataIn1 = 32'd1090
; 
32'd152812: dataIn1 = 32'd2664
; 
32'd152813: dataIn1 = 32'd3529
; 
32'd152814: dataIn1 = 32'd4999
; 
32'd152815: dataIn1 = 32'd5003
; 
32'd152816: dataIn1 = 32'd5004
; 
32'd152817: dataIn1 = 32'd1090
; 
32'd152818: dataIn1 = 32'd2662
; 
32'd152819: dataIn1 = 32'd4743
; 
32'd152820: dataIn1 = 32'd4999
; 
32'd152821: dataIn1 = 32'd5003
; 
32'd152822: dataIn1 = 32'd5004
; 
32'd152823: dataIn1 = 32'd5008
; 
32'd152824: dataIn1 = 32'd1113
; 
32'd152825: dataIn1 = 32'd2663
; 
32'd152826: dataIn1 = 32'd5000
; 
32'd152827: dataIn1 = 32'd5005
; 
32'd152828: dataIn1 = 32'd5006
; 
32'd152829: dataIn1 = 32'd5014
; 
32'd152830: dataIn1 = 32'd5016
; 
32'd152831: dataIn1 = 32'd8231
; 
32'd152832: dataIn1 = 32'd1113
; 
32'd152833: dataIn1 = 32'd2662
; 
32'd152834: dataIn1 = 32'd5000
; 
32'd152835: dataIn1 = 32'd5005
; 
32'd152836: dataIn1 = 32'd5006
; 
32'd152837: dataIn1 = 32'd5009
; 
32'd152838: dataIn1 = 32'd5011
; 
32'd152839: dataIn1 = 32'd8253
; 
32'd152840: dataIn1 = 32'd2591
; 
32'd152841: dataIn1 = 32'd2665
; 
32'd152842: dataIn1 = 32'd4741
; 
32'd152843: dataIn1 = 32'd5007
; 
32'd152844: dataIn1 = 32'd5008
; 
32'd152845: dataIn1 = 32'd5009
; 
32'd152846: dataIn1 = 32'd5010
; 
32'd152847: dataIn1 = 32'd8247
; 
32'd152848: dataIn1 = 32'd2591
; 
32'd152849: dataIn1 = 32'd2662
; 
32'd152850: dataIn1 = 32'd4743
; 
32'd152851: dataIn1 = 32'd5004
; 
32'd152852: dataIn1 = 32'd5007
; 
32'd152853: dataIn1 = 32'd5008
; 
32'd152854: dataIn1 = 32'd5009
; 
32'd152855: dataIn1 = 32'd2662
; 
32'd152856: dataIn1 = 32'd2665
; 
32'd152857: dataIn1 = 32'd5006
; 
32'd152858: dataIn1 = 32'd5007
; 
32'd152859: dataIn1 = 32'd5008
; 
32'd152860: dataIn1 = 32'd5009
; 
32'd152861: dataIn1 = 32'd5011
; 
32'd152862: dataIn1 = 32'd8252
; 
32'd152863: dataIn1 = 32'd4741
; 
32'd152864: dataIn1 = 32'd5007
; 
32'd152865: dataIn1 = 32'd5010
; 
32'd152866: dataIn1 = 32'd8244
; 
32'd152867: dataIn1 = 32'd8245
; 
32'd152868: dataIn1 = 32'd8247
; 
32'd152869: dataIn1 = 32'd8248
; 
32'd152870: dataIn1 = 32'd5006
; 
32'd152871: dataIn1 = 32'd5009
; 
32'd152872: dataIn1 = 32'd5011
; 
32'd152873: dataIn1 = 32'd8249
; 
32'd152874: dataIn1 = 32'd8251
; 
32'd152875: dataIn1 = 32'd8252
; 
32'd152876: dataIn1 = 32'd8253
; 
32'd152877: dataIn1 = 32'd2586
; 
32'd152878: dataIn1 = 32'd2663
; 
32'd152879: dataIn1 = 32'd4737
; 
32'd152880: dataIn1 = 32'd5002
; 
32'd152881: dataIn1 = 32'd5012
; 
32'd152882: dataIn1 = 32'd5013
; 
32'd152883: dataIn1 = 32'd5014
; 
32'd152884: dataIn1 = 32'd2586
; 
32'd152885: dataIn1 = 32'd2666
; 
32'd152886: dataIn1 = 32'd4735
; 
32'd152887: dataIn1 = 32'd5012
; 
32'd152888: dataIn1 = 32'd5013
; 
32'd152889: dataIn1 = 32'd5014
; 
32'd152890: dataIn1 = 32'd5015
; 
32'd152891: dataIn1 = 32'd8220
; 
32'd152892: dataIn1 = 32'd2663
; 
32'd152893: dataIn1 = 32'd2666
; 
32'd152894: dataIn1 = 32'd5005
; 
32'd152895: dataIn1 = 32'd5012
; 
32'd152896: dataIn1 = 32'd5013
; 
32'd152897: dataIn1 = 32'd5014
; 
32'd152898: dataIn1 = 32'd5016
; 
32'd152899: dataIn1 = 32'd8230
; 
32'd152900: dataIn1 = 32'd4735
; 
32'd152901: dataIn1 = 32'd5013
; 
32'd152902: dataIn1 = 32'd5015
; 
32'd152903: dataIn1 = 32'd8215
; 
32'd152904: dataIn1 = 32'd8216
; 
32'd152905: dataIn1 = 32'd8218
; 
32'd152906: dataIn1 = 32'd8220
; 
32'd152907: dataIn1 = 32'd5005
; 
32'd152908: dataIn1 = 32'd5014
; 
32'd152909: dataIn1 = 32'd5016
; 
32'd152910: dataIn1 = 32'd8228
; 
32'd152911: dataIn1 = 32'd8229
; 
32'd152912: dataIn1 = 32'd8230
; 
32'd152913: dataIn1 = 32'd8231
; 
32'd152914: dataIn1 = 32'd2668
; 
32'd152915: dataIn1 = 32'd2669
; 
32'd152916: dataIn1 = 32'd5017
; 
32'd152917: dataIn1 = 32'd5018
; 
32'd152918: dataIn1 = 32'd5019
; 
32'd152919: dataIn1 = 32'd5020
; 
32'd152920: dataIn1 = 32'd5021
; 
32'd152921: dataIn1 = 32'd2667
; 
32'd152922: dataIn1 = 32'd2669
; 
32'd152923: dataIn1 = 32'd5017
; 
32'd152924: dataIn1 = 32'd5018
; 
32'd152925: dataIn1 = 32'd5019
; 
32'd152926: dataIn1 = 32'd5022
; 
32'd152927: dataIn1 = 32'd5023
; 
32'd152928: dataIn1 = 32'd2667
; 
32'd152929: dataIn1 = 32'd2668
; 
32'd152930: dataIn1 = 32'd5017
; 
32'd152931: dataIn1 = 32'd5018
; 
32'd152932: dataIn1 = 32'd5019
; 
32'd152933: dataIn1 = 32'd5024
; 
32'd152934: dataIn1 = 32'd5025
; 
32'd152935: dataIn1 = 32'd1092
; 
32'd152936: dataIn1 = 32'd2669
; 
32'd152937: dataIn1 = 32'd4750
; 
32'd152938: dataIn1 = 32'd5017
; 
32'd152939: dataIn1 = 32'd5020
; 
32'd152940: dataIn1 = 32'd5021
; 
32'd152941: dataIn1 = 32'd5031
; 
32'd152942: dataIn1 = 32'd1092
; 
32'd152943: dataIn1 = 32'd2668
; 
32'd152944: dataIn1 = 32'd3537
; 
32'd152945: dataIn1 = 32'd5017
; 
32'd152946: dataIn1 = 32'd5020
; 
32'd152947: dataIn1 = 32'd5021
; 
32'd152948: dataIn1 = 32'd1114
; 
32'd152949: dataIn1 = 32'd2669
; 
32'd152950: dataIn1 = 32'd5018
; 
32'd152951: dataIn1 = 32'd5022
; 
32'd152952: dataIn1 = 32'd5023
; 
32'd152953: dataIn1 = 32'd5032
; 
32'd152954: dataIn1 = 32'd5034
; 
32'd152955: dataIn1 = 32'd8351
; 
32'd152956: dataIn1 = 32'd1114
; 
32'd152957: dataIn1 = 32'd2667
; 
32'd152958: dataIn1 = 32'd5018
; 
32'd152959: dataIn1 = 32'd5022
; 
32'd152960: dataIn1 = 32'd5023
; 
32'd152961: dataIn1 = 32'd5027
; 
32'd152962: dataIn1 = 32'd5030
; 
32'd152963: dataIn1 = 32'd8329
; 
32'd152964: dataIn1 = 32'd1091
; 
32'd152965: dataIn1 = 32'd2668
; 
32'd152966: dataIn1 = 32'd3535
; 
32'd152967: dataIn1 = 32'd5019
; 
32'd152968: dataIn1 = 32'd5024
; 
32'd152969: dataIn1 = 32'd5025
; 
32'd152970: dataIn1 = 32'd1091
; 
32'd152971: dataIn1 = 32'd2667
; 
32'd152972: dataIn1 = 32'd4745
; 
32'd152973: dataIn1 = 32'd5019
; 
32'd152974: dataIn1 = 32'd5024
; 
32'd152975: dataIn1 = 32'd5025
; 
32'd152976: dataIn1 = 32'd5028
; 
32'd152977: dataIn1 = 32'd2590
; 
32'd152978: dataIn1 = 32'd2670
; 
32'd152979: dataIn1 = 32'd4742
; 
32'd152980: dataIn1 = 32'd5026
; 
32'd152981: dataIn1 = 32'd5027
; 
32'd152982: dataIn1 = 32'd5028
; 
32'd152983: dataIn1 = 32'd5029
; 
32'd152984: dataIn1 = 32'd8335
; 
32'd152985: dataIn1 = 32'd2667
; 
32'd152986: dataIn1 = 32'd2670
; 
32'd152987: dataIn1 = 32'd5023
; 
32'd152988: dataIn1 = 32'd5026
; 
32'd152989: dataIn1 = 32'd5027
; 
32'd152990: dataIn1 = 32'd5028
; 
32'd152991: dataIn1 = 32'd5030
; 
32'd152992: dataIn1 = 32'd8330
; 
32'd152993: dataIn1 = 32'd2590
; 
32'd152994: dataIn1 = 32'd2667
; 
32'd152995: dataIn1 = 32'd4745
; 
32'd152996: dataIn1 = 32'd5025
; 
32'd152997: dataIn1 = 32'd5026
; 
32'd152998: dataIn1 = 32'd5027
; 
32'd152999: dataIn1 = 32'd5028
; 
32'd153000: dataIn1 = 32'd4742
; 
32'd153001: dataIn1 = 32'd5026
; 
32'd153002: dataIn1 = 32'd5029
; 
32'd153003: dataIn1 = 32'd8332
; 
32'd153004: dataIn1 = 32'd8333
; 
32'd153005: dataIn1 = 32'd8334
; 
32'd153006: dataIn1 = 32'd8335
; 
32'd153007: dataIn1 = 32'd5023
; 
32'd153008: dataIn1 = 32'd5027
; 
32'd153009: dataIn1 = 32'd5030
; 
32'd153010: dataIn1 = 32'd8326
; 
32'd153011: dataIn1 = 32'd8328
; 
32'd153012: dataIn1 = 32'd8329
; 
32'd153013: dataIn1 = 32'd8330
; 
32'd153014: dataIn1 = 32'd2594
; 
32'd153015: dataIn1 = 32'd2669
; 
32'd153016: dataIn1 = 32'd4750
; 
32'd153017: dataIn1 = 32'd5020
; 
32'd153018: dataIn1 = 32'd5031
; 
32'd153019: dataIn1 = 32'd5032
; 
32'd153020: dataIn1 = 32'd5033
; 
32'd153021: dataIn1 = 32'd2669
; 
32'd153022: dataIn1 = 32'd2671
; 
32'd153023: dataIn1 = 32'd5022
; 
32'd153024: dataIn1 = 32'd5031
; 
32'd153025: dataIn1 = 32'd5032
; 
32'd153026: dataIn1 = 32'd5033
; 
32'd153027: dataIn1 = 32'd5034
; 
32'd153028: dataIn1 = 32'd8352
; 
32'd153029: dataIn1 = 32'd2594
; 
32'd153030: dataIn1 = 32'd2671
; 
32'd153031: dataIn1 = 32'd4752
; 
32'd153032: dataIn1 = 32'd5031
; 
32'd153033: dataIn1 = 32'd5032
; 
32'd153034: dataIn1 = 32'd5033
; 
32'd153035: dataIn1 = 32'd5035
; 
32'd153036: dataIn1 = 32'd8362
; 
32'd153037: dataIn1 = 32'd5022
; 
32'd153038: dataIn1 = 32'd5032
; 
32'd153039: dataIn1 = 32'd5034
; 
32'd153040: dataIn1 = 32'd8348
; 
32'd153041: dataIn1 = 32'd8349
; 
32'd153042: dataIn1 = 32'd8351
; 
32'd153043: dataIn1 = 32'd8352
; 
32'd153044: dataIn1 = 32'd4752
; 
32'd153045: dataIn1 = 32'd5033
; 
32'd153046: dataIn1 = 32'd5035
; 
32'd153047: dataIn1 = 32'd8359
; 
32'd153048: dataIn1 = 32'd8360
; 
32'd153049: dataIn1 = 32'd8362
; 
32'd153050: dataIn1 = 32'd8364
; 
32'd153051: dataIn1 = 32'd2673
; 
32'd153052: dataIn1 = 32'd2674
; 
32'd153053: dataIn1 = 32'd5036
; 
32'd153054: dataIn1 = 32'd5037
; 
32'd153055: dataIn1 = 32'd5038
; 
32'd153056: dataIn1 = 32'd5039
; 
32'd153057: dataIn1 = 32'd5040
; 
32'd153058: dataIn1 = 32'd2672
; 
32'd153059: dataIn1 = 32'd2674
; 
32'd153060: dataIn1 = 32'd5036
; 
32'd153061: dataIn1 = 32'd5037
; 
32'd153062: dataIn1 = 32'd5038
; 
32'd153063: dataIn1 = 32'd5041
; 
32'd153064: dataIn1 = 32'd5042
; 
32'd153065: dataIn1 = 32'd2672
; 
32'd153066: dataIn1 = 32'd2673
; 
32'd153067: dataIn1 = 32'd5036
; 
32'd153068: dataIn1 = 32'd5037
; 
32'd153069: dataIn1 = 32'd5038
; 
32'd153070: dataIn1 = 32'd5043
; 
32'd153071: dataIn1 = 32'd5044
; 
32'd153072: dataIn1 = 32'd1093
; 
32'd153073: dataIn1 = 32'd2674
; 
32'd153074: dataIn1 = 32'd3543
; 
32'd153075: dataIn1 = 32'd5036
; 
32'd153076: dataIn1 = 32'd5039
; 
32'd153077: dataIn1 = 32'd5040
; 
32'd153078: dataIn1 = 32'd1093
; 
32'd153079: dataIn1 = 32'd2673
; 
32'd153080: dataIn1 = 32'd4755
; 
32'd153081: dataIn1 = 32'd5036
; 
32'd153082: dataIn1 = 32'd5039
; 
32'd153083: dataIn1 = 32'd5040
; 
32'd153084: dataIn1 = 32'd5050
; 
32'd153085: dataIn1 = 32'd1094
; 
32'd153086: dataIn1 = 32'd2674
; 
32'd153087: dataIn1 = 32'd3545
; 
32'd153088: dataIn1 = 32'd5037
; 
32'd153089: dataIn1 = 32'd5041
; 
32'd153090: dataIn1 = 32'd5042
; 
32'd153091: dataIn1 = 32'd1094
; 
32'd153092: dataIn1 = 32'd2672
; 
32'd153093: dataIn1 = 32'd4761
; 
32'd153094: dataIn1 = 32'd5037
; 
32'd153095: dataIn1 = 32'd5041
; 
32'd153096: dataIn1 = 32'd5042
; 
32'd153097: dataIn1 = 32'd5046
; 
32'd153098: dataIn1 = 32'd1115
; 
32'd153099: dataIn1 = 32'd2673
; 
32'd153100: dataIn1 = 32'd5038
; 
32'd153101: dataIn1 = 32'd5043
; 
32'd153102: dataIn1 = 32'd5044
; 
32'd153103: dataIn1 = 32'd5052
; 
32'd153104: dataIn1 = 32'd5054
; 
32'd153105: dataIn1 = 32'd8483
; 
32'd153106: dataIn1 = 32'd1115
; 
32'd153107: dataIn1 = 32'd2672
; 
32'd153108: dataIn1 = 32'd5038
; 
32'd153109: dataIn1 = 32'd5043
; 
32'd153110: dataIn1 = 32'd5044
; 
32'd153111: dataIn1 = 32'd5047
; 
32'd153112: dataIn1 = 32'd5049
; 
32'd153113: dataIn1 = 32'd8505
; 
32'd153114: dataIn1 = 32'd2597
; 
32'd153115: dataIn1 = 32'd2675
; 
32'd153116: dataIn1 = 32'd4759
; 
32'd153117: dataIn1 = 32'd5045
; 
32'd153118: dataIn1 = 32'd5046
; 
32'd153119: dataIn1 = 32'd5047
; 
32'd153120: dataIn1 = 32'd5048
; 
32'd153121: dataIn1 = 32'd8499
; 
32'd153122: dataIn1 = 32'd2597
; 
32'd153123: dataIn1 = 32'd2672
; 
32'd153124: dataIn1 = 32'd4761
; 
32'd153125: dataIn1 = 32'd5042
; 
32'd153126: dataIn1 = 32'd5045
; 
32'd153127: dataIn1 = 32'd5046
; 
32'd153128: dataIn1 = 32'd5047
; 
32'd153129: dataIn1 = 32'd2672
; 
32'd153130: dataIn1 = 32'd2675
; 
32'd153131: dataIn1 = 32'd5044
; 
32'd153132: dataIn1 = 32'd5045
; 
32'd153133: dataIn1 = 32'd5046
; 
32'd153134: dataIn1 = 32'd5047
; 
32'd153135: dataIn1 = 32'd5049
; 
32'd153136: dataIn1 = 32'd8504
; 
32'd153137: dataIn1 = 32'd4759
; 
32'd153138: dataIn1 = 32'd5045
; 
32'd153139: dataIn1 = 32'd5048
; 
32'd153140: dataIn1 = 32'd8496
; 
32'd153141: dataIn1 = 32'd8497
; 
32'd153142: dataIn1 = 32'd8499
; 
32'd153143: dataIn1 = 32'd8500
; 
32'd153144: dataIn1 = 32'd5044
; 
32'd153145: dataIn1 = 32'd5047
; 
32'd153146: dataIn1 = 32'd5049
; 
32'd153147: dataIn1 = 32'd8501
; 
32'd153148: dataIn1 = 32'd8503
; 
32'd153149: dataIn1 = 32'd8504
; 
32'd153150: dataIn1 = 32'd8505
; 
32'd153151: dataIn1 = 32'd2592
; 
32'd153152: dataIn1 = 32'd2673
; 
32'd153153: dataIn1 = 32'd4755
; 
32'd153154: dataIn1 = 32'd5040
; 
32'd153155: dataIn1 = 32'd5050
; 
32'd153156: dataIn1 = 32'd5051
; 
32'd153157: dataIn1 = 32'd5052
; 
32'd153158: dataIn1 = 32'd2592
; 
32'd153159: dataIn1 = 32'd2676
; 
32'd153160: dataIn1 = 32'd4753
; 
32'd153161: dataIn1 = 32'd5050
; 
32'd153162: dataIn1 = 32'd5051
; 
32'd153163: dataIn1 = 32'd5052
; 
32'd153164: dataIn1 = 32'd5053
; 
32'd153165: dataIn1 = 32'd8472
; 
32'd153166: dataIn1 = 32'd2673
; 
32'd153167: dataIn1 = 32'd2676
; 
32'd153168: dataIn1 = 32'd5043
; 
32'd153169: dataIn1 = 32'd5050
; 
32'd153170: dataIn1 = 32'd5051
; 
32'd153171: dataIn1 = 32'd5052
; 
32'd153172: dataIn1 = 32'd5054
; 
32'd153173: dataIn1 = 32'd8482
; 
32'd153174: dataIn1 = 32'd4753
; 
32'd153175: dataIn1 = 32'd5051
; 
32'd153176: dataIn1 = 32'd5053
; 
32'd153177: dataIn1 = 32'd8467
; 
32'd153178: dataIn1 = 32'd8468
; 
32'd153179: dataIn1 = 32'd8470
; 
32'd153180: dataIn1 = 32'd8472
; 
32'd153181: dataIn1 = 32'd5043
; 
32'd153182: dataIn1 = 32'd5052
; 
32'd153183: dataIn1 = 32'd5054
; 
32'd153184: dataIn1 = 32'd8480
; 
32'd153185: dataIn1 = 32'd8481
; 
32'd153186: dataIn1 = 32'd8482
; 
32'd153187: dataIn1 = 32'd8483
; 
32'd153188: dataIn1 = 32'd2678
; 
32'd153189: dataIn1 = 32'd2679
; 
32'd153190: dataIn1 = 32'd5055
; 
32'd153191: dataIn1 = 32'd5056
; 
32'd153192: dataIn1 = 32'd5057
; 
32'd153193: dataIn1 = 32'd5058
; 
32'd153194: dataIn1 = 32'd5059
; 
32'd153195: dataIn1 = 32'd2677
; 
32'd153196: dataIn1 = 32'd2679
; 
32'd153197: dataIn1 = 32'd5055
; 
32'd153198: dataIn1 = 32'd5056
; 
32'd153199: dataIn1 = 32'd5057
; 
32'd153200: dataIn1 = 32'd5060
; 
32'd153201: dataIn1 = 32'd5061
; 
32'd153202: dataIn1 = 32'd2677
; 
32'd153203: dataIn1 = 32'd2678
; 
32'd153204: dataIn1 = 32'd5055
; 
32'd153205: dataIn1 = 32'd5056
; 
32'd153206: dataIn1 = 32'd5057
; 
32'd153207: dataIn1 = 32'd5062
; 
32'd153208: dataIn1 = 32'd5063
; 
32'd153209: dataIn1 = 32'd1096
; 
32'd153210: dataIn1 = 32'd2679
; 
32'd153211: dataIn1 = 32'd4768
; 
32'd153212: dataIn1 = 32'd5055
; 
32'd153213: dataIn1 = 32'd5058
; 
32'd153214: dataIn1 = 32'd5059
; 
32'd153215: dataIn1 = 32'd5069
; 
32'd153216: dataIn1 = 32'd1096
; 
32'd153217: dataIn1 = 32'd2678
; 
32'd153218: dataIn1 = 32'd3553
; 
32'd153219: dataIn1 = 32'd5055
; 
32'd153220: dataIn1 = 32'd5058
; 
32'd153221: dataIn1 = 32'd5059
; 
32'd153222: dataIn1 = 32'd1116
; 
32'd153223: dataIn1 = 32'd2679
; 
32'd153224: dataIn1 = 32'd5056
; 
32'd153225: dataIn1 = 32'd5060
; 
32'd153226: dataIn1 = 32'd5061
; 
32'd153227: dataIn1 = 32'd5070
; 
32'd153228: dataIn1 = 32'd5072
; 
32'd153229: dataIn1 = 32'd8604
; 
32'd153230: dataIn1 = 32'd1116
; 
32'd153231: dataIn1 = 32'd2677
; 
32'd153232: dataIn1 = 32'd5056
; 
32'd153233: dataIn1 = 32'd5060
; 
32'd153234: dataIn1 = 32'd5061
; 
32'd153235: dataIn1 = 32'd5065
; 
32'd153236: dataIn1 = 32'd5068
; 
32'd153237: dataIn1 = 32'd8582
; 
32'd153238: dataIn1 = 32'd1095
; 
32'd153239: dataIn1 = 32'd2678
; 
32'd153240: dataIn1 = 32'd3551
; 
32'd153241: dataIn1 = 32'd5057
; 
32'd153242: dataIn1 = 32'd5062
; 
32'd153243: dataIn1 = 32'd5063
; 
32'd153244: dataIn1 = 32'd1095
; 
32'd153245: dataIn1 = 32'd2677
; 
32'd153246: dataIn1 = 32'd4763
; 
32'd153247: dataIn1 = 32'd5057
; 
32'd153248: dataIn1 = 32'd5062
; 
32'd153249: dataIn1 = 32'd5063
; 
32'd153250: dataIn1 = 32'd5066
; 
32'd153251: dataIn1 = 32'd2596
; 
32'd153252: dataIn1 = 32'd2680
; 
32'd153253: dataIn1 = 32'd4760
; 
32'd153254: dataIn1 = 32'd5064
; 
32'd153255: dataIn1 = 32'd5065
; 
32'd153256: dataIn1 = 32'd5066
; 
32'd153257: dataIn1 = 32'd5067
; 
32'd153258: dataIn1 = 32'd8588
; 
32'd153259: dataIn1 = 32'd2677
; 
32'd153260: dataIn1 = 32'd2680
; 
32'd153261: dataIn1 = 32'd5061
; 
32'd153262: dataIn1 = 32'd5064
; 
32'd153263: dataIn1 = 32'd5065
; 
32'd153264: dataIn1 = 32'd5066
; 
32'd153265: dataIn1 = 32'd5068
; 
32'd153266: dataIn1 = 32'd8583
; 
32'd153267: dataIn1 = 32'd2596
; 
32'd153268: dataIn1 = 32'd2677
; 
32'd153269: dataIn1 = 32'd4763
; 
32'd153270: dataIn1 = 32'd5063
; 
32'd153271: dataIn1 = 32'd5064
; 
32'd153272: dataIn1 = 32'd5065
; 
32'd153273: dataIn1 = 32'd5066
; 
32'd153274: dataIn1 = 32'd4760
; 
32'd153275: dataIn1 = 32'd5064
; 
32'd153276: dataIn1 = 32'd5067
; 
32'd153277: dataIn1 = 32'd8585
; 
32'd153278: dataIn1 = 32'd8586
; 
32'd153279: dataIn1 = 32'd8587
; 
32'd153280: dataIn1 = 32'd8588
; 
32'd153281: dataIn1 = 32'd5061
; 
32'd153282: dataIn1 = 32'd5065
; 
32'd153283: dataIn1 = 32'd5068
; 
32'd153284: dataIn1 = 32'd8579
; 
32'd153285: dataIn1 = 32'd8581
; 
32'd153286: dataIn1 = 32'd8582
; 
32'd153287: dataIn1 = 32'd8583
; 
32'd153288: dataIn1 = 32'd2600
; 
32'd153289: dataIn1 = 32'd2679
; 
32'd153290: dataIn1 = 32'd4768
; 
32'd153291: dataIn1 = 32'd5058
; 
32'd153292: dataIn1 = 32'd5069
; 
32'd153293: dataIn1 = 32'd5070
; 
32'd153294: dataIn1 = 32'd5071
; 
32'd153295: dataIn1 = 32'd2679
; 
32'd153296: dataIn1 = 32'd2681
; 
32'd153297: dataIn1 = 32'd5060
; 
32'd153298: dataIn1 = 32'd5069
; 
32'd153299: dataIn1 = 32'd5070
; 
32'd153300: dataIn1 = 32'd5071
; 
32'd153301: dataIn1 = 32'd5072
; 
32'd153302: dataIn1 = 32'd8605
; 
32'd153303: dataIn1 = 32'd2600
; 
32'd153304: dataIn1 = 32'd2681
; 
32'd153305: dataIn1 = 32'd4770
; 
32'd153306: dataIn1 = 32'd5069
; 
32'd153307: dataIn1 = 32'd5070
; 
32'd153308: dataIn1 = 32'd5071
; 
32'd153309: dataIn1 = 32'd5073
; 
32'd153310: dataIn1 = 32'd8615
; 
32'd153311: dataIn1 = 32'd5060
; 
32'd153312: dataIn1 = 32'd5070
; 
32'd153313: dataIn1 = 32'd5072
; 
32'd153314: dataIn1 = 32'd8601
; 
32'd153315: dataIn1 = 32'd8602
; 
32'd153316: dataIn1 = 32'd8604
; 
32'd153317: dataIn1 = 32'd8605
; 
32'd153318: dataIn1 = 32'd4770
; 
32'd153319: dataIn1 = 32'd5071
; 
32'd153320: dataIn1 = 32'd5073
; 
32'd153321: dataIn1 = 32'd8612
; 
32'd153322: dataIn1 = 32'd8613
; 
32'd153323: dataIn1 = 32'd8615
; 
32'd153324: dataIn1 = 32'd8617
; 
32'd153325: dataIn1 = 32'd2683
; 
32'd153326: dataIn1 = 32'd2684
; 
32'd153327: dataIn1 = 32'd5074
; 
32'd153328: dataIn1 = 32'd5075
; 
32'd153329: dataIn1 = 32'd5076
; 
32'd153330: dataIn1 = 32'd5077
; 
32'd153331: dataIn1 = 32'd5078
; 
32'd153332: dataIn1 = 32'd2682
; 
32'd153333: dataIn1 = 32'd2684
; 
32'd153334: dataIn1 = 32'd5074
; 
32'd153335: dataIn1 = 32'd5075
; 
32'd153336: dataIn1 = 32'd5076
; 
32'd153337: dataIn1 = 32'd5079
; 
32'd153338: dataIn1 = 32'd5080
; 
32'd153339: dataIn1 = 32'd2682
; 
32'd153340: dataIn1 = 32'd2683
; 
32'd153341: dataIn1 = 32'd5074
; 
32'd153342: dataIn1 = 32'd5075
; 
32'd153343: dataIn1 = 32'd5076
; 
32'd153344: dataIn1 = 32'd5081
; 
32'd153345: dataIn1 = 32'd5082
; 
32'd153346: dataIn1 = 32'd1097
; 
32'd153347: dataIn1 = 32'd2684
; 
32'd153348: dataIn1 = 32'd3559
; 
32'd153349: dataIn1 = 32'd5074
; 
32'd153350: dataIn1 = 32'd5077
; 
32'd153351: dataIn1 = 32'd5078
; 
32'd153352: dataIn1 = 32'd1097
; 
32'd153353: dataIn1 = 32'd2683
; 
32'd153354: dataIn1 = 32'd4773
; 
32'd153355: dataIn1 = 32'd5074
; 
32'd153356: dataIn1 = 32'd5077
; 
32'd153357: dataIn1 = 32'd5078
; 
32'd153358: dataIn1 = 32'd5088
; 
32'd153359: dataIn1 = 32'd1098
; 
32'd153360: dataIn1 = 32'd2684
; 
32'd153361: dataIn1 = 32'd3561
; 
32'd153362: dataIn1 = 32'd5075
; 
32'd153363: dataIn1 = 32'd5079
; 
32'd153364: dataIn1 = 32'd5080
; 
32'd153365: dataIn1 = 32'd1098
; 
32'd153366: dataIn1 = 32'd2682
; 
32'd153367: dataIn1 = 32'd4779
; 
32'd153368: dataIn1 = 32'd5075
; 
32'd153369: dataIn1 = 32'd5079
; 
32'd153370: dataIn1 = 32'd5080
; 
32'd153371: dataIn1 = 32'd5084
; 
32'd153372: dataIn1 = 32'd1117
; 
32'd153373: dataIn1 = 32'd2683
; 
32'd153374: dataIn1 = 32'd5076
; 
32'd153375: dataIn1 = 32'd5081
; 
32'd153376: dataIn1 = 32'd5082
; 
32'd153377: dataIn1 = 32'd5090
; 
32'd153378: dataIn1 = 32'd5092
; 
32'd153379: dataIn1 = 32'd8736
; 
32'd153380: dataIn1 = 32'd1117
; 
32'd153381: dataIn1 = 32'd2682
; 
32'd153382: dataIn1 = 32'd5076
; 
32'd153383: dataIn1 = 32'd5081
; 
32'd153384: dataIn1 = 32'd5082
; 
32'd153385: dataIn1 = 32'd5085
; 
32'd153386: dataIn1 = 32'd5087
; 
32'd153387: dataIn1 = 32'd8758
; 
32'd153388: dataIn1 = 32'd2603
; 
32'd153389: dataIn1 = 32'd2685
; 
32'd153390: dataIn1 = 32'd4777
; 
32'd153391: dataIn1 = 32'd5083
; 
32'd153392: dataIn1 = 32'd5084
; 
32'd153393: dataIn1 = 32'd5085
; 
32'd153394: dataIn1 = 32'd5086
; 
32'd153395: dataIn1 = 32'd8752
; 
32'd153396: dataIn1 = 32'd2603
; 
32'd153397: dataIn1 = 32'd2682
; 
32'd153398: dataIn1 = 32'd4779
; 
32'd153399: dataIn1 = 32'd5080
; 
32'd153400: dataIn1 = 32'd5083
; 
32'd153401: dataIn1 = 32'd5084
; 
32'd153402: dataIn1 = 32'd5085
; 
32'd153403: dataIn1 = 32'd2682
; 
32'd153404: dataIn1 = 32'd2685
; 
32'd153405: dataIn1 = 32'd5082
; 
32'd153406: dataIn1 = 32'd5083
; 
32'd153407: dataIn1 = 32'd5084
; 
32'd153408: dataIn1 = 32'd5085
; 
32'd153409: dataIn1 = 32'd5087
; 
32'd153410: dataIn1 = 32'd8757
; 
32'd153411: dataIn1 = 32'd4777
; 
32'd153412: dataIn1 = 32'd5083
; 
32'd153413: dataIn1 = 32'd5086
; 
32'd153414: dataIn1 = 32'd8749
; 
32'd153415: dataIn1 = 32'd8750
; 
32'd153416: dataIn1 = 32'd8752
; 
32'd153417: dataIn1 = 32'd8753
; 
32'd153418: dataIn1 = 32'd5082
; 
32'd153419: dataIn1 = 32'd5085
; 
32'd153420: dataIn1 = 32'd5087
; 
32'd153421: dataIn1 = 32'd8754
; 
32'd153422: dataIn1 = 32'd8756
; 
32'd153423: dataIn1 = 32'd8757
; 
32'd153424: dataIn1 = 32'd8758
; 
32'd153425: dataIn1 = 32'd2598
; 
32'd153426: dataIn1 = 32'd2683
; 
32'd153427: dataIn1 = 32'd4773
; 
32'd153428: dataIn1 = 32'd5078
; 
32'd153429: dataIn1 = 32'd5088
; 
32'd153430: dataIn1 = 32'd5089
; 
32'd153431: dataIn1 = 32'd5090
; 
32'd153432: dataIn1 = 32'd2598
; 
32'd153433: dataIn1 = 32'd2686
; 
32'd153434: dataIn1 = 32'd4771
; 
32'd153435: dataIn1 = 32'd5088
; 
32'd153436: dataIn1 = 32'd5089
; 
32'd153437: dataIn1 = 32'd5090
; 
32'd153438: dataIn1 = 32'd5091
; 
32'd153439: dataIn1 = 32'd8725
; 
32'd153440: dataIn1 = 32'd2683
; 
32'd153441: dataIn1 = 32'd2686
; 
32'd153442: dataIn1 = 32'd5081
; 
32'd153443: dataIn1 = 32'd5088
; 
32'd153444: dataIn1 = 32'd5089
; 
32'd153445: dataIn1 = 32'd5090
; 
32'd153446: dataIn1 = 32'd5092
; 
32'd153447: dataIn1 = 32'd8735
; 
32'd153448: dataIn1 = 32'd4771
; 
32'd153449: dataIn1 = 32'd5089
; 
32'd153450: dataIn1 = 32'd5091
; 
32'd153451: dataIn1 = 32'd8720
; 
32'd153452: dataIn1 = 32'd8721
; 
32'd153453: dataIn1 = 32'd8723
; 
32'd153454: dataIn1 = 32'd8725
; 
32'd153455: dataIn1 = 32'd5081
; 
32'd153456: dataIn1 = 32'd5090
; 
32'd153457: dataIn1 = 32'd5092
; 
32'd153458: dataIn1 = 32'd8733
; 
32'd153459: dataIn1 = 32'd8734
; 
32'd153460: dataIn1 = 32'd8735
; 
32'd153461: dataIn1 = 32'd8736
; 
32'd153462: dataIn1 = 32'd2688
; 
32'd153463: dataIn1 = 32'd2689
; 
32'd153464: dataIn1 = 32'd5093
; 
32'd153465: dataIn1 = 32'd5094
; 
32'd153466: dataIn1 = 32'd5095
; 
32'd153467: dataIn1 = 32'd5096
; 
32'd153468: dataIn1 = 32'd5097
; 
32'd153469: dataIn1 = 32'd2687
; 
32'd153470: dataIn1 = 32'd2689
; 
32'd153471: dataIn1 = 32'd5093
; 
32'd153472: dataIn1 = 32'd5094
; 
32'd153473: dataIn1 = 32'd5095
; 
32'd153474: dataIn1 = 32'd5098
; 
32'd153475: dataIn1 = 32'd5099
; 
32'd153476: dataIn1 = 32'd2687
; 
32'd153477: dataIn1 = 32'd2688
; 
32'd153478: dataIn1 = 32'd5093
; 
32'd153479: dataIn1 = 32'd5094
; 
32'd153480: dataIn1 = 32'd5095
; 
32'd153481: dataIn1 = 32'd5100
; 
32'd153482: dataIn1 = 32'd5101
; 
32'd153483: dataIn1 = 32'd1100
; 
32'd153484: dataIn1 = 32'd2689
; 
32'd153485: dataIn1 = 32'd4786
; 
32'd153486: dataIn1 = 32'd5093
; 
32'd153487: dataIn1 = 32'd5096
; 
32'd153488: dataIn1 = 32'd5097
; 
32'd153489: dataIn1 = 32'd5107
; 
32'd153490: dataIn1 = 32'd1100
; 
32'd153491: dataIn1 = 32'd2688
; 
32'd153492: dataIn1 = 32'd3569
; 
32'd153493: dataIn1 = 32'd5093
; 
32'd153494: dataIn1 = 32'd5096
; 
32'd153495: dataIn1 = 32'd5097
; 
32'd153496: dataIn1 = 32'd1118
; 
32'd153497: dataIn1 = 32'd2689
; 
32'd153498: dataIn1 = 32'd5094
; 
32'd153499: dataIn1 = 32'd5098
; 
32'd153500: dataIn1 = 32'd5099
; 
32'd153501: dataIn1 = 32'd5108
; 
32'd153502: dataIn1 = 32'd5110
; 
32'd153503: dataIn1 = 32'd8856
; 
32'd153504: dataIn1 = 32'd1118
; 
32'd153505: dataIn1 = 32'd2687
; 
32'd153506: dataIn1 = 32'd5094
; 
32'd153507: dataIn1 = 32'd5098
; 
32'd153508: dataIn1 = 32'd5099
; 
32'd153509: dataIn1 = 32'd5103
; 
32'd153510: dataIn1 = 32'd5106
; 
32'd153511: dataIn1 = 32'd8834
; 
32'd153512: dataIn1 = 32'd1099
; 
32'd153513: dataIn1 = 32'd2688
; 
32'd153514: dataIn1 = 32'd3567
; 
32'd153515: dataIn1 = 32'd5095
; 
32'd153516: dataIn1 = 32'd5100
; 
32'd153517: dataIn1 = 32'd5101
; 
32'd153518: dataIn1 = 32'd1099
; 
32'd153519: dataIn1 = 32'd2687
; 
32'd153520: dataIn1 = 32'd4781
; 
32'd153521: dataIn1 = 32'd5095
; 
32'd153522: dataIn1 = 32'd5100
; 
32'd153523: dataIn1 = 32'd5101
; 
32'd153524: dataIn1 = 32'd5104
; 
32'd153525: dataIn1 = 32'd2602
; 
32'd153526: dataIn1 = 32'd2690
; 
32'd153527: dataIn1 = 32'd4778
; 
32'd153528: dataIn1 = 32'd5102
; 
32'd153529: dataIn1 = 32'd5103
; 
32'd153530: dataIn1 = 32'd5104
; 
32'd153531: dataIn1 = 32'd5105
; 
32'd153532: dataIn1 = 32'd8840
; 
32'd153533: dataIn1 = 32'd2687
; 
32'd153534: dataIn1 = 32'd2690
; 
32'd153535: dataIn1 = 32'd5099
; 
32'd153536: dataIn1 = 32'd5102
; 
32'd153537: dataIn1 = 32'd5103
; 
32'd153538: dataIn1 = 32'd5104
; 
32'd153539: dataIn1 = 32'd5106
; 
32'd153540: dataIn1 = 32'd8835
; 
32'd153541: dataIn1 = 32'd2602
; 
32'd153542: dataIn1 = 32'd2687
; 
32'd153543: dataIn1 = 32'd4781
; 
32'd153544: dataIn1 = 32'd5101
; 
32'd153545: dataIn1 = 32'd5102
; 
32'd153546: dataIn1 = 32'd5103
; 
32'd153547: dataIn1 = 32'd5104
; 
32'd153548: dataIn1 = 32'd4778
; 
32'd153549: dataIn1 = 32'd5102
; 
32'd153550: dataIn1 = 32'd5105
; 
32'd153551: dataIn1 = 32'd8837
; 
32'd153552: dataIn1 = 32'd8838
; 
32'd153553: dataIn1 = 32'd8839
; 
32'd153554: dataIn1 = 32'd8840
; 
32'd153555: dataIn1 = 32'd5099
; 
32'd153556: dataIn1 = 32'd5103
; 
32'd153557: dataIn1 = 32'd5106
; 
32'd153558: dataIn1 = 32'd8831
; 
32'd153559: dataIn1 = 32'd8833
; 
32'd153560: dataIn1 = 32'd8834
; 
32'd153561: dataIn1 = 32'd8835
; 
32'd153562: dataIn1 = 32'd2606
; 
32'd153563: dataIn1 = 32'd2689
; 
32'd153564: dataIn1 = 32'd4786
; 
32'd153565: dataIn1 = 32'd5096
; 
32'd153566: dataIn1 = 32'd5107
; 
32'd153567: dataIn1 = 32'd5108
; 
32'd153568: dataIn1 = 32'd5109
; 
32'd153569: dataIn1 = 32'd2689
; 
32'd153570: dataIn1 = 32'd2691
; 
32'd153571: dataIn1 = 32'd5098
; 
32'd153572: dataIn1 = 32'd5107
; 
32'd153573: dataIn1 = 32'd5108
; 
32'd153574: dataIn1 = 32'd5109
; 
32'd153575: dataIn1 = 32'd5110
; 
32'd153576: dataIn1 = 32'd8857
; 
32'd153577: dataIn1 = 32'd2606
; 
32'd153578: dataIn1 = 32'd2691
; 
32'd153579: dataIn1 = 32'd4788
; 
32'd153580: dataIn1 = 32'd5107
; 
32'd153581: dataIn1 = 32'd5108
; 
32'd153582: dataIn1 = 32'd5109
; 
32'd153583: dataIn1 = 32'd5111
; 
32'd153584: dataIn1 = 32'd8867
; 
32'd153585: dataIn1 = 32'd5098
; 
32'd153586: dataIn1 = 32'd5108
; 
32'd153587: dataIn1 = 32'd5110
; 
32'd153588: dataIn1 = 32'd8853
; 
32'd153589: dataIn1 = 32'd8854
; 
32'd153590: dataIn1 = 32'd8856
; 
32'd153591: dataIn1 = 32'd8857
; 
32'd153592: dataIn1 = 32'd4788
; 
32'd153593: dataIn1 = 32'd5109
; 
32'd153594: dataIn1 = 32'd5111
; 
32'd153595: dataIn1 = 32'd8864
; 
32'd153596: dataIn1 = 32'd8865
; 
32'd153597: dataIn1 = 32'd8867
; 
32'd153598: dataIn1 = 32'd8869
; 
32'd153599: dataIn1 = 32'd5112
; 
32'd153600: dataIn1 = 32'd6073
; 
32'd153601: dataIn1 = 32'd6077
; 
32'd153602: dataIn1 = 32'd7058
; 
32'd153603: dataIn1 = 32'd7059
; 
32'd153604: dataIn1 = 32'd7074
; 
32'd153605: dataIn1 = 32'd7081
; 
32'd153606: dataIn1 = 32'd5113
; 
32'd153607: dataIn1 = 32'd7060
; 
32'd153608: dataIn1 = 32'd7061
; 
32'd153609: dataIn1 = 32'd7069
; 
32'd153610: dataIn1 = 32'd7075
; 
32'd153611: dataIn1 = 32'd7090
; 
32'd153612: dataIn1 = 32'd7091
; 
32'd153613: dataIn1 = 32'd5114
; 
32'd153614: dataIn1 = 32'd6072
; 
32'd153615: dataIn1 = 32'd6091
; 
32'd153616: dataIn1 = 32'd7062
; 
32'd153617: dataIn1 = 32'd7063
; 
32'd153618: dataIn1 = 32'd7070
; 
32'd153619: dataIn1 = 32'd7110
; 
32'd153620: dataIn1 = 32'd5115
; 
32'd153621: dataIn1 = 32'd6076
; 
32'd153622: dataIn1 = 32'd6080
; 
32'd153623: dataIn1 = 32'd7082
; 
32'd153624: dataIn1 = 32'd7083
; 
32'd153625: dataIn1 = 32'd7191
; 
32'd153626: dataIn1 = 32'd7192
; 
32'd153627: dataIn1 = 32'd5116
; 
32'd153628: dataIn1 = 32'd6076
; 
32'd153629: dataIn1 = 32'd6077
; 
32'd153630: dataIn1 = 32'd6079
; 
32'd153631: dataIn1 = 32'd6081
; 
32'd153632: dataIn1 = 32'd6704
; 
32'd153633: dataIn1 = 32'd6705
; 
32'd153634: dataIn1 = 32'd5117
; 
32'd153635: dataIn1 = 32'd7088
; 
32'd153636: dataIn1 = 32'd7089
; 
32'd153637: dataIn1 = 32'd7102
; 
32'd153638: dataIn1 = 32'd7206
; 
32'd153639: dataIn1 = 32'd9790
; 
32'd153640: dataIn1 = 32'd9791
; 
32'd153641: dataIn1 = 32'd5118
; 
32'd153642: dataIn1 = 32'd7092
; 
32'd153643: dataIn1 = 32'd7093
; 
32'd153644: dataIn1 = 32'd7098
; 
32'd153645: dataIn1 = 32'd7145
; 
32'd153646: dataIn1 = 32'd9794
; 
32'd153647: dataIn1 = 32'd9795
; 
32'd153648: dataIn1 = 32'd5119
; 
32'd153649: dataIn1 = 32'd6091
; 
32'd153650: dataIn1 = 32'd6092
; 
32'd153651: dataIn1 = 32'd6094
; 
32'd153652: dataIn1 = 32'd6096
; 
32'd153653: dataIn1 = 32'd6706
; 
32'd153654: dataIn1 = 32'd6707
; 
32'd153655: dataIn1 = 32'd5120
; 
32'd153656: dataIn1 = 32'd6092
; 
32'd153657: dataIn1 = 32'd6095
; 
32'd153658: dataIn1 = 32'd7108
; 
32'd153659: dataIn1 = 32'd7109
; 
32'd153660: dataIn1 = 32'd7151
; 
32'd153661: dataIn1 = 32'd7152
; 
32'd153662: dataIn1 = 32'd5121
; 
32'd153663: dataIn1 = 32'd7114
; 
32'd153664: dataIn1 = 32'd7115
; 
32'd153665: dataIn1 = 32'd7130
; 
32'd153666: dataIn1 = 32'd7137
; 
32'd153667: dataIn1 = 32'd9802
; 
32'd153668: dataIn1 = 32'd9803
; 
32'd153669: dataIn1 = 32'd5122
; 
32'd153670: dataIn1 = 32'd7116
; 
32'd153671: dataIn1 = 32'd7117
; 
32'd153672: dataIn1 = 32'd7125
; 
32'd153673: dataIn1 = 32'd7144
; 
32'd153674: dataIn1 = 32'd9798
; 
32'd153675: dataIn1 = 32'd9799
; 
32'd153676: dataIn1 = 32'd5123
; 
32'd153677: dataIn1 = 32'd7118
; 
32'd153678: dataIn1 = 32'd7119
; 
32'd153679: dataIn1 = 32'd7126
; 
32'd153680: dataIn1 = 32'd7133
; 
32'd153681: dataIn1 = 32'd7153
; 
32'd153682: dataIn1 = 32'd7154
; 
32'd153683: dataIn1 = 32'd5124
; 
32'd153684: dataIn1 = 32'd7139
; 
32'd153685: dataIn1 = 32'd7140
; 
32'd153686: dataIn1 = 32'd9368
; 
32'd153687: dataIn1 = 32'd9369
; 
32'd153688: dataIn1 = 32'd9806
; 
32'd153689: dataIn1 = 32'd9807
; 
32'd153690: dataIn1 = 32'd5125
; 
32'd153691: dataIn1 = 32'd6118
; 
32'd153692: dataIn1 = 32'd6817
; 
32'd153693: dataIn1 = 32'd7149
; 
32'd153694: dataIn1 = 32'd7150
; 
32'd153695: dataIn1 = 32'd7161
; 
32'd153696: dataIn1 = 32'd9446
; 
32'd153697: dataIn1 = 32'd5126
; 
32'd153698: dataIn1 = 32'd7166
; 
32'd153699: dataIn1 = 32'd7167
; 
32'd153700: dataIn1 = 32'd7175
; 
32'd153701: dataIn1 = 32'd7182
; 
32'd153702: dataIn1 = 32'd7189
; 
32'd153703: dataIn1 = 32'd7190
; 
32'd153704: dataIn1 = 32'd5127
; 
32'd153705: dataIn1 = 32'd7168
; 
32'd153706: dataIn1 = 32'd7169
; 
32'd153707: dataIn1 = 32'd7183
; 
32'd153708: dataIn1 = 32'd7207
; 
32'd153709: dataIn1 = 32'd9786
; 
32'd153710: dataIn1 = 32'd9787
; 
32'd153711: dataIn1 = 32'd5128
; 
32'd153712: dataIn1 = 32'd7170
; 
32'd153713: dataIn1 = 32'd7171
; 
32'd153714: dataIn1 = 32'd7178
; 
32'd153715: dataIn1 = 32'd7213
; 
32'd153716: dataIn1 = 32'd7214
; 
32'd153717: dataIn1 = 32'd9759
; 
32'd153718: dataIn1 = 32'd5129
; 
32'd153719: dataIn1 = 32'd6131
; 
32'd153720: dataIn1 = 32'd6592
; 
32'd153721: dataIn1 = 32'd7193
; 
32'd153722: dataIn1 = 32'd7194
; 
32'd153723: dataIn1 = 32'd7199
; 
32'd153724: dataIn1 = 32'd8919
; 
32'd153725: dataIn1 = 32'd5130
; 
32'd153726: dataIn1 = 32'd7211
; 
32'd153727: dataIn1 = 32'd7212
; 
32'd153728: dataIn1 = 32'd7218
; 
32'd153729: dataIn1 = 32'd7221
; 
32'd153730: dataIn1 = 32'd8900
; 
32'd153731: dataIn1 = 32'd8901
; 
32'd153732: dataIn1 = 32'd2698
; 
32'd153733: dataIn1 = 32'd5131
; 
32'd153734: dataIn1 = 32'd5133
; 
32'd153735: dataIn1 = 32'd5135
; 
32'd153736: dataIn1 = 32'd6142
; 
32'd153737: dataIn1 = 32'd6143
; 
32'd153738: dataIn1 = 32'd6145
; 
32'd153739: dataIn1 = 32'd5132
; 
32'd153740: dataIn1 = 32'd5133
; 
32'd153741: dataIn1 = 32'd6143
; 
32'd153742: dataIn1 = 32'd6150
; 
32'd153743: dataIn1 = 32'd7227
; 
32'd153744: dataIn1 = 32'd7228
; 
32'd153745: dataIn1 = 32'd7244
; 
32'd153746: dataIn1 = 32'd2697
; 
32'd153747: dataIn1 = 32'd2698
; 
32'd153748: dataIn1 = 32'd5131
; 
32'd153749: dataIn1 = 32'd5132
; 
32'd153750: dataIn1 = 32'd5133
; 
32'd153751: dataIn1 = 32'd5138
; 
32'd153752: dataIn1 = 32'd5139
; 
32'd153753: dataIn1 = 32'd6143
; 
32'd153754: dataIn1 = 32'd6150
; 
32'd153755: dataIn1 = 32'd1121
; 
32'd153756: dataIn1 = 32'd5134
; 
32'd153757: dataIn1 = 32'd5135
; 
32'd153758: dataIn1 = 32'd6144
; 
32'd153759: dataIn1 = 32'd6145
; 
32'd153760: dataIn1 = 32'd6177
; 
32'd153761: dataIn1 = 32'd6179
; 
32'd153762: dataIn1 = 32'd1121
; 
32'd153763: dataIn1 = 32'd2698
; 
32'd153764: dataIn1 = 32'd2702
; 
32'd153765: dataIn1 = 32'd5131
; 
32'd153766: dataIn1 = 32'd5134
; 
32'd153767: dataIn1 = 32'd5135
; 
32'd153768: dataIn1 = 32'd6145
; 
32'd153769: dataIn1 = 32'd5136
; 
32'd153770: dataIn1 = 32'd7225
; 
32'd153771: dataIn1 = 32'd7226
; 
32'd153772: dataIn1 = 32'd7236
; 
32'd153773: dataIn1 = 32'd7243
; 
32'd153774: dataIn1 = 32'd7320
; 
32'd153775: dataIn1 = 32'd7321
; 
32'd153776: dataIn1 = 32'd5137
; 
32'd153777: dataIn1 = 32'd7229
; 
32'd153778: dataIn1 = 32'd7230
; 
32'd153779: dataIn1 = 32'd7231
; 
32'd153780: dataIn1 = 32'd7239
; 
32'd153781: dataIn1 = 32'd7270
; 
32'd153782: dataIn1 = 32'd7271
; 
32'd153783: dataIn1 = 32'd1122
; 
32'd153784: dataIn1 = 32'd2698
; 
32'd153785: dataIn1 = 32'd2701
; 
32'd153786: dataIn1 = 32'd5133
; 
32'd153787: dataIn1 = 32'd5138
; 
32'd153788: dataIn1 = 32'd5139
; 
32'd153789: dataIn1 = 32'd1122
; 
32'd153790: dataIn1 = 32'd2697
; 
32'd153791: dataIn1 = 32'd5133
; 
32'd153792: dataIn1 = 32'd5138
; 
32'd153793: dataIn1 = 32'd5139
; 
32'd153794: dataIn1 = 32'd5142
; 
32'd153795: dataIn1 = 32'd5144
; 
32'd153796: dataIn1 = 32'd6157
; 
32'd153797: dataIn1 = 32'd5140
; 
32'd153798: dataIn1 = 32'd7250
; 
32'd153799: dataIn1 = 32'd7251
; 
32'd153800: dataIn1 = 32'd7262
; 
32'd153801: dataIn1 = 32'd9760
; 
32'd153802: dataIn1 = 32'd10122
; 
32'd153803: dataIn1 = 32'd10123
; 
32'd153804: dataIn1 = 32'd5141
; 
32'd153805: dataIn1 = 32'd7252
; 
32'd153806: dataIn1 = 32'd7253
; 
32'd153807: dataIn1 = 32'd7268
; 
32'd153808: dataIn1 = 32'd7269
; 
32'd153809: dataIn1 = 32'd7275
; 
32'd153810: dataIn1 = 32'd9761
; 
32'd153811: dataIn1 = 32'd5139
; 
32'd153812: dataIn1 = 32'd5142
; 
32'd153813: dataIn1 = 32'd5144
; 
32'd153814: dataIn1 = 32'd6154
; 
32'd153815: dataIn1 = 32'd6155
; 
32'd153816: dataIn1 = 32'd6157
; 
32'd153817: dataIn1 = 32'd9668
; 
32'd153818: dataIn1 = 32'd9734
; 
32'd153819: dataIn1 = 32'd5143
; 
32'd153820: dataIn1 = 32'd9745
; 
32'd153821: dataIn1 = 32'd9746
; 
32'd153822: dataIn1 = 32'd9767
; 
32'd153823: dataIn1 = 32'd9778
; 
32'd153824: dataIn1 = 32'd10124
; 
32'd153825: dataIn1 = 32'd10125
; 
32'd153826: dataIn1 = 32'd1122
; 
32'd153827: dataIn1 = 32'd2700
; 
32'd153828: dataIn1 = 32'd5139
; 
32'd153829: dataIn1 = 32'd5142
; 
32'd153830: dataIn1 = 32'd5144
; 
32'd153831: dataIn1 = 32'd5270
; 
32'd153832: dataIn1 = 32'd5272
; 
32'd153833: dataIn1 = 32'd9668
; 
32'd153834: dataIn1 = 32'd5145
; 
32'd153835: dataIn1 = 32'd6179
; 
32'd153836: dataIn1 = 32'd7285
; 
32'd153837: dataIn1 = 32'd7286
; 
32'd153838: dataIn1 = 32'd7301
; 
32'd153839: dataIn1 = 32'd7308
; 
32'd153840: dataIn1 = 32'd7315
; 
32'd153841: dataIn1 = 32'd5146
; 
32'd153842: dataIn1 = 32'd7287
; 
32'd153843: dataIn1 = 32'd7288
; 
32'd153844: dataIn1 = 32'd7296
; 
32'd153845: dataIn1 = 32'd7309
; 
32'd153846: dataIn1 = 32'd7322
; 
32'd153847: dataIn1 = 32'd7323
; 
32'd153848: dataIn1 = 32'd5147
; 
32'd153849: dataIn1 = 32'd7289
; 
32'd153850: dataIn1 = 32'd7290
; 
32'd153851: dataIn1 = 32'd7297
; 
32'd153852: dataIn1 = 32'd7304
; 
32'd153853: dataIn1 = 32'd7342
; 
32'd153854: dataIn1 = 32'd7343
; 
32'd153855: dataIn1 = 32'd1121
; 
32'd153856: dataIn1 = 32'd5148
; 
32'd153857: dataIn1 = 32'd5278
; 
32'd153858: dataIn1 = 32'd6177
; 
32'd153859: dataIn1 = 32'd6178
; 
32'd153860: dataIn1 = 32'd6180
; 
32'd153861: dataIn1 = 32'd6610
; 
32'd153862: dataIn1 = 32'd7314
; 
32'd153863: dataIn1 = 32'd5149
; 
32'd153864: dataIn1 = 32'd7338
; 
32'd153865: dataIn1 = 32'd7339
; 
32'd153866: dataIn1 = 32'd7350
; 
32'd153867: dataIn1 = 32'd7355
; 
32'd153868: dataIn1 = 32'd8957
; 
32'd153869: dataIn1 = 32'd8958
; 
32'd153870: dataIn1 = 32'd5150
; 
32'd153871: dataIn1 = 32'd6745
; 
32'd153872: dataIn1 = 32'd6747
; 
32'd153873: dataIn1 = 32'd7359
; 
32'd153874: dataIn1 = 32'd7360
; 
32'd153875: dataIn1 = 32'd7375
; 
32'd153876: dataIn1 = 32'd7382
; 
32'd153877: dataIn1 = 32'd5151
; 
32'd153878: dataIn1 = 32'd7361
; 
32'd153879: dataIn1 = 32'd7362
; 
32'd153880: dataIn1 = 32'd7370
; 
32'd153881: dataIn1 = 32'd7376
; 
32'd153882: dataIn1 = 32'd7391
; 
32'd153883: dataIn1 = 32'd7392
; 
32'd153884: dataIn1 = 32'd5152
; 
32'd153885: dataIn1 = 32'd6744
; 
32'd153886: dataIn1 = 32'd6748
; 
32'd153887: dataIn1 = 32'd7363
; 
32'd153888: dataIn1 = 32'd7364
; 
32'd153889: dataIn1 = 32'd7371
; 
32'd153890: dataIn1 = 32'd7418
; 
32'd153891: dataIn1 = 32'd5153
; 
32'd153892: dataIn1 = 32'd6746
; 
32'd153893: dataIn1 = 32'd6753
; 
32'd153894: dataIn1 = 32'd7383
; 
32'd153895: dataIn1 = 32'd7384
; 
32'd153896: dataIn1 = 32'd7547
; 
32'd153897: dataIn1 = 32'd7548
; 
32'd153898: dataIn1 = 32'd5154
; 
32'd153899: dataIn1 = 32'd6746
; 
32'd153900: dataIn1 = 32'd6747
; 
32'd153901: dataIn1 = 32'd9235
; 
32'd153902: dataIn1 = 32'd9237
; 
32'd153903: dataIn1 = 32'd9287
; 
32'd153904: dataIn1 = 32'd9288
; 
32'd153905: dataIn1 = 32'd5155
; 
32'd153906: dataIn1 = 32'd7389
; 
32'd153907: dataIn1 = 32'd7390
; 
32'd153908: dataIn1 = 32'd7403
; 
32'd153909: dataIn1 = 32'd7410
; 
32'd153910: dataIn1 = 32'd7562
; 
32'd153911: dataIn1 = 32'd7563
; 
32'd153912: dataIn1 = 32'd5156
; 
32'd153913: dataIn1 = 32'd7393
; 
32'd153914: dataIn1 = 32'd7394
; 
32'd153915: dataIn1 = 32'd7399
; 
32'd153916: dataIn1 = 32'd7406
; 
32'd153917: dataIn1 = 32'd7480
; 
32'd153918: dataIn1 = 32'd7481
; 
32'd153919: dataIn1 = 32'd5157
; 
32'd153920: dataIn1 = 32'd6748
; 
32'd153921: dataIn1 = 32'd6749
; 
32'd153922: dataIn1 = 32'd9236
; 
32'd153923: dataIn1 = 32'd9238
; 
32'd153924: dataIn1 = 32'd9289
; 
32'd153925: dataIn1 = 32'd9290
; 
32'd153926: dataIn1 = 32'd5158
; 
32'd153927: dataIn1 = 32'd6749
; 
32'd153928: dataIn1 = 32'd6750
; 
32'd153929: dataIn1 = 32'd7416
; 
32'd153930: dataIn1 = 32'd7417
; 
32'd153931: dataIn1 = 32'd7500
; 
32'd153932: dataIn1 = 32'd7501
; 
32'd153933: dataIn1 = 32'd5159
; 
32'd153934: dataIn1 = 32'd7422
; 
32'd153935: dataIn1 = 32'd7423
; 
32'd153936: dataIn1 = 32'd7438
; 
32'd153937: dataIn1 = 32'd7445
; 
32'd153938: dataIn1 = 32'd7452
; 
32'd153939: dataIn1 = 32'd7453
; 
32'd153940: dataIn1 = 32'd5160
; 
32'd153941: dataIn1 = 32'd7424
; 
32'd153942: dataIn1 = 32'd7425
; 
32'd153943: dataIn1 = 32'd7433
; 
32'd153944: dataIn1 = 32'd7446
; 
32'd153945: dataIn1 = 32'd7478
; 
32'd153946: dataIn1 = 32'd7479
; 
32'd153947: dataIn1 = 32'd5161
; 
32'd153948: dataIn1 = 32'd7426
; 
32'd153949: dataIn1 = 32'd7427
; 
32'd153950: dataIn1 = 32'd7434
; 
32'd153951: dataIn1 = 32'd7441
; 
32'd153952: dataIn1 = 32'd7502
; 
32'd153953: dataIn1 = 32'd7503
; 
32'd153954: dataIn1 = 32'd5162
; 
32'd153955: dataIn1 = 32'd7456
; 
32'd153956: dataIn1 = 32'd7457
; 
32'd153957: dataIn1 = 32'd7462
; 
32'd153958: dataIn1 = 32'd7467
; 
32'd153959: dataIn1 = 32'd8955
; 
32'd153960: dataIn1 = 32'd8956
; 
32'd153961: dataIn1 = 32'd5163
; 
32'd153962: dataIn1 = 32'd6751
; 
32'd153963: dataIn1 = 32'd7498
; 
32'd153964: dataIn1 = 32'd7499
; 
32'd153965: dataIn1 = 32'd7510
; 
32'd153966: dataIn1 = 32'd8973
; 
32'd153967: dataIn1 = 32'd9280
; 
32'd153968: dataIn1 = 32'd5164
; 
32'd153969: dataIn1 = 32'd7515
; 
32'd153970: dataIn1 = 32'd7516
; 
32'd153971: dataIn1 = 32'd7531
; 
32'd153972: dataIn1 = 32'd7538
; 
32'd153973: dataIn1 = 32'd7545
; 
32'd153974: dataIn1 = 32'd7546
; 
32'd153975: dataIn1 = 32'd5165
; 
32'd153976: dataIn1 = 32'd7517
; 
32'd153977: dataIn1 = 32'd7518
; 
32'd153978: dataIn1 = 32'd7526
; 
32'd153979: dataIn1 = 32'd7539
; 
32'd153980: dataIn1 = 32'd7564
; 
32'd153981: dataIn1 = 32'd7565
; 
32'd153982: dataIn1 = 32'd5166
; 
32'd153983: dataIn1 = 32'd7519
; 
32'd153984: dataIn1 = 32'd7520
; 
32'd153985: dataIn1 = 32'd7527
; 
32'd153986: dataIn1 = 32'd7534
; 
32'd153987: dataIn1 = 32'd7588
; 
32'd153988: dataIn1 = 32'd7589
; 
32'd153989: dataIn1 = 32'd5167
; 
32'd153990: dataIn1 = 32'd6752
; 
32'd153991: dataIn1 = 32'd6791
; 
32'd153992: dataIn1 = 32'd7549
; 
32'd153993: dataIn1 = 32'd7550
; 
32'd153994: dataIn1 = 32'd7555
; 
32'd153995: dataIn1 = 32'd9025
; 
32'd153996: dataIn1 = 32'd5168
; 
32'd153997: dataIn1 = 32'd7584
; 
32'd153998: dataIn1 = 32'd7585
; 
32'd153999: dataIn1 = 32'd7598
; 
32'd154000: dataIn1 = 32'd7603
; 
32'd154001: dataIn1 = 32'd9006
; 
32'd154002: dataIn1 = 32'd9007
; 
32'd154003: dataIn1 = 32'd5169
; 
32'd154004: dataIn1 = 32'd6755
; 
32'd154005: dataIn1 = 32'd6757
; 
32'd154006: dataIn1 = 32'd7610
; 
32'd154007: dataIn1 = 32'd7611
; 
32'd154008: dataIn1 = 32'd7626
; 
32'd154009: dataIn1 = 32'd7633
; 
32'd154010: dataIn1 = 32'd5170
; 
32'd154011: dataIn1 = 32'd7612
; 
32'd154012: dataIn1 = 32'd7613
; 
32'd154013: dataIn1 = 32'd7621
; 
32'd154014: dataIn1 = 32'd7627
; 
32'd154015: dataIn1 = 32'd7642
; 
32'd154016: dataIn1 = 32'd7643
; 
32'd154017: dataIn1 = 32'd5171
; 
32'd154018: dataIn1 = 32'd6754
; 
32'd154019: dataIn1 = 32'd6758
; 
32'd154020: dataIn1 = 32'd7614
; 
32'd154021: dataIn1 = 32'd7615
; 
32'd154022: dataIn1 = 32'd7622
; 
32'd154023: dataIn1 = 32'd7669
; 
32'd154024: dataIn1 = 32'd5172
; 
32'd154025: dataIn1 = 32'd6756
; 
32'd154026: dataIn1 = 32'd6763
; 
32'd154027: dataIn1 = 32'd7634
; 
32'd154028: dataIn1 = 32'd7635
; 
32'd154029: dataIn1 = 32'd7800
; 
32'd154030: dataIn1 = 32'd7801
; 
32'd154031: dataIn1 = 32'd5173
; 
32'd154032: dataIn1 = 32'd6756
; 
32'd154033: dataIn1 = 32'd6757
; 
32'd154034: dataIn1 = 32'd9240
; 
32'd154035: dataIn1 = 32'd9242
; 
32'd154036: dataIn1 = 32'd9293
; 
32'd154037: dataIn1 = 32'd9294
; 
32'd154038: dataIn1 = 32'd5174
; 
32'd154039: dataIn1 = 32'd7640
; 
32'd154040: dataIn1 = 32'd7641
; 
32'd154041: dataIn1 = 32'd7654
; 
32'd154042: dataIn1 = 32'd7661
; 
32'd154043: dataIn1 = 32'd7815
; 
32'd154044: dataIn1 = 32'd7816
; 
32'd154045: dataIn1 = 32'd5175
; 
32'd154046: dataIn1 = 32'd7644
; 
32'd154047: dataIn1 = 32'd7645
; 
32'd154048: dataIn1 = 32'd7650
; 
32'd154049: dataIn1 = 32'd7657
; 
32'd154050: dataIn1 = 32'd7733
; 
32'd154051: dataIn1 = 32'd7734
; 
32'd154052: dataIn1 = 32'd5176
; 
32'd154053: dataIn1 = 32'd6758
; 
32'd154054: dataIn1 = 32'd6759
; 
32'd154055: dataIn1 = 32'd9241
; 
32'd154056: dataIn1 = 32'd9243
; 
32'd154057: dataIn1 = 32'd9295
; 
32'd154058: dataIn1 = 32'd9296
; 
32'd154059: dataIn1 = 32'd5177
; 
32'd154060: dataIn1 = 32'd6759
; 
32'd154061: dataIn1 = 32'd6760
; 
32'd154062: dataIn1 = 32'd7667
; 
32'd154063: dataIn1 = 32'd7668
; 
32'd154064: dataIn1 = 32'd7753
; 
32'd154065: dataIn1 = 32'd7754
; 
32'd154066: dataIn1 = 32'd5178
; 
32'd154067: dataIn1 = 32'd7673
; 
32'd154068: dataIn1 = 32'd7674
; 
32'd154069: dataIn1 = 32'd7689
; 
32'd154070: dataIn1 = 32'd7696
; 
32'd154071: dataIn1 = 32'd7703
; 
32'd154072: dataIn1 = 32'd7704
; 
32'd154073: dataIn1 = 32'd5179
; 
32'd154074: dataIn1 = 32'd7675
; 
32'd154075: dataIn1 = 32'd7676
; 
32'd154076: dataIn1 = 32'd7684
; 
32'd154077: dataIn1 = 32'd7697
; 
32'd154078: dataIn1 = 32'd7731
; 
32'd154079: dataIn1 = 32'd7732
; 
32'd154080: dataIn1 = 32'd5180
; 
32'd154081: dataIn1 = 32'd7677
; 
32'd154082: dataIn1 = 32'd7678
; 
32'd154083: dataIn1 = 32'd7685
; 
32'd154084: dataIn1 = 32'd7692
; 
32'd154085: dataIn1 = 32'd7755
; 
32'd154086: dataIn1 = 32'd7756
; 
32'd154087: dataIn1 = 32'd5181
; 
32'd154088: dataIn1 = 32'd7707
; 
32'd154089: dataIn1 = 32'd7708
; 
32'd154090: dataIn1 = 32'd7715
; 
32'd154091: dataIn1 = 32'd7720
; 
32'd154092: dataIn1 = 32'd9004
; 
32'd154093: dataIn1 = 32'd9005
; 
32'd154094: dataIn1 = 32'd5182
; 
32'd154095: dataIn1 = 32'd6761
; 
32'd154096: dataIn1 = 32'd6789
; 
32'd154097: dataIn1 = 32'd7751
; 
32'd154098: dataIn1 = 32'd7752
; 
32'd154099: dataIn1 = 32'd7763
; 
32'd154100: dataIn1 = 32'd9020
; 
32'd154101: dataIn1 = 32'd5183
; 
32'd154102: dataIn1 = 32'd7768
; 
32'd154103: dataIn1 = 32'd7769
; 
32'd154104: dataIn1 = 32'd7784
; 
32'd154105: dataIn1 = 32'd7791
; 
32'd154106: dataIn1 = 32'd7798
; 
32'd154107: dataIn1 = 32'd7799
; 
32'd154108: dataIn1 = 32'd5184
; 
32'd154109: dataIn1 = 32'd7770
; 
32'd154110: dataIn1 = 32'd7771
; 
32'd154111: dataIn1 = 32'd7779
; 
32'd154112: dataIn1 = 32'd7792
; 
32'd154113: dataIn1 = 32'd7817
; 
32'd154114: dataIn1 = 32'd7818
; 
32'd154115: dataIn1 = 32'd5185
; 
32'd154116: dataIn1 = 32'd7772
; 
32'd154117: dataIn1 = 32'd7773
; 
32'd154118: dataIn1 = 32'd7780
; 
32'd154119: dataIn1 = 32'd7787
; 
32'd154120: dataIn1 = 32'd7841
; 
32'd154121: dataIn1 = 32'd7842
; 
32'd154122: dataIn1 = 32'd5186
; 
32'd154123: dataIn1 = 32'd6762
; 
32'd154124: dataIn1 = 32'd6793
; 
32'd154125: dataIn1 = 32'd7802
; 
32'd154126: dataIn1 = 32'd7803
; 
32'd154127: dataIn1 = 32'd7808
; 
32'd154128: dataIn1 = 32'd9077
; 
32'd154129: dataIn1 = 32'd5187
; 
32'd154130: dataIn1 = 32'd7837
; 
32'd154131: dataIn1 = 32'd7838
; 
32'd154132: dataIn1 = 32'd7851
; 
32'd154133: dataIn1 = 32'd7856
; 
32'd154134: dataIn1 = 32'd9058
; 
32'd154135: dataIn1 = 32'd9059
; 
32'd154136: dataIn1 = 32'd5188
; 
32'd154137: dataIn1 = 32'd6315
; 
32'd154138: dataIn1 = 32'd6322
; 
32'd154139: dataIn1 = 32'd7863
; 
32'd154140: dataIn1 = 32'd7864
; 
32'd154141: dataIn1 = 32'd7879
; 
32'd154142: dataIn1 = 32'd7886
; 
32'd154143: dataIn1 = 32'd5189
; 
32'd154144: dataIn1 = 32'd7865
; 
32'd154145: dataIn1 = 32'd7866
; 
32'd154146: dataIn1 = 32'd7874
; 
32'd154147: dataIn1 = 32'd7880
; 
32'd154148: dataIn1 = 32'd7895
; 
32'd154149: dataIn1 = 32'd7896
; 
32'd154150: dataIn1 = 32'd5190
; 
32'd154151: dataIn1 = 32'd6314
; 
32'd154152: dataIn1 = 32'd6334
; 
32'd154153: dataIn1 = 32'd7867
; 
32'd154154: dataIn1 = 32'd7868
; 
32'd154155: dataIn1 = 32'd7875
; 
32'd154156: dataIn1 = 32'd7922
; 
32'd154157: dataIn1 = 32'd5191
; 
32'd154158: dataIn1 = 32'd6318
; 
32'd154159: dataIn1 = 32'd6320
; 
32'd154160: dataIn1 = 32'd7887
; 
32'd154161: dataIn1 = 32'd7888
; 
32'd154162: dataIn1 = 32'd8053
; 
32'd154163: dataIn1 = 32'd8054
; 
32'd154164: dataIn1 = 32'd5192
; 
32'd154165: dataIn1 = 32'd6318
; 
32'd154166: dataIn1 = 32'd6319
; 
32'd154167: dataIn1 = 32'd6321
; 
32'd154168: dataIn1 = 32'd6322
; 
32'd154169: dataIn1 = 32'd6708
; 
32'd154170: dataIn1 = 32'd6709
; 
32'd154171: dataIn1 = 32'd5193
; 
32'd154172: dataIn1 = 32'd7893
; 
32'd154173: dataIn1 = 32'd7894
; 
32'd154174: dataIn1 = 32'd7907
; 
32'd154175: dataIn1 = 32'd7914
; 
32'd154176: dataIn1 = 32'd8068
; 
32'd154177: dataIn1 = 32'd8069
; 
32'd154178: dataIn1 = 32'd5194
; 
32'd154179: dataIn1 = 32'd7897
; 
32'd154180: dataIn1 = 32'd7898
; 
32'd154181: dataIn1 = 32'd7903
; 
32'd154182: dataIn1 = 32'd7910
; 
32'd154183: dataIn1 = 32'd7986
; 
32'd154184: dataIn1 = 32'd7987
; 
32'd154185: dataIn1 = 32'd5195
; 
32'd154186: dataIn1 = 32'd6334
; 
32'd154187: dataIn1 = 32'd6335
; 
32'd154188: dataIn1 = 32'd6337
; 
32'd154189: dataIn1 = 32'd6338
; 
32'd154190: dataIn1 = 32'd6710
; 
32'd154191: dataIn1 = 32'd6711
; 
32'd154192: dataIn1 = 32'd5196
; 
32'd154193: dataIn1 = 32'd6336
; 
32'd154194: dataIn1 = 32'd6338
; 
32'd154195: dataIn1 = 32'd7920
; 
32'd154196: dataIn1 = 32'd7921
; 
32'd154197: dataIn1 = 32'd8006
; 
32'd154198: dataIn1 = 32'd8007
; 
32'd154199: dataIn1 = 32'd5197
; 
32'd154200: dataIn1 = 32'd7926
; 
32'd154201: dataIn1 = 32'd7927
; 
32'd154202: dataIn1 = 32'd7942
; 
32'd154203: dataIn1 = 32'd7949
; 
32'd154204: dataIn1 = 32'd7956
; 
32'd154205: dataIn1 = 32'd7957
; 
32'd154206: dataIn1 = 32'd5198
; 
32'd154207: dataIn1 = 32'd7928
; 
32'd154208: dataIn1 = 32'd7929
; 
32'd154209: dataIn1 = 32'd7937
; 
32'd154210: dataIn1 = 32'd7950
; 
32'd154211: dataIn1 = 32'd7984
; 
32'd154212: dataIn1 = 32'd7985
; 
32'd154213: dataIn1 = 32'd5199
; 
32'd154214: dataIn1 = 32'd7930
; 
32'd154215: dataIn1 = 32'd7931
; 
32'd154216: dataIn1 = 32'd7938
; 
32'd154217: dataIn1 = 32'd7945
; 
32'd154218: dataIn1 = 32'd8008
; 
32'd154219: dataIn1 = 32'd8009
; 
32'd154220: dataIn1 = 32'd5200
; 
32'd154221: dataIn1 = 32'd7960
; 
32'd154222: dataIn1 = 32'd7961
; 
32'd154223: dataIn1 = 32'd7968
; 
32'd154224: dataIn1 = 32'd7973
; 
32'd154225: dataIn1 = 32'd9056
; 
32'd154226: dataIn1 = 32'd9057
; 
32'd154227: dataIn1 = 32'd5201
; 
32'd154228: dataIn1 = 32'd6360
; 
32'd154229: dataIn1 = 32'd6638
; 
32'd154230: dataIn1 = 32'd8004
; 
32'd154231: dataIn1 = 32'd8005
; 
32'd154232: dataIn1 = 32'd8016
; 
32'd154233: dataIn1 = 32'd9072
; 
32'd154234: dataIn1 = 32'd5202
; 
32'd154235: dataIn1 = 32'd8021
; 
32'd154236: dataIn1 = 32'd8022
; 
32'd154237: dataIn1 = 32'd8037
; 
32'd154238: dataIn1 = 32'd8044
; 
32'd154239: dataIn1 = 32'd8051
; 
32'd154240: dataIn1 = 32'd8052
; 
32'd154241: dataIn1 = 32'd5203
; 
32'd154242: dataIn1 = 32'd8023
; 
32'd154243: dataIn1 = 32'd8024
; 
32'd154244: dataIn1 = 32'd8032
; 
32'd154245: dataIn1 = 32'd8045
; 
32'd154246: dataIn1 = 32'd8070
; 
32'd154247: dataIn1 = 32'd8071
; 
32'd154248: dataIn1 = 32'd5204
; 
32'd154249: dataIn1 = 32'd8025
; 
32'd154250: dataIn1 = 32'd8026
; 
32'd154251: dataIn1 = 32'd8033
; 
32'd154252: dataIn1 = 32'd8040
; 
32'd154253: dataIn1 = 32'd8094
; 
32'd154254: dataIn1 = 32'd8095
; 
32'd154255: dataIn1 = 32'd5205
; 
32'd154256: dataIn1 = 32'd6373
; 
32'd154257: dataIn1 = 32'd6660
; 
32'd154258: dataIn1 = 32'd8055
; 
32'd154259: dataIn1 = 32'd8056
; 
32'd154260: dataIn1 = 32'd8061
; 
32'd154261: dataIn1 = 32'd9128
; 
32'd154262: dataIn1 = 32'd5206
; 
32'd154263: dataIn1 = 32'd8090
; 
32'd154264: dataIn1 = 32'd8091
; 
32'd154265: dataIn1 = 32'd8104
; 
32'd154266: dataIn1 = 32'd8109
; 
32'd154267: dataIn1 = 32'd9109
; 
32'd154268: dataIn1 = 32'd9110
; 
32'd154269: dataIn1 = 32'd5207
; 
32'd154270: dataIn1 = 32'd6389
; 
32'd154271: dataIn1 = 32'd8116
; 
32'd154272: dataIn1 = 32'd8117
; 
32'd154273: dataIn1 = 32'd8132
; 
32'd154274: dataIn1 = 32'd8139
; 
32'd154275: dataIn1 = 32'd9765
; 
32'd154276: dataIn1 = 32'd5208
; 
32'd154277: dataIn1 = 32'd8118
; 
32'd154278: dataIn1 = 32'd8119
; 
32'd154279: dataIn1 = 32'd8127
; 
32'd154280: dataIn1 = 32'd8133
; 
32'd154281: dataIn1 = 32'd8148
; 
32'd154282: dataIn1 = 32'd8149
; 
32'd154283: dataIn1 = 32'd5209
; 
32'd154284: dataIn1 = 32'd6388
; 
32'd154285: dataIn1 = 32'd6408
; 
32'd154286: dataIn1 = 32'd8120
; 
32'd154287: dataIn1 = 32'd8121
; 
32'd154288: dataIn1 = 32'd8128
; 
32'd154289: dataIn1 = 32'd8175
; 
32'd154290: dataIn1 = 32'd5210
; 
32'd154291: dataIn1 = 32'd8140
; 
32'd154292: dataIn1 = 32'd8141
; 
32'd154293: dataIn1 = 32'd8306
; 
32'd154294: dataIn1 = 32'd8307
; 
32'd154295: dataIn1 = 32'd9766
; 
32'd154296: dataIn1 = 32'd10278
; 
32'd154297: dataIn1 = 32'd5211
; 
32'd154298: dataIn1 = 32'd6397
; 
32'd154299: dataIn1 = 32'd9738
; 
32'd154300: dataIn1 = 32'd9739
; 
32'd154301: dataIn1 = 32'd9740
; 
32'd154302: dataIn1 = 32'd9748
; 
32'd154303: dataIn1 = 32'd10221
; 
32'd154304: dataIn1 = 32'd5212
; 
32'd154305: dataIn1 = 32'd8146
; 
32'd154306: dataIn1 = 32'd8147
; 
32'd154307: dataIn1 = 32'd8160
; 
32'd154308: dataIn1 = 32'd8167
; 
32'd154309: dataIn1 = 32'd8320
; 
32'd154310: dataIn1 = 32'd8321
; 
32'd154311: dataIn1 = 32'd5213
; 
32'd154312: dataIn1 = 32'd8150
; 
32'd154313: dataIn1 = 32'd8151
; 
32'd154314: dataIn1 = 32'd8156
; 
32'd154315: dataIn1 = 32'd8163
; 
32'd154316: dataIn1 = 32'd8239
; 
32'd154317: dataIn1 = 32'd8240
; 
32'd154318: dataIn1 = 32'd5214
; 
32'd154319: dataIn1 = 32'd6408
; 
32'd154320: dataIn1 = 32'd6409
; 
32'd154321: dataIn1 = 32'd6714
; 
32'd154322: dataIn1 = 32'd6715
; 
32'd154323: dataIn1 = 32'd6716
; 
32'd154324: dataIn1 = 32'd9233
; 
32'd154325: dataIn1 = 32'd5215
; 
32'd154326: dataIn1 = 32'd6714
; 
32'd154327: dataIn1 = 32'd6764
; 
32'd154328: dataIn1 = 32'd8173
; 
32'd154329: dataIn1 = 32'd8174
; 
32'd154330: dataIn1 = 32'd8259
; 
32'd154331: dataIn1 = 32'd8260
; 
32'd154332: dataIn1 = 32'd5216
; 
32'd154333: dataIn1 = 32'd8179
; 
32'd154334: dataIn1 = 32'd8180
; 
32'd154335: dataIn1 = 32'd8195
; 
32'd154336: dataIn1 = 32'd8202
; 
32'd154337: dataIn1 = 32'd8209
; 
32'd154338: dataIn1 = 32'd8210
; 
32'd154339: dataIn1 = 32'd5217
; 
32'd154340: dataIn1 = 32'd8181
; 
32'd154341: dataIn1 = 32'd8182
; 
32'd154342: dataIn1 = 32'd8190
; 
32'd154343: dataIn1 = 32'd8203
; 
32'd154344: dataIn1 = 32'd8237
; 
32'd154345: dataIn1 = 32'd8238
; 
32'd154346: dataIn1 = 32'd5218
; 
32'd154347: dataIn1 = 32'd8183
; 
32'd154348: dataIn1 = 32'd8184
; 
32'd154349: dataIn1 = 32'd8191
; 
32'd154350: dataIn1 = 32'd8198
; 
32'd154351: dataIn1 = 32'd8261
; 
32'd154352: dataIn1 = 32'd8262
; 
32'd154353: dataIn1 = 32'd5219
; 
32'd154354: dataIn1 = 32'd8213
; 
32'd154355: dataIn1 = 32'd8214
; 
32'd154356: dataIn1 = 32'd8221
; 
32'd154357: dataIn1 = 32'd8226
; 
32'd154358: dataIn1 = 32'd9107
; 
32'd154359: dataIn1 = 32'd9108
; 
32'd154360: dataIn1 = 32'd5220
; 
32'd154361: dataIn1 = 32'd6725
; 
32'd154362: dataIn1 = 32'd6765
; 
32'd154363: dataIn1 = 32'd8257
; 
32'd154364: dataIn1 = 32'd8258
; 
32'd154365: dataIn1 = 32'd8269
; 
32'd154366: dataIn1 = 32'd9123
; 
32'd154367: dataIn1 = 32'd5221
; 
32'd154368: dataIn1 = 32'd8274
; 
32'd154369: dataIn1 = 32'd8275
; 
32'd154370: dataIn1 = 32'd8290
; 
32'd154371: dataIn1 = 32'd8297
; 
32'd154372: dataIn1 = 32'd8304
; 
32'd154373: dataIn1 = 32'd8305
; 
32'd154374: dataIn1 = 32'd5222
; 
32'd154375: dataIn1 = 32'd8276
; 
32'd154376: dataIn1 = 32'd8277
; 
32'd154377: dataIn1 = 32'd8285
; 
32'd154378: dataIn1 = 32'd8298
; 
32'd154379: dataIn1 = 32'd8322
; 
32'd154380: dataIn1 = 32'd8323
; 
32'd154381: dataIn1 = 32'd5223
; 
32'd154382: dataIn1 = 32'd8278
; 
32'd154383: dataIn1 = 32'd8279
; 
32'd154384: dataIn1 = 32'd8286
; 
32'd154385: dataIn1 = 32'd8293
; 
32'd154386: dataIn1 = 32'd8346
; 
32'd154387: dataIn1 = 32'd8347
; 
32'd154388: dataIn1 = 32'd5224
; 
32'd154389: dataIn1 = 32'd6443
; 
32'd154390: dataIn1 = 32'd6676
; 
32'd154391: dataIn1 = 32'd8308
; 
32'd154392: dataIn1 = 32'd8309
; 
32'd154393: dataIn1 = 32'd9275
; 
32'd154394: dataIn1 = 32'd9285
; 
32'd154395: dataIn1 = 32'd5225
; 
32'd154396: dataIn1 = 32'd8342
; 
32'd154397: dataIn1 = 32'd8343
; 
32'd154398: dataIn1 = 32'd8356
; 
32'd154399: dataIn1 = 32'd8361
; 
32'd154400: dataIn1 = 32'd9161
; 
32'd154401: dataIn1 = 32'd9162
; 
32'd154402: dataIn1 = 32'd5226
; 
32'd154403: dataIn1 = 32'd6767
; 
32'd154404: dataIn1 = 32'd6769
; 
32'd154405: dataIn1 = 32'd8368
; 
32'd154406: dataIn1 = 32'd8369
; 
32'd154407: dataIn1 = 32'd8384
; 
32'd154408: dataIn1 = 32'd8391
; 
32'd154409: dataIn1 = 32'd5227
; 
32'd154410: dataIn1 = 32'd8370
; 
32'd154411: dataIn1 = 32'd8371
; 
32'd154412: dataIn1 = 32'd8379
; 
32'd154413: dataIn1 = 32'd8385
; 
32'd154414: dataIn1 = 32'd8400
; 
32'd154415: dataIn1 = 32'd8401
; 
32'd154416: dataIn1 = 32'd5228
; 
32'd154417: dataIn1 = 32'd6766
; 
32'd154418: dataIn1 = 32'd6770
; 
32'd154419: dataIn1 = 32'd8372
; 
32'd154420: dataIn1 = 32'd8373
; 
32'd154421: dataIn1 = 32'd8380
; 
32'd154422: dataIn1 = 32'd8427
; 
32'd154423: dataIn1 = 32'd5229
; 
32'd154424: dataIn1 = 32'd6768
; 
32'd154425: dataIn1 = 32'd6775
; 
32'd154426: dataIn1 = 32'd8392
; 
32'd154427: dataIn1 = 32'd8393
; 
32'd154428: dataIn1 = 32'd8558
; 
32'd154429: dataIn1 = 32'd8559
; 
32'd154430: dataIn1 = 32'd5230
; 
32'd154431: dataIn1 = 32'd6768
; 
32'd154432: dataIn1 = 32'd6769
; 
32'd154433: dataIn1 = 32'd9246
; 
32'd154434: dataIn1 = 32'd9248
; 
32'd154435: dataIn1 = 32'd9299
; 
32'd154436: dataIn1 = 32'd9300
; 
32'd154437: dataIn1 = 32'd5231
; 
32'd154438: dataIn1 = 32'd8398
; 
32'd154439: dataIn1 = 32'd8399
; 
32'd154440: dataIn1 = 32'd8412
; 
32'd154441: dataIn1 = 32'd8419
; 
32'd154442: dataIn1 = 32'd8573
; 
32'd154443: dataIn1 = 32'd8574
; 
32'd154444: dataIn1 = 32'd5232
; 
32'd154445: dataIn1 = 32'd8402
; 
32'd154446: dataIn1 = 32'd8403
; 
32'd154447: dataIn1 = 32'd8408
; 
32'd154448: dataIn1 = 32'd8415
; 
32'd154449: dataIn1 = 32'd8491
; 
32'd154450: dataIn1 = 32'd8492
; 
32'd154451: dataIn1 = 32'd5233
; 
32'd154452: dataIn1 = 32'd6770
; 
32'd154453: dataIn1 = 32'd6771
; 
32'd154454: dataIn1 = 32'd9247
; 
32'd154455: dataIn1 = 32'd9249
; 
32'd154456: dataIn1 = 32'd9301
; 
32'd154457: dataIn1 = 32'd9302
; 
32'd154458: dataIn1 = 32'd5234
; 
32'd154459: dataIn1 = 32'd6771
; 
32'd154460: dataIn1 = 32'd6772
; 
32'd154461: dataIn1 = 32'd8425
; 
32'd154462: dataIn1 = 32'd8426
; 
32'd154463: dataIn1 = 32'd8511
; 
32'd154464: dataIn1 = 32'd8512
; 
32'd154465: dataIn1 = 32'd5235
; 
32'd154466: dataIn1 = 32'd8431
; 
32'd154467: dataIn1 = 32'd8432
; 
32'd154468: dataIn1 = 32'd8447
; 
32'd154469: dataIn1 = 32'd8454
; 
32'd154470: dataIn1 = 32'd8461
; 
32'd154471: dataIn1 = 32'd8462
; 
32'd154472: dataIn1 = 32'd5236
; 
32'd154473: dataIn1 = 32'd8433
; 
32'd154474: dataIn1 = 32'd8434
; 
32'd154475: dataIn1 = 32'd8442
; 
32'd154476: dataIn1 = 32'd8455
; 
32'd154477: dataIn1 = 32'd8489
; 
32'd154478: dataIn1 = 32'd8490
; 
32'd154479: dataIn1 = 32'd5237
; 
32'd154480: dataIn1 = 32'd8435
; 
32'd154481: dataIn1 = 32'd8436
; 
32'd154482: dataIn1 = 32'd8443
; 
32'd154483: dataIn1 = 32'd8450
; 
32'd154484: dataIn1 = 32'd8513
; 
32'd154485: dataIn1 = 32'd8514
; 
32'd154486: dataIn1 = 32'd5238
; 
32'd154487: dataIn1 = 32'd8465
; 
32'd154488: dataIn1 = 32'd8466
; 
32'd154489: dataIn1 = 32'd8473
; 
32'd154490: dataIn1 = 32'd8478
; 
32'd154491: dataIn1 = 32'd9159
; 
32'd154492: dataIn1 = 32'd9160
; 
32'd154493: dataIn1 = 32'd5239
; 
32'd154494: dataIn1 = 32'd6773
; 
32'd154495: dataIn1 = 32'd6795
; 
32'd154496: dataIn1 = 32'd8509
; 
32'd154497: dataIn1 = 32'd8510
; 
32'd154498: dataIn1 = 32'd8521
; 
32'd154499: dataIn1 = 32'd9175
; 
32'd154500: dataIn1 = 32'd5240
; 
32'd154501: dataIn1 = 32'd8526
; 
32'd154502: dataIn1 = 32'd8527
; 
32'd154503: dataIn1 = 32'd8542
; 
32'd154504: dataIn1 = 32'd8549
; 
32'd154505: dataIn1 = 32'd8556
; 
32'd154506: dataIn1 = 32'd8557
; 
32'd154507: dataIn1 = 32'd5241
; 
32'd154508: dataIn1 = 32'd8528
; 
32'd154509: dataIn1 = 32'd8529
; 
32'd154510: dataIn1 = 32'd8537
; 
32'd154511: dataIn1 = 32'd8550
; 
32'd154512: dataIn1 = 32'd8575
; 
32'd154513: dataIn1 = 32'd8576
; 
32'd154514: dataIn1 = 32'd5242
; 
32'd154515: dataIn1 = 32'd8530
; 
32'd154516: dataIn1 = 32'd8531
; 
32'd154517: dataIn1 = 32'd8538
; 
32'd154518: dataIn1 = 32'd8545
; 
32'd154519: dataIn1 = 32'd8599
; 
32'd154520: dataIn1 = 32'd8600
; 
32'd154521: dataIn1 = 32'd5243
; 
32'd154522: dataIn1 = 32'd6774
; 
32'd154523: dataIn1 = 32'd6801
; 
32'd154524: dataIn1 = 32'd8560
; 
32'd154525: dataIn1 = 32'd8561
; 
32'd154526: dataIn1 = 32'd8566
; 
32'd154527: dataIn1 = 32'd9230
; 
32'd154528: dataIn1 = 32'd5244
; 
32'd154529: dataIn1 = 32'd8595
; 
32'd154530: dataIn1 = 32'd8596
; 
32'd154531: dataIn1 = 32'd8609
; 
32'd154532: dataIn1 = 32'd8614
; 
32'd154533: dataIn1 = 32'd9211
; 
32'd154534: dataIn1 = 32'd9212
; 
32'd154535: dataIn1 = 32'd5245
; 
32'd154536: dataIn1 = 32'd6777
; 
32'd154537: dataIn1 = 32'd6779
; 
32'd154538: dataIn1 = 32'd8621
; 
32'd154539: dataIn1 = 32'd8622
; 
32'd154540: dataIn1 = 32'd8637
; 
32'd154541: dataIn1 = 32'd8644
; 
32'd154542: dataIn1 = 32'd5246
; 
32'd154543: dataIn1 = 32'd8623
; 
32'd154544: dataIn1 = 32'd8624
; 
32'd154545: dataIn1 = 32'd8632
; 
32'd154546: dataIn1 = 32'd8638
; 
32'd154547: dataIn1 = 32'd8653
; 
32'd154548: dataIn1 = 32'd8654
; 
32'd154549: dataIn1 = 32'd5247
; 
32'd154550: dataIn1 = 32'd6776
; 
32'd154551: dataIn1 = 32'd6780
; 
32'd154552: dataIn1 = 32'd8625
; 
32'd154553: dataIn1 = 32'd8626
; 
32'd154554: dataIn1 = 32'd8633
; 
32'd154555: dataIn1 = 32'd8680
; 
32'd154556: dataIn1 = 32'd5248
; 
32'd154557: dataIn1 = 32'd6778
; 
32'd154558: dataIn1 = 32'd6785
; 
32'd154559: dataIn1 = 32'd8645
; 
32'd154560: dataIn1 = 32'd8646
; 
32'd154561: dataIn1 = 32'd8811
; 
32'd154562: dataIn1 = 32'd8812
; 
32'd154563: dataIn1 = 32'd5249
; 
32'd154564: dataIn1 = 32'd6778
; 
32'd154565: dataIn1 = 32'd6779
; 
32'd154566: dataIn1 = 32'd9252
; 
32'd154567: dataIn1 = 32'd9254
; 
32'd154568: dataIn1 = 32'd9305
; 
32'd154569: dataIn1 = 32'd9306
; 
32'd154570: dataIn1 = 32'd5250
; 
32'd154571: dataIn1 = 32'd8651
; 
32'd154572: dataIn1 = 32'd8652
; 
32'd154573: dataIn1 = 32'd8665
; 
32'd154574: dataIn1 = 32'd8672
; 
32'd154575: dataIn1 = 32'd8825
; 
32'd154576: dataIn1 = 32'd8826
; 
32'd154577: dataIn1 = 32'd5251
; 
32'd154578: dataIn1 = 32'd8655
; 
32'd154579: dataIn1 = 32'd8656
; 
32'd154580: dataIn1 = 32'd8661
; 
32'd154581: dataIn1 = 32'd8668
; 
32'd154582: dataIn1 = 32'd8744
; 
32'd154583: dataIn1 = 32'd8745
; 
32'd154584: dataIn1 = 32'd5252
; 
32'd154585: dataIn1 = 32'd6780
; 
32'd154586: dataIn1 = 32'd6781
; 
32'd154587: dataIn1 = 32'd9253
; 
32'd154588: dataIn1 = 32'd9255
; 
32'd154589: dataIn1 = 32'd9307
; 
32'd154590: dataIn1 = 32'd9308
; 
32'd154591: dataIn1 = 32'd5253
; 
32'd154592: dataIn1 = 32'd6781
; 
32'd154593: dataIn1 = 32'd6782
; 
32'd154594: dataIn1 = 32'd8678
; 
32'd154595: dataIn1 = 32'd8679
; 
32'd154596: dataIn1 = 32'd8764
; 
32'd154597: dataIn1 = 32'd8765
; 
32'd154598: dataIn1 = 32'd5254
; 
32'd154599: dataIn1 = 32'd8684
; 
32'd154600: dataIn1 = 32'd8685
; 
32'd154601: dataIn1 = 32'd8700
; 
32'd154602: dataIn1 = 32'd8707
; 
32'd154603: dataIn1 = 32'd8714
; 
32'd154604: dataIn1 = 32'd8715
; 
32'd154605: dataIn1 = 32'd5255
; 
32'd154606: dataIn1 = 32'd8686
; 
32'd154607: dataIn1 = 32'd8687
; 
32'd154608: dataIn1 = 32'd8695
; 
32'd154609: dataIn1 = 32'd8708
; 
32'd154610: dataIn1 = 32'd8742
; 
32'd154611: dataIn1 = 32'd8743
; 
32'd154612: dataIn1 = 32'd5256
; 
32'd154613: dataIn1 = 32'd8688
; 
32'd154614: dataIn1 = 32'd8689
; 
32'd154615: dataIn1 = 32'd8696
; 
32'd154616: dataIn1 = 32'd8703
; 
32'd154617: dataIn1 = 32'd8766
; 
32'd154618: dataIn1 = 32'd8767
; 
32'd154619: dataIn1 = 32'd5257
; 
32'd154620: dataIn1 = 32'd8718
; 
32'd154621: dataIn1 = 32'd8719
; 
32'd154622: dataIn1 = 32'd8726
; 
32'd154623: dataIn1 = 32'd8731
; 
32'd154624: dataIn1 = 32'd9209
; 
32'd154625: dataIn1 = 32'd9210
; 
32'd154626: dataIn1 = 32'd5258
; 
32'd154627: dataIn1 = 32'd6783
; 
32'd154628: dataIn1 = 32'd6799
; 
32'd154629: dataIn1 = 32'd8762
; 
32'd154630: dataIn1 = 32'd8763
; 
32'd154631: dataIn1 = 32'd8774
; 
32'd154632: dataIn1 = 32'd9225
; 
32'd154633: dataIn1 = 32'd5259
; 
32'd154634: dataIn1 = 32'd8779
; 
32'd154635: dataIn1 = 32'd8780
; 
32'd154636: dataIn1 = 32'd8795
; 
32'd154637: dataIn1 = 32'd8802
; 
32'd154638: dataIn1 = 32'd8809
; 
32'd154639: dataIn1 = 32'd8810
; 
32'd154640: dataIn1 = 32'd5260
; 
32'd154641: dataIn1 = 32'd8781
; 
32'd154642: dataIn1 = 32'd8782
; 
32'd154643: dataIn1 = 32'd8790
; 
32'd154644: dataIn1 = 32'd8803
; 
32'd154645: dataIn1 = 32'd8827
; 
32'd154646: dataIn1 = 32'd8828
; 
32'd154647: dataIn1 = 32'd5261
; 
32'd154648: dataIn1 = 32'd8783
; 
32'd154649: dataIn1 = 32'd8784
; 
32'd154650: dataIn1 = 32'd8791
; 
32'd154651: dataIn1 = 32'd8798
; 
32'd154652: dataIn1 = 32'd8851
; 
32'd154653: dataIn1 = 32'd8852
; 
32'd154654: dataIn1 = 32'd5262
; 
32'd154655: dataIn1 = 32'd6784
; 
32'd154656: dataIn1 = 32'd6849
; 
32'd154657: dataIn1 = 32'd8813
; 
32'd154658: dataIn1 = 32'd8814
; 
32'd154659: dataIn1 = 32'd8818
; 
32'd154660: dataIn1 = 32'd9447
; 
32'd154661: dataIn1 = 32'd5263
; 
32'd154662: dataIn1 = 32'd8847
; 
32'd154663: dataIn1 = 32'd8848
; 
32'd154664: dataIn1 = 32'd8861
; 
32'd154665: dataIn1 = 32'd8866
; 
32'd154666: dataIn1 = 32'd9421
; 
32'd154667: dataIn1 = 32'd9422
; 
32'd154668: dataIn1 = 32'd5264
; 
32'd154669: dataIn1 = 32'd8873
; 
32'd154670: dataIn1 = 32'd8874
; 
32'd154671: dataIn1 = 32'd8882
; 
32'd154672: dataIn1 = 32'd8889
; 
32'd154673: dataIn1 = 32'd8896
; 
32'd154674: dataIn1 = 32'd8897
; 
32'd154675: dataIn1 = 32'd5265
; 
32'd154676: dataIn1 = 32'd6577
; 
32'd154677: dataIn1 = 32'd6585
; 
32'd154678: dataIn1 = 32'd8875
; 
32'd154679: dataIn1 = 32'd8876
; 
32'd154680: dataIn1 = 32'd8890
; 
32'd154681: dataIn1 = 32'd8915
; 
32'd154682: dataIn1 = 32'd5266
; 
32'd154683: dataIn1 = 32'd6576
; 
32'd154684: dataIn1 = 32'd6590
; 
32'd154685: dataIn1 = 32'd8877
; 
32'd154686: dataIn1 = 32'd8878
; 
32'd154687: dataIn1 = 32'd8885
; 
32'd154688: dataIn1 = 32'd8920
; 
32'd154689: dataIn1 = 32'd5267
; 
32'd154690: dataIn1 = 32'd6585
; 
32'd154691: dataIn1 = 32'd6586
; 
32'd154692: dataIn1 = 32'd6588
; 
32'd154693: dataIn1 = 32'd6589
; 
32'd154694: dataIn1 = 32'd6717
; 
32'd154695: dataIn1 = 32'd6718
; 
32'd154696: dataIn1 = 32'd5268
; 
32'd154697: dataIn1 = 32'd6590
; 
32'd154698: dataIn1 = 32'd6592
; 
32'd154699: dataIn1 = 32'd6593
; 
32'd154700: dataIn1 = 32'd6594
; 
32'd154701: dataIn1 = 32'd6719
; 
32'd154702: dataIn1 = 32'd6720
; 
32'd154703: dataIn1 = 32'd5269
; 
32'd154704: dataIn1 = 32'd5270
; 
32'd154705: dataIn1 = 32'd5271
; 
32'd154706: dataIn1 = 32'd6596
; 
32'd154707: dataIn1 = 32'd6597
; 
32'd154708: dataIn1 = 32'd6598
; 
32'd154709: dataIn1 = 32'd9671
; 
32'd154710: dataIn1 = 32'd9742
; 
32'd154711: dataIn1 = 32'd2700
; 
32'd154712: dataIn1 = 32'd2738
; 
32'd154713: dataIn1 = 32'd5144
; 
32'd154714: dataIn1 = 32'd5269
; 
32'd154715: dataIn1 = 32'd5270
; 
32'd154716: dataIn1 = 32'd5271
; 
32'd154717: dataIn1 = 32'd5272
; 
32'd154718: dataIn1 = 32'd9671
; 
32'd154719: dataIn1 = 32'd2325
; 
32'd154720: dataIn1 = 32'd2738
; 
32'd154721: dataIn1 = 32'd3984
; 
32'd154722: dataIn1 = 32'd5269
; 
32'd154723: dataIn1 = 32'd5270
; 
32'd154724: dataIn1 = 32'd5271
; 
32'd154725: dataIn1 = 32'd5273
; 
32'd154726: dataIn1 = 32'd6598
; 
32'd154727: dataIn1 = 32'd9272
; 
32'd154728: dataIn1 = 32'd1122
; 
32'd154729: dataIn1 = 32'd2738
; 
32'd154730: dataIn1 = 32'd2740
; 
32'd154731: dataIn1 = 32'd5144
; 
32'd154732: dataIn1 = 32'd5270
; 
32'd154733: dataIn1 = 32'd5272
; 
32'd154734: dataIn1 = 32'd451
; 
32'd154735: dataIn1 = 32'd2738
; 
32'd154736: dataIn1 = 32'd3984
; 
32'd154737: dataIn1 = 32'd5271
; 
32'd154738: dataIn1 = 32'd5273
; 
32'd154739: dataIn1 = 32'd5633
; 
32'd154740: dataIn1 = 32'd5634
; 
32'd154741: dataIn1 = 32'd5274
; 
32'd154742: dataIn1 = 32'd8930
; 
32'd154743: dataIn1 = 32'd8931
; 
32'd154744: dataIn1 = 32'd8939
; 
32'd154745: dataIn1 = 32'd8946
; 
32'd154746: dataIn1 = 32'd8953
; 
32'd154747: dataIn1 = 32'd8954
; 
32'd154748: dataIn1 = 32'd5275
; 
32'd154749: dataIn1 = 32'd8932
; 
32'd154750: dataIn1 = 32'd8933
; 
32'd154751: dataIn1 = 32'd8947
; 
32'd154752: dataIn1 = 32'd8974
; 
32'd154753: dataIn1 = 32'd9278
; 
32'd154754: dataIn1 = 32'd9279
; 
32'd154755: dataIn1 = 32'd5276
; 
32'd154756: dataIn1 = 32'd5278
; 
32'd154757: dataIn1 = 32'd6610
; 
32'd154758: dataIn1 = 32'd8934
; 
32'd154759: dataIn1 = 32'd8935
; 
32'd154760: dataIn1 = 32'd8942
; 
32'd154761: dataIn1 = 32'd9277
; 
32'd154762: dataIn1 = 32'd5277
; 
32'd154763: dataIn1 = 32'd9279
; 
32'd154764: dataIn1 = 32'd9280
; 
32'd154765: dataIn1 = 32'd9321
; 
32'd154766: dataIn1 = 32'd9322
; 
32'd154767: dataIn1 = 32'd9337
; 
32'd154768: dataIn1 = 32'd9338
; 
32'd154769: dataIn1 = 32'd1121
; 
32'd154770: dataIn1 = 32'd2743
; 
32'd154771: dataIn1 = 32'd2744
; 
32'd154772: dataIn1 = 32'd5148
; 
32'd154773: dataIn1 = 32'd5276
; 
32'd154774: dataIn1 = 32'd5278
; 
32'd154775: dataIn1 = 32'd6610
; 
32'd154776: dataIn1 = 32'd9277
; 
32'd154777: dataIn1 = 32'd5279
; 
32'd154778: dataIn1 = 32'd8979
; 
32'd154779: dataIn1 = 32'd8980
; 
32'd154780: dataIn1 = 32'd8988
; 
32'd154781: dataIn1 = 32'd8995
; 
32'd154782: dataIn1 = 32'd9002
; 
32'd154783: dataIn1 = 32'd9003
; 
32'd154784: dataIn1 = 32'd5280
; 
32'd154785: dataIn1 = 32'd6787
; 
32'd154786: dataIn1 = 32'd6788
; 
32'd154787: dataIn1 = 32'd8981
; 
32'd154788: dataIn1 = 32'd8982
; 
32'd154789: dataIn1 = 32'd8996
; 
32'd154790: dataIn1 = 32'd9021
; 
32'd154791: dataIn1 = 32'd5281
; 
32'd154792: dataIn1 = 32'd6786
; 
32'd154793: dataIn1 = 32'd6790
; 
32'd154794: dataIn1 = 32'd8983
; 
32'd154795: dataIn1 = 32'd8984
; 
32'd154796: dataIn1 = 32'd8991
; 
32'd154797: dataIn1 = 32'd9026
; 
32'd154798: dataIn1 = 32'd5282
; 
32'd154799: dataIn1 = 32'd6788
; 
32'd154800: dataIn1 = 32'd6789
; 
32'd154801: dataIn1 = 32'd9244
; 
32'd154802: dataIn1 = 32'd9258
; 
32'd154803: dataIn1 = 32'd9297
; 
32'd154804: dataIn1 = 32'd9298
; 
32'd154805: dataIn1 = 32'd5283
; 
32'd154806: dataIn1 = 32'd6790
; 
32'd154807: dataIn1 = 32'd6791
; 
32'd154808: dataIn1 = 32'd9239
; 
32'd154809: dataIn1 = 32'd9259
; 
32'd154810: dataIn1 = 32'd9291
; 
32'd154811: dataIn1 = 32'd9292
; 
32'd154812: dataIn1 = 32'd5284
; 
32'd154813: dataIn1 = 32'd9030
; 
32'd154814: dataIn1 = 32'd9031
; 
32'd154815: dataIn1 = 32'd9040
; 
32'd154816: dataIn1 = 32'd9047
; 
32'd154817: dataIn1 = 32'd9054
; 
32'd154818: dataIn1 = 32'd9055
; 
32'd154819: dataIn1 = 32'd5285
; 
32'd154820: dataIn1 = 32'd6627
; 
32'd154821: dataIn1 = 32'd6635
; 
32'd154822: dataIn1 = 32'd9032
; 
32'd154823: dataIn1 = 32'd9033
; 
32'd154824: dataIn1 = 32'd9048
; 
32'd154825: dataIn1 = 32'd9073
; 
32'd154826: dataIn1 = 32'd5286
; 
32'd154827: dataIn1 = 32'd6626
; 
32'd154828: dataIn1 = 32'd6792
; 
32'd154829: dataIn1 = 32'd9034
; 
32'd154830: dataIn1 = 32'd9035
; 
32'd154831: dataIn1 = 32'd9043
; 
32'd154832: dataIn1 = 32'd9078
; 
32'd154833: dataIn1 = 32'd5287
; 
32'd154834: dataIn1 = 32'd6635
; 
32'd154835: dataIn1 = 32'd6636
; 
32'd154836: dataIn1 = 32'd6637
; 
32'd154837: dataIn1 = 32'd6638
; 
32'd154838: dataIn1 = 32'd6721
; 
32'd154839: dataIn1 = 32'd6722
; 
32'd154840: dataIn1 = 32'd5288
; 
32'd154841: dataIn1 = 32'd6792
; 
32'd154842: dataIn1 = 32'd6793
; 
32'd154843: dataIn1 = 32'd9036
; 
32'd154844: dataIn1 = 32'd9245
; 
32'd154845: dataIn1 = 32'd9281
; 
32'd154846: dataIn1 = 32'd9282
; 
32'd154847: dataIn1 = 32'd5289
; 
32'd154848: dataIn1 = 32'd9082
; 
32'd154849: dataIn1 = 32'd9083
; 
32'd154850: dataIn1 = 32'd9091
; 
32'd154851: dataIn1 = 32'd9098
; 
32'd154852: dataIn1 = 32'd9105
; 
32'd154853: dataIn1 = 32'd9106
; 
32'd154854: dataIn1 = 32'd5290
; 
32'd154855: dataIn1 = 32'd6645
; 
32'd154856: dataIn1 = 32'd6653
; 
32'd154857: dataIn1 = 32'd9084
; 
32'd154858: dataIn1 = 32'd9085
; 
32'd154859: dataIn1 = 32'd9099
; 
32'd154860: dataIn1 = 32'd9124
; 
32'd154861: dataIn1 = 32'd5291
; 
32'd154862: dataIn1 = 32'd6644
; 
32'd154863: dataIn1 = 32'd6656
; 
32'd154864: dataIn1 = 32'd9086
; 
32'd154865: dataIn1 = 32'd9087
; 
32'd154866: dataIn1 = 32'd9094
; 
32'd154867: dataIn1 = 32'd9129
; 
32'd154868: dataIn1 = 32'd5292
; 
32'd154869: dataIn1 = 32'd6653
; 
32'd154870: dataIn1 = 32'd6654
; 
32'd154871: dataIn1 = 32'd6723
; 
32'd154872: dataIn1 = 32'd6724
; 
32'd154873: dataIn1 = 32'd6725
; 
32'd154874: dataIn1 = 32'd9234
; 
32'd154875: dataIn1 = 32'd5293
; 
32'd154876: dataIn1 = 32'd6656
; 
32'd154877: dataIn1 = 32'd6657
; 
32'd154878: dataIn1 = 32'd6659
; 
32'd154879: dataIn1 = 32'd6660
; 
32'd154880: dataIn1 = 32'd6726
; 
32'd154881: dataIn1 = 32'd6727
; 
32'd154882: dataIn1 = 32'd5294
; 
32'd154883: dataIn1 = 32'd9133
; 
32'd154884: dataIn1 = 32'd9134
; 
32'd154885: dataIn1 = 32'd9143
; 
32'd154886: dataIn1 = 32'd9150
; 
32'd154887: dataIn1 = 32'd9157
; 
32'd154888: dataIn1 = 32'd9158
; 
32'd154889: dataIn1 = 32'd5295
; 
32'd154890: dataIn1 = 32'd6665
; 
32'd154891: dataIn1 = 32'd6794
; 
32'd154892: dataIn1 = 32'd9135
; 
32'd154893: dataIn1 = 32'd9136
; 
32'd154894: dataIn1 = 32'd9151
; 
32'd154895: dataIn1 = 32'd9176
; 
32'd154896: dataIn1 = 32'd5296
; 
32'd154897: dataIn1 = 32'd6664
; 
32'd154898: dataIn1 = 32'd6674
; 
32'd154899: dataIn1 = 32'd9137
; 
32'd154900: dataIn1 = 32'd9138
; 
32'd154901: dataIn1 = 32'd9146
; 
32'd154902: dataIn1 = 32'd9180
; 
32'd154903: dataIn1 = 32'd5297
; 
32'd154904: dataIn1 = 32'd6794
; 
32'd154905: dataIn1 = 32'd6795
; 
32'd154906: dataIn1 = 32'd9139
; 
32'd154907: dataIn1 = 32'd9250
; 
32'd154908: dataIn1 = 32'd9283
; 
32'd154909: dataIn1 = 32'd9284
; 
32'd154910: dataIn1 = 32'd5298
; 
32'd154911: dataIn1 = 32'd6674
; 
32'd154912: dataIn1 = 32'd6676
; 
32'd154913: dataIn1 = 32'd6677
; 
32'd154914: dataIn1 = 32'd6678
; 
32'd154915: dataIn1 = 32'd6729
; 
32'd154916: dataIn1 = 32'd10246
; 
32'd154917: dataIn1 = 32'd5299
; 
32'd154918: dataIn1 = 32'd9184
; 
32'd154919: dataIn1 = 32'd9185
; 
32'd154920: dataIn1 = 32'd9193
; 
32'd154921: dataIn1 = 32'd9200
; 
32'd154922: dataIn1 = 32'd9207
; 
32'd154923: dataIn1 = 32'd9208
; 
32'd154924: dataIn1 = 32'd5300
; 
32'd154925: dataIn1 = 32'd6797
; 
32'd154926: dataIn1 = 32'd6798
; 
32'd154927: dataIn1 = 32'd9186
; 
32'd154928: dataIn1 = 32'd9187
; 
32'd154929: dataIn1 = 32'd9201
; 
32'd154930: dataIn1 = 32'd9226
; 
32'd154931: dataIn1 = 32'd5301
; 
32'd154932: dataIn1 = 32'd6796
; 
32'd154933: dataIn1 = 32'd6800
; 
32'd154934: dataIn1 = 32'd9188
; 
32'd154935: dataIn1 = 32'd9189
; 
32'd154936: dataIn1 = 32'd9196
; 
32'd154937: dataIn1 = 32'd9231
; 
32'd154938: dataIn1 = 32'd5302
; 
32'd154939: dataIn1 = 32'd6798
; 
32'd154940: dataIn1 = 32'd6799
; 
32'd154941: dataIn1 = 32'd9256
; 
32'd154942: dataIn1 = 32'd9260
; 
32'd154943: dataIn1 = 32'd9309
; 
32'd154944: dataIn1 = 32'd9310
; 
32'd154945: dataIn1 = 32'd5303
; 
32'd154946: dataIn1 = 32'd6800
; 
32'd154947: dataIn1 = 32'd6801
; 
32'd154948: dataIn1 = 32'd9251
; 
32'd154949: dataIn1 = 32'd9261
; 
32'd154950: dataIn1 = 32'd9303
; 
32'd154951: dataIn1 = 32'd9304
; 
32'd154952: dataIn1 = 32'd285
; 
32'd154953: dataIn1 = 32'd2295
; 
32'd154954: dataIn1 = 32'd2769
; 
32'd154955: dataIn1 = 32'd3421
; 
32'd154956: dataIn1 = 32'd3868
; 
32'd154957: dataIn1 = 32'd5304
; 
32'd154958: dataIn1 = 32'd193
; 
32'd154959: dataIn1 = 32'd2479
; 
32'd154960: dataIn1 = 32'd3401
; 
32'd154961: dataIn1 = 32'd4595
; 
32'd154962: dataIn1 = 32'd5305
; 
32'd154963: dataIn1 = 32'd2039
; 
32'd154964: dataIn1 = 32'd2533
; 
32'd154965: dataIn1 = 32'd2534
; 
32'd154966: dataIn1 = 32'd3408
; 
32'd154967: dataIn1 = 32'd4612
; 
32'd154968: dataIn1 = 32'd5306
; 
32'd154969: dataIn1 = 32'd980
; 
32'd154970: dataIn1 = 32'd2544
; 
32'd154971: dataIn1 = 32'd3417
; 
32'd154972: dataIn1 = 32'd4625
; 
32'd154973: dataIn1 = 32'd5307
; 
32'd154974: dataIn1 = 32'd5428
; 
32'd154975: dataIn1 = 32'd43
; 
32'd154976: dataIn1 = 32'd2154
; 
32'd154977: dataIn1 = 32'd2183
; 
32'd154978: dataIn1 = 32'd3606
; 
32'd154979: dataIn1 = 32'd3607
; 
32'd154980: dataIn1 = 32'd5308
; 
32'd154981: dataIn1 = 32'd54
; 
32'd154982: dataIn1 = 32'd2182
; 
32'd154983: dataIn1 = 32'd2212
; 
32'd154984: dataIn1 = 32'd3653
; 
32'd154985: dataIn1 = 32'd3654
; 
32'd154986: dataIn1 = 32'd5309
; 
32'd154987: dataIn1 = 32'd2215
; 
32'd154988: dataIn1 = 32'd2217
; 
32'd154989: dataIn1 = 32'd3658
; 
32'd154990: dataIn1 = 32'd3744
; 
32'd154991: dataIn1 = 32'd5310
; 
32'd154992: dataIn1 = 32'd9568
; 
32'd154993: dataIn1 = 32'd9773
; 
32'd154994: dataIn1 = 32'd9782
; 
32'd154995: dataIn1 = 32'd10204
; 
32'd154996: dataIn1 = 32'd74
; 
32'd154997: dataIn1 = 32'd75
; 
32'd154998: dataIn1 = 32'd85
; 
32'd154999: dataIn1 = 32'd2240
; 
32'd155000: dataIn1 = 32'd5311
; 
32'd155001: dataIn1 = 32'd5312
; 
32'd155002: dataIn1 = 32'd64
; 
32'd155003: dataIn1 = 32'd75
; 
32'd155004: dataIn1 = 32'd2213
; 
32'd155005: dataIn1 = 32'd2240
; 
32'd155006: dataIn1 = 32'd3731
; 
32'd155007: dataIn1 = 32'd5311
; 
32'd155008: dataIn1 = 32'd5312
; 
32'd155009: dataIn1 = 32'd5455
; 
32'd155010: dataIn1 = 32'd87
; 
32'd155011: dataIn1 = 32'd2266
; 
32'd155012: dataIn1 = 32'd2268
; 
32'd155013: dataIn1 = 32'd3826
; 
32'd155014: dataIn1 = 32'd3830
; 
32'd155015: dataIn1 = 32'd5313
; 
32'd155016: dataIn1 = 32'd88
; 
32'd155017: dataIn1 = 32'd98
; 
32'd155018: dataIn1 = 32'd2268
; 
32'd155019: dataIn1 = 32'd3829
; 
32'd155020: dataIn1 = 32'd5314
; 
32'd155021: dataIn1 = 32'd5315
; 
32'd155022: dataIn1 = 32'd5317
; 
32'd155023: dataIn1 = 32'd5456
; 
32'd155024: dataIn1 = 32'd87
; 
32'd155025: dataIn1 = 32'd97
; 
32'd155026: dataIn1 = 32'd98
; 
32'd155027: dataIn1 = 32'd2268
; 
32'd155028: dataIn1 = 32'd5314
; 
32'd155029: dataIn1 = 32'd5315
; 
32'd155030: dataIn1 = 32'd10288
; 
32'd155031: dataIn1 = 32'd89
; 
32'd155032: dataIn1 = 32'd99
; 
32'd155033: dataIn1 = 32'd100
; 
32'd155034: dataIn1 = 32'd2271
; 
32'd155035: dataIn1 = 32'd3841
; 
32'd155036: dataIn1 = 32'd5316
; 
32'd155037: dataIn1 = 32'd5317
; 
32'd155038: dataIn1 = 32'd10289
; 
32'd155039: dataIn1 = 32'd88
; 
32'd155040: dataIn1 = 32'd99
; 
32'd155041: dataIn1 = 32'd2271
; 
32'd155042: dataIn1 = 32'd3839
; 
32'd155043: dataIn1 = 32'd5314
; 
32'd155044: dataIn1 = 32'd5316
; 
32'd155045: dataIn1 = 32'd5317
; 
32'd155046: dataIn1 = 32'd5456
; 
32'd155047: dataIn1 = 32'd2302
; 
32'd155048: dataIn1 = 32'd2619
; 
32'd155049: dataIn1 = 32'd3898
; 
32'd155050: dataIn1 = 32'd4823
; 
32'd155051: dataIn1 = 32'd4838
; 
32'd155052: dataIn1 = 32'd5318
; 
32'd155053: dataIn1 = 32'd5430
; 
32'd155054: dataIn1 = 32'd5950
; 
32'd155055: dataIn1 = 32'd276
; 
32'd155056: dataIn1 = 32'd443
; 
32'd155057: dataIn1 = 32'd2310
; 
32'd155058: dataIn1 = 32'd3502
; 
32'd155059: dataIn1 = 32'd5319
; 
32'd155060: dataIn1 = 32'd5320
; 
32'd155061: dataIn1 = 32'd5457
; 
32'd155062: dataIn1 = 32'd276
; 
32'd155063: dataIn1 = 32'd448
; 
32'd155064: dataIn1 = 32'd2310
; 
32'd155065: dataIn1 = 32'd3931
; 
32'd155066: dataIn1 = 32'd5319
; 
32'd155067: dataIn1 = 32'd5320
; 
32'd155068: dataIn1 = 32'd5527
; 
32'd155069: dataIn1 = 32'd5528
; 
32'd155070: dataIn1 = 32'd284
; 
32'd155071: dataIn1 = 32'd450
; 
32'd155072: dataIn1 = 32'd2318
; 
32'd155073: dataIn1 = 32'd3961
; 
32'd155074: dataIn1 = 32'd5321
; 
32'd155075: dataIn1 = 32'd5322
; 
32'd155076: dataIn1 = 32'd5324
; 
32'd155077: dataIn1 = 32'd5458
; 
32'd155078: dataIn1 = 32'd284
; 
32'd155079: dataIn1 = 32'd448
; 
32'd155080: dataIn1 = 32'd2318
; 
32'd155081: dataIn1 = 32'd3959
; 
32'd155082: dataIn1 = 32'd5321
; 
32'd155083: dataIn1 = 32'd5322
; 
32'd155084: dataIn1 = 32'd5528
; 
32'd155085: dataIn1 = 32'd5529
; 
32'd155086: dataIn1 = 32'd451
; 
32'd155087: dataIn1 = 32'd2324
; 
32'd155088: dataIn1 = 32'd3967
; 
32'd155089: dataIn1 = 32'd3977
; 
32'd155090: dataIn1 = 32'd5323
; 
32'd155091: dataIn1 = 32'd5633
; 
32'd155092: dataIn1 = 32'd6691
; 
32'd155093: dataIn1 = 32'd153
; 
32'd155094: dataIn1 = 32'd450
; 
32'd155095: dataIn1 = 32'd2326
; 
32'd155096: dataIn1 = 32'd3994
; 
32'd155097: dataIn1 = 32'd5321
; 
32'd155098: dataIn1 = 32'd5324
; 
32'd155099: dataIn1 = 32'd5325
; 
32'd155100: dataIn1 = 32'd5458
; 
32'd155101: dataIn1 = 32'd153
; 
32'd155102: dataIn1 = 32'd453
; 
32'd155103: dataIn1 = 32'd2326
; 
32'd155104: dataIn1 = 32'd3992
; 
32'd155105: dataIn1 = 32'd5324
; 
32'd155106: dataIn1 = 32'd5325
; 
32'd155107: dataIn1 = 32'd5326
; 
32'd155108: dataIn1 = 32'd5459
; 
32'd155109: dataIn1 = 32'd283
; 
32'd155110: dataIn1 = 32'd453
; 
32'd155111: dataIn1 = 32'd2331
; 
32'd155112: dataIn1 = 32'd4007
; 
32'd155113: dataIn1 = 32'd5325
; 
32'd155114: dataIn1 = 32'd5326
; 
32'd155115: dataIn1 = 32'd5327
; 
32'd155116: dataIn1 = 32'd5459
; 
32'd155117: dataIn1 = 32'd283
; 
32'd155118: dataIn1 = 32'd454
; 
32'd155119: dataIn1 = 32'd2331
; 
32'd155120: dataIn1 = 32'd4005
; 
32'd155121: dataIn1 = 32'd5326
; 
32'd155122: dataIn1 = 32'd5327
; 
32'd155123: dataIn1 = 32'd5329
; 
32'd155124: dataIn1 = 32'd5460
; 
32'd155125: dataIn1 = 32'd109
; 
32'd155126: dataIn1 = 32'd455
; 
32'd155127: dataIn1 = 32'd2333
; 
32'd155128: dataIn1 = 32'd4017
; 
32'd155129: dataIn1 = 32'd5328
; 
32'd155130: dataIn1 = 32'd5329
; 
32'd155131: dataIn1 = 32'd5331
; 
32'd155132: dataIn1 = 32'd5461
; 
32'd155133: dataIn1 = 32'd109
; 
32'd155134: dataIn1 = 32'd454
; 
32'd155135: dataIn1 = 32'd2333
; 
32'd155136: dataIn1 = 32'd4014
; 
32'd155137: dataIn1 = 32'd5327
; 
32'd155138: dataIn1 = 32'd5328
; 
32'd155139: dataIn1 = 32'd5329
; 
32'd155140: dataIn1 = 32'd5460
; 
32'd155141: dataIn1 = 32'd291
; 
32'd155142: dataIn1 = 32'd456
; 
32'd155143: dataIn1 = 32'd2336
; 
32'd155144: dataIn1 = 32'd4033
; 
32'd155145: dataIn1 = 32'd5330
; 
32'd155146: dataIn1 = 32'd5331
; 
32'd155147: dataIn1 = 32'd5332
; 
32'd155148: dataIn1 = 32'd5462
; 
32'd155149: dataIn1 = 32'd291
; 
32'd155150: dataIn1 = 32'd455
; 
32'd155151: dataIn1 = 32'd2336
; 
32'd155152: dataIn1 = 32'd4031
; 
32'd155153: dataIn1 = 32'd5328
; 
32'd155154: dataIn1 = 32'd5330
; 
32'd155155: dataIn1 = 32'd5331
; 
32'd155156: dataIn1 = 32'd5461
; 
32'd155157: dataIn1 = 32'd158
; 
32'd155158: dataIn1 = 32'd456
; 
32'd155159: dataIn1 = 32'd2339
; 
32'd155160: dataIn1 = 32'd4041
; 
32'd155161: dataIn1 = 32'd5330
; 
32'd155162: dataIn1 = 32'd5332
; 
32'd155163: dataIn1 = 32'd5333
; 
32'd155164: dataIn1 = 32'd5462
; 
32'd155165: dataIn1 = 32'd158
; 
32'd155166: dataIn1 = 32'd457
; 
32'd155167: dataIn1 = 32'd2339
; 
32'd155168: dataIn1 = 32'd4038
; 
32'd155169: dataIn1 = 32'd5332
; 
32'd155170: dataIn1 = 32'd5333
; 
32'd155171: dataIn1 = 32'd5335
; 
32'd155172: dataIn1 = 32'd5463
; 
32'd155173: dataIn1 = 32'd290
; 
32'd155174: dataIn1 = 32'd458
; 
32'd155175: dataIn1 = 32'd2343
; 
32'd155176: dataIn1 = 32'd4054
; 
32'd155177: dataIn1 = 32'd5334
; 
32'd155178: dataIn1 = 32'd5335
; 
32'd155179: dataIn1 = 32'd5336
; 
32'd155180: dataIn1 = 32'd5464
; 
32'd155181: dataIn1 = 32'd290
; 
32'd155182: dataIn1 = 32'd457
; 
32'd155183: dataIn1 = 32'd2343
; 
32'd155184: dataIn1 = 32'd4053
; 
32'd155185: dataIn1 = 32'd5333
; 
32'd155186: dataIn1 = 32'd5334
; 
32'd155187: dataIn1 = 32'd5335
; 
32'd155188: dataIn1 = 32'd5463
; 
32'd155189: dataIn1 = 32'd110
; 
32'd155190: dataIn1 = 32'd458
; 
32'd155191: dataIn1 = 32'd2346
; 
32'd155192: dataIn1 = 32'd4063
; 
32'd155193: dataIn1 = 32'd5334
; 
32'd155194: dataIn1 = 32'd5336
; 
32'd155195: dataIn1 = 32'd5337
; 
32'd155196: dataIn1 = 32'd5464
; 
32'd155197: dataIn1 = 32'd110
; 
32'd155198: dataIn1 = 32'd459
; 
32'd155199: dataIn1 = 32'd2346
; 
32'd155200: dataIn1 = 32'd4061
; 
32'd155201: dataIn1 = 32'd5336
; 
32'd155202: dataIn1 = 32'd5337
; 
32'd155203: dataIn1 = 32'd5339
; 
32'd155204: dataIn1 = 32'd5465
; 
32'd155205: dataIn1 = 32'd300
; 
32'd155206: dataIn1 = 32'd460
; 
32'd155207: dataIn1 = 32'd2349
; 
32'd155208: dataIn1 = 32'd4080
; 
32'd155209: dataIn1 = 32'd5338
; 
32'd155210: dataIn1 = 32'd5339
; 
32'd155211: dataIn1 = 32'd5340
; 
32'd155212: dataIn1 = 32'd5466
; 
32'd155213: dataIn1 = 32'd300
; 
32'd155214: dataIn1 = 32'd459
; 
32'd155215: dataIn1 = 32'd2349
; 
32'd155216: dataIn1 = 32'd4077
; 
32'd155217: dataIn1 = 32'd5337
; 
32'd155218: dataIn1 = 32'd5338
; 
32'd155219: dataIn1 = 32'd5339
; 
32'd155220: dataIn1 = 32'd5465
; 
32'd155221: dataIn1 = 32'd160
; 
32'd155222: dataIn1 = 32'd460
; 
32'd155223: dataIn1 = 32'd2350
; 
32'd155224: dataIn1 = 32'd4090
; 
32'd155225: dataIn1 = 32'd5338
; 
32'd155226: dataIn1 = 32'd5340
; 
32'd155227: dataIn1 = 32'd5341
; 
32'd155228: dataIn1 = 32'd5466
; 
32'd155229: dataIn1 = 32'd160
; 
32'd155230: dataIn1 = 32'd461
; 
32'd155231: dataIn1 = 32'd2350
; 
32'd155232: dataIn1 = 32'd4088
; 
32'd155233: dataIn1 = 32'd5340
; 
32'd155234: dataIn1 = 32'd5341
; 
32'd155235: dataIn1 = 32'd5342
; 
32'd155236: dataIn1 = 32'd5467
; 
32'd155237: dataIn1 = 32'd299
; 
32'd155238: dataIn1 = 32'd461
; 
32'd155239: dataIn1 = 32'd2355
; 
32'd155240: dataIn1 = 32'd4103
; 
32'd155241: dataIn1 = 32'd5341
; 
32'd155242: dataIn1 = 32'd5342
; 
32'd155243: dataIn1 = 32'd5343
; 
32'd155244: dataIn1 = 32'd5467
; 
32'd155245: dataIn1 = 32'd299
; 
32'd155246: dataIn1 = 32'd462
; 
32'd155247: dataIn1 = 32'd2355
; 
32'd155248: dataIn1 = 32'd4101
; 
32'd155249: dataIn1 = 32'd5342
; 
32'd155250: dataIn1 = 32'd5343
; 
32'd155251: dataIn1 = 32'd5345
; 
32'd155252: dataIn1 = 32'd5468
; 
32'd155253: dataIn1 = 32'd111
; 
32'd155254: dataIn1 = 32'd463
; 
32'd155255: dataIn1 = 32'd2357
; 
32'd155256: dataIn1 = 32'd4113
; 
32'd155257: dataIn1 = 32'd5344
; 
32'd155258: dataIn1 = 32'd5345
; 
32'd155259: dataIn1 = 32'd5347
; 
32'd155260: dataIn1 = 32'd5469
; 
32'd155261: dataIn1 = 32'd111
; 
32'd155262: dataIn1 = 32'd462
; 
32'd155263: dataIn1 = 32'd2357
; 
32'd155264: dataIn1 = 32'd4110
; 
32'd155265: dataIn1 = 32'd5343
; 
32'd155266: dataIn1 = 32'd5344
; 
32'd155267: dataIn1 = 32'd5345
; 
32'd155268: dataIn1 = 32'd5468
; 
32'd155269: dataIn1 = 32'd307
; 
32'd155270: dataIn1 = 32'd464
; 
32'd155271: dataIn1 = 32'd2360
; 
32'd155272: dataIn1 = 32'd4129
; 
32'd155273: dataIn1 = 32'd5346
; 
32'd155274: dataIn1 = 32'd5347
; 
32'd155275: dataIn1 = 32'd5348
; 
32'd155276: dataIn1 = 32'd5470
; 
32'd155277: dataIn1 = 32'd307
; 
32'd155278: dataIn1 = 32'd463
; 
32'd155279: dataIn1 = 32'd2360
; 
32'd155280: dataIn1 = 32'd4127
; 
32'd155281: dataIn1 = 32'd5344
; 
32'd155282: dataIn1 = 32'd5346
; 
32'd155283: dataIn1 = 32'd5347
; 
32'd155284: dataIn1 = 32'd5469
; 
32'd155285: dataIn1 = 32'd164
; 
32'd155286: dataIn1 = 32'd464
; 
32'd155287: dataIn1 = 32'd2363
; 
32'd155288: dataIn1 = 32'd4137
; 
32'd155289: dataIn1 = 32'd5346
; 
32'd155290: dataIn1 = 32'd5348
; 
32'd155291: dataIn1 = 32'd5349
; 
32'd155292: dataIn1 = 32'd5470
; 
32'd155293: dataIn1 = 32'd164
; 
32'd155294: dataIn1 = 32'd465
; 
32'd155295: dataIn1 = 32'd2363
; 
32'd155296: dataIn1 = 32'd4134
; 
32'd155297: dataIn1 = 32'd5348
; 
32'd155298: dataIn1 = 32'd5349
; 
32'd155299: dataIn1 = 32'd5351
; 
32'd155300: dataIn1 = 32'd5471
; 
32'd155301: dataIn1 = 32'd306
; 
32'd155302: dataIn1 = 32'd466
; 
32'd155303: dataIn1 = 32'd2367
; 
32'd155304: dataIn1 = 32'd4150
; 
32'd155305: dataIn1 = 32'd5350
; 
32'd155306: dataIn1 = 32'd5351
; 
32'd155307: dataIn1 = 32'd5352
; 
32'd155308: dataIn1 = 32'd5472
; 
32'd155309: dataIn1 = 32'd306
; 
32'd155310: dataIn1 = 32'd465
; 
32'd155311: dataIn1 = 32'd2367
; 
32'd155312: dataIn1 = 32'd4149
; 
32'd155313: dataIn1 = 32'd5349
; 
32'd155314: dataIn1 = 32'd5350
; 
32'd155315: dataIn1 = 32'd5351
; 
32'd155316: dataIn1 = 32'd5471
; 
32'd155317: dataIn1 = 32'd112
; 
32'd155318: dataIn1 = 32'd466
; 
32'd155319: dataIn1 = 32'd2370
; 
32'd155320: dataIn1 = 32'd4159
; 
32'd155321: dataIn1 = 32'd5350
; 
32'd155322: dataIn1 = 32'd5352
; 
32'd155323: dataIn1 = 32'd5353
; 
32'd155324: dataIn1 = 32'd5472
; 
32'd155325: dataIn1 = 32'd112
; 
32'd155326: dataIn1 = 32'd467
; 
32'd155327: dataIn1 = 32'd2370
; 
32'd155328: dataIn1 = 32'd4157
; 
32'd155329: dataIn1 = 32'd5352
; 
32'd155330: dataIn1 = 32'd5353
; 
32'd155331: dataIn1 = 32'd5355
; 
32'd155332: dataIn1 = 32'd5473
; 
32'd155333: dataIn1 = 32'd316
; 
32'd155334: dataIn1 = 32'd468
; 
32'd155335: dataIn1 = 32'd2373
; 
32'd155336: dataIn1 = 32'd4176
; 
32'd155337: dataIn1 = 32'd5354
; 
32'd155338: dataIn1 = 32'd5355
; 
32'd155339: dataIn1 = 32'd5356
; 
32'd155340: dataIn1 = 32'd5474
; 
32'd155341: dataIn1 = 32'd316
; 
32'd155342: dataIn1 = 32'd467
; 
32'd155343: dataIn1 = 32'd2373
; 
32'd155344: dataIn1 = 32'd4173
; 
32'd155345: dataIn1 = 32'd5353
; 
32'd155346: dataIn1 = 32'd5354
; 
32'd155347: dataIn1 = 32'd5355
; 
32'd155348: dataIn1 = 32'd5473
; 
32'd155349: dataIn1 = 32'd166
; 
32'd155350: dataIn1 = 32'd468
; 
32'd155351: dataIn1 = 32'd2374
; 
32'd155352: dataIn1 = 32'd4186
; 
32'd155353: dataIn1 = 32'd5354
; 
32'd155354: dataIn1 = 32'd5356
; 
32'd155355: dataIn1 = 32'd5357
; 
32'd155356: dataIn1 = 32'd5474
; 
32'd155357: dataIn1 = 32'd166
; 
32'd155358: dataIn1 = 32'd469
; 
32'd155359: dataIn1 = 32'd2374
; 
32'd155360: dataIn1 = 32'd4184
; 
32'd155361: dataIn1 = 32'd5356
; 
32'd155362: dataIn1 = 32'd5357
; 
32'd155363: dataIn1 = 32'd5358
; 
32'd155364: dataIn1 = 32'd5475
; 
32'd155365: dataIn1 = 32'd315
; 
32'd155366: dataIn1 = 32'd469
; 
32'd155367: dataIn1 = 32'd2379
; 
32'd155368: dataIn1 = 32'd4199
; 
32'd155369: dataIn1 = 32'd5357
; 
32'd155370: dataIn1 = 32'd5358
; 
32'd155371: dataIn1 = 32'd5359
; 
32'd155372: dataIn1 = 32'd5475
; 
32'd155373: dataIn1 = 32'd315
; 
32'd155374: dataIn1 = 32'd470
; 
32'd155375: dataIn1 = 32'd2379
; 
32'd155376: dataIn1 = 32'd4197
; 
32'd155377: dataIn1 = 32'd5358
; 
32'd155378: dataIn1 = 32'd5359
; 
32'd155379: dataIn1 = 32'd5361
; 
32'd155380: dataIn1 = 32'd5476
; 
32'd155381: dataIn1 = 32'd113
; 
32'd155382: dataIn1 = 32'd471
; 
32'd155383: dataIn1 = 32'd2381
; 
32'd155384: dataIn1 = 32'd4209
; 
32'd155385: dataIn1 = 32'd5360
; 
32'd155386: dataIn1 = 32'd5361
; 
32'd155387: dataIn1 = 32'd5363
; 
32'd155388: dataIn1 = 32'd5477
; 
32'd155389: dataIn1 = 32'd113
; 
32'd155390: dataIn1 = 32'd470
; 
32'd155391: dataIn1 = 32'd2381
; 
32'd155392: dataIn1 = 32'd4206
; 
32'd155393: dataIn1 = 32'd5359
; 
32'd155394: dataIn1 = 32'd5360
; 
32'd155395: dataIn1 = 32'd5361
; 
32'd155396: dataIn1 = 32'd5476
; 
32'd155397: dataIn1 = 32'd323
; 
32'd155398: dataIn1 = 32'd472
; 
32'd155399: dataIn1 = 32'd2384
; 
32'd155400: dataIn1 = 32'd4225
; 
32'd155401: dataIn1 = 32'd5362
; 
32'd155402: dataIn1 = 32'd5363
; 
32'd155403: dataIn1 = 32'd5364
; 
32'd155404: dataIn1 = 32'd5478
; 
32'd155405: dataIn1 = 32'd323
; 
32'd155406: dataIn1 = 32'd471
; 
32'd155407: dataIn1 = 32'd2384
; 
32'd155408: dataIn1 = 32'd4223
; 
32'd155409: dataIn1 = 32'd5360
; 
32'd155410: dataIn1 = 32'd5362
; 
32'd155411: dataIn1 = 32'd5363
; 
32'd155412: dataIn1 = 32'd5477
; 
32'd155413: dataIn1 = 32'd170
; 
32'd155414: dataIn1 = 32'd472
; 
32'd155415: dataIn1 = 32'd2387
; 
32'd155416: dataIn1 = 32'd4233
; 
32'd155417: dataIn1 = 32'd5362
; 
32'd155418: dataIn1 = 32'd5364
; 
32'd155419: dataIn1 = 32'd5365
; 
32'd155420: dataIn1 = 32'd5478
; 
32'd155421: dataIn1 = 32'd170
; 
32'd155422: dataIn1 = 32'd473
; 
32'd155423: dataIn1 = 32'd2387
; 
32'd155424: dataIn1 = 32'd4230
; 
32'd155425: dataIn1 = 32'd5364
; 
32'd155426: dataIn1 = 32'd5365
; 
32'd155427: dataIn1 = 32'd5367
; 
32'd155428: dataIn1 = 32'd5479
; 
32'd155429: dataIn1 = 32'd322
; 
32'd155430: dataIn1 = 32'd474
; 
32'd155431: dataIn1 = 32'd2391
; 
32'd155432: dataIn1 = 32'd4246
; 
32'd155433: dataIn1 = 32'd5366
; 
32'd155434: dataIn1 = 32'd5367
; 
32'd155435: dataIn1 = 32'd5368
; 
32'd155436: dataIn1 = 32'd5480
; 
32'd155437: dataIn1 = 32'd322
; 
32'd155438: dataIn1 = 32'd473
; 
32'd155439: dataIn1 = 32'd2391
; 
32'd155440: dataIn1 = 32'd4245
; 
32'd155441: dataIn1 = 32'd5365
; 
32'd155442: dataIn1 = 32'd5366
; 
32'd155443: dataIn1 = 32'd5367
; 
32'd155444: dataIn1 = 32'd5479
; 
32'd155445: dataIn1 = 32'd114
; 
32'd155446: dataIn1 = 32'd474
; 
32'd155447: dataIn1 = 32'd2394
; 
32'd155448: dataIn1 = 32'd4255
; 
32'd155449: dataIn1 = 32'd5366
; 
32'd155450: dataIn1 = 32'd5368
; 
32'd155451: dataIn1 = 32'd5369
; 
32'd155452: dataIn1 = 32'd5480
; 
32'd155453: dataIn1 = 32'd114
; 
32'd155454: dataIn1 = 32'd475
; 
32'd155455: dataIn1 = 32'd2394
; 
32'd155456: dataIn1 = 32'd4253
; 
32'd155457: dataIn1 = 32'd5368
; 
32'd155458: dataIn1 = 32'd5369
; 
32'd155459: dataIn1 = 32'd5371
; 
32'd155460: dataIn1 = 32'd5481
; 
32'd155461: dataIn1 = 32'd332
; 
32'd155462: dataIn1 = 32'd476
; 
32'd155463: dataIn1 = 32'd2397
; 
32'd155464: dataIn1 = 32'd4272
; 
32'd155465: dataIn1 = 32'd5370
; 
32'd155466: dataIn1 = 32'd5371
; 
32'd155467: dataIn1 = 32'd5372
; 
32'd155468: dataIn1 = 32'd5482
; 
32'd155469: dataIn1 = 32'd332
; 
32'd155470: dataIn1 = 32'd475
; 
32'd155471: dataIn1 = 32'd2397
; 
32'd155472: dataIn1 = 32'd4269
; 
32'd155473: dataIn1 = 32'd5369
; 
32'd155474: dataIn1 = 32'd5370
; 
32'd155475: dataIn1 = 32'd5371
; 
32'd155476: dataIn1 = 32'd5481
; 
32'd155477: dataIn1 = 32'd172
; 
32'd155478: dataIn1 = 32'd476
; 
32'd155479: dataIn1 = 32'd2398
; 
32'd155480: dataIn1 = 32'd4282
; 
32'd155481: dataIn1 = 32'd5370
; 
32'd155482: dataIn1 = 32'd5372
; 
32'd155483: dataIn1 = 32'd5373
; 
32'd155484: dataIn1 = 32'd5482
; 
32'd155485: dataIn1 = 32'd172
; 
32'd155486: dataIn1 = 32'd477
; 
32'd155487: dataIn1 = 32'd2398
; 
32'd155488: dataIn1 = 32'd4280
; 
32'd155489: dataIn1 = 32'd5372
; 
32'd155490: dataIn1 = 32'd5373
; 
32'd155491: dataIn1 = 32'd5374
; 
32'd155492: dataIn1 = 32'd5483
; 
32'd155493: dataIn1 = 32'd331
; 
32'd155494: dataIn1 = 32'd477
; 
32'd155495: dataIn1 = 32'd2403
; 
32'd155496: dataIn1 = 32'd4295
; 
32'd155497: dataIn1 = 32'd5373
; 
32'd155498: dataIn1 = 32'd5374
; 
32'd155499: dataIn1 = 32'd5375
; 
32'd155500: dataIn1 = 32'd5483
; 
32'd155501: dataIn1 = 32'd331
; 
32'd155502: dataIn1 = 32'd478
; 
32'd155503: dataIn1 = 32'd2403
; 
32'd155504: dataIn1 = 32'd4293
; 
32'd155505: dataIn1 = 32'd5374
; 
32'd155506: dataIn1 = 32'd5375
; 
32'd155507: dataIn1 = 32'd5377
; 
32'd155508: dataIn1 = 32'd5484
; 
32'd155509: dataIn1 = 32'd115
; 
32'd155510: dataIn1 = 32'd479
; 
32'd155511: dataIn1 = 32'd2405
; 
32'd155512: dataIn1 = 32'd4305
; 
32'd155513: dataIn1 = 32'd5376
; 
32'd155514: dataIn1 = 32'd5377
; 
32'd155515: dataIn1 = 32'd5379
; 
32'd155516: dataIn1 = 32'd5485
; 
32'd155517: dataIn1 = 32'd115
; 
32'd155518: dataIn1 = 32'd478
; 
32'd155519: dataIn1 = 32'd2405
; 
32'd155520: dataIn1 = 32'd4302
; 
32'd155521: dataIn1 = 32'd5375
; 
32'd155522: dataIn1 = 32'd5376
; 
32'd155523: dataIn1 = 32'd5377
; 
32'd155524: dataIn1 = 32'd5484
; 
32'd155525: dataIn1 = 32'd339
; 
32'd155526: dataIn1 = 32'd480
; 
32'd155527: dataIn1 = 32'd2408
; 
32'd155528: dataIn1 = 32'd4321
; 
32'd155529: dataIn1 = 32'd5378
; 
32'd155530: dataIn1 = 32'd5379
; 
32'd155531: dataIn1 = 32'd5380
; 
32'd155532: dataIn1 = 32'd5486
; 
32'd155533: dataIn1 = 32'd339
; 
32'd155534: dataIn1 = 32'd479
; 
32'd155535: dataIn1 = 32'd2408
; 
32'd155536: dataIn1 = 32'd4319
; 
32'd155537: dataIn1 = 32'd5376
; 
32'd155538: dataIn1 = 32'd5378
; 
32'd155539: dataIn1 = 32'd5379
; 
32'd155540: dataIn1 = 32'd5485
; 
32'd155541: dataIn1 = 32'd176
; 
32'd155542: dataIn1 = 32'd480
; 
32'd155543: dataIn1 = 32'd2411
; 
32'd155544: dataIn1 = 32'd4329
; 
32'd155545: dataIn1 = 32'd5378
; 
32'd155546: dataIn1 = 32'd5380
; 
32'd155547: dataIn1 = 32'd5381
; 
32'd155548: dataIn1 = 32'd5486
; 
32'd155549: dataIn1 = 32'd176
; 
32'd155550: dataIn1 = 32'd481
; 
32'd155551: dataIn1 = 32'd2411
; 
32'd155552: dataIn1 = 32'd4326
; 
32'd155553: dataIn1 = 32'd5380
; 
32'd155554: dataIn1 = 32'd5381
; 
32'd155555: dataIn1 = 32'd5383
; 
32'd155556: dataIn1 = 32'd5487
; 
32'd155557: dataIn1 = 32'd338
; 
32'd155558: dataIn1 = 32'd482
; 
32'd155559: dataIn1 = 32'd2415
; 
32'd155560: dataIn1 = 32'd4342
; 
32'd155561: dataIn1 = 32'd5382
; 
32'd155562: dataIn1 = 32'd5383
; 
32'd155563: dataIn1 = 32'd5384
; 
32'd155564: dataIn1 = 32'd5488
; 
32'd155565: dataIn1 = 32'd338
; 
32'd155566: dataIn1 = 32'd481
; 
32'd155567: dataIn1 = 32'd2415
; 
32'd155568: dataIn1 = 32'd4341
; 
32'd155569: dataIn1 = 32'd5381
; 
32'd155570: dataIn1 = 32'd5382
; 
32'd155571: dataIn1 = 32'd5383
; 
32'd155572: dataIn1 = 32'd5487
; 
32'd155573: dataIn1 = 32'd116
; 
32'd155574: dataIn1 = 32'd482
; 
32'd155575: dataIn1 = 32'd2418
; 
32'd155576: dataIn1 = 32'd4351
; 
32'd155577: dataIn1 = 32'd5382
; 
32'd155578: dataIn1 = 32'd5384
; 
32'd155579: dataIn1 = 32'd5385
; 
32'd155580: dataIn1 = 32'd5488
; 
32'd155581: dataIn1 = 32'd116
; 
32'd155582: dataIn1 = 32'd483
; 
32'd155583: dataIn1 = 32'd2418
; 
32'd155584: dataIn1 = 32'd4349
; 
32'd155585: dataIn1 = 32'd5384
; 
32'd155586: dataIn1 = 32'd5385
; 
32'd155587: dataIn1 = 32'd5387
; 
32'd155588: dataIn1 = 32'd5489
; 
32'd155589: dataIn1 = 32'd348
; 
32'd155590: dataIn1 = 32'd484
; 
32'd155591: dataIn1 = 32'd2421
; 
32'd155592: dataIn1 = 32'd4368
; 
32'd155593: dataIn1 = 32'd5386
; 
32'd155594: dataIn1 = 32'd5387
; 
32'd155595: dataIn1 = 32'd5388
; 
32'd155596: dataIn1 = 32'd5490
; 
32'd155597: dataIn1 = 32'd348
; 
32'd155598: dataIn1 = 32'd483
; 
32'd155599: dataIn1 = 32'd2421
; 
32'd155600: dataIn1 = 32'd4365
; 
32'd155601: dataIn1 = 32'd5385
; 
32'd155602: dataIn1 = 32'd5386
; 
32'd155603: dataIn1 = 32'd5387
; 
32'd155604: dataIn1 = 32'd5489
; 
32'd155605: dataIn1 = 32'd178
; 
32'd155606: dataIn1 = 32'd484
; 
32'd155607: dataIn1 = 32'd2422
; 
32'd155608: dataIn1 = 32'd4378
; 
32'd155609: dataIn1 = 32'd5386
; 
32'd155610: dataIn1 = 32'd5388
; 
32'd155611: dataIn1 = 32'd5389
; 
32'd155612: dataIn1 = 32'd5490
; 
32'd155613: dataIn1 = 32'd178
; 
32'd155614: dataIn1 = 32'd485
; 
32'd155615: dataIn1 = 32'd2422
; 
32'd155616: dataIn1 = 32'd4376
; 
32'd155617: dataIn1 = 32'd5388
; 
32'd155618: dataIn1 = 32'd5389
; 
32'd155619: dataIn1 = 32'd5390
; 
32'd155620: dataIn1 = 32'd5491
; 
32'd155621: dataIn1 = 32'd347
; 
32'd155622: dataIn1 = 32'd485
; 
32'd155623: dataIn1 = 32'd2427
; 
32'd155624: dataIn1 = 32'd4391
; 
32'd155625: dataIn1 = 32'd5389
; 
32'd155626: dataIn1 = 32'd5390
; 
32'd155627: dataIn1 = 32'd5391
; 
32'd155628: dataIn1 = 32'd5491
; 
32'd155629: dataIn1 = 32'd347
; 
32'd155630: dataIn1 = 32'd486
; 
32'd155631: dataIn1 = 32'd2427
; 
32'd155632: dataIn1 = 32'd4389
; 
32'd155633: dataIn1 = 32'd5390
; 
32'd155634: dataIn1 = 32'd5391
; 
32'd155635: dataIn1 = 32'd5393
; 
32'd155636: dataIn1 = 32'd5492
; 
32'd155637: dataIn1 = 32'd117
; 
32'd155638: dataIn1 = 32'd487
; 
32'd155639: dataIn1 = 32'd2429
; 
32'd155640: dataIn1 = 32'd4401
; 
32'd155641: dataIn1 = 32'd5392
; 
32'd155642: dataIn1 = 32'd5393
; 
32'd155643: dataIn1 = 32'd5395
; 
32'd155644: dataIn1 = 32'd5493
; 
32'd155645: dataIn1 = 32'd117
; 
32'd155646: dataIn1 = 32'd486
; 
32'd155647: dataIn1 = 32'd2429
; 
32'd155648: dataIn1 = 32'd4398
; 
32'd155649: dataIn1 = 32'd5391
; 
32'd155650: dataIn1 = 32'd5392
; 
32'd155651: dataIn1 = 32'd5393
; 
32'd155652: dataIn1 = 32'd5492
; 
32'd155653: dataIn1 = 32'd355
; 
32'd155654: dataIn1 = 32'd488
; 
32'd155655: dataIn1 = 32'd2432
; 
32'd155656: dataIn1 = 32'd4417
; 
32'd155657: dataIn1 = 32'd5394
; 
32'd155658: dataIn1 = 32'd5395
; 
32'd155659: dataIn1 = 32'd5396
; 
32'd155660: dataIn1 = 32'd5494
; 
32'd155661: dataIn1 = 32'd355
; 
32'd155662: dataIn1 = 32'd487
; 
32'd155663: dataIn1 = 32'd2432
; 
32'd155664: dataIn1 = 32'd4415
; 
32'd155665: dataIn1 = 32'd5392
; 
32'd155666: dataIn1 = 32'd5394
; 
32'd155667: dataIn1 = 32'd5395
; 
32'd155668: dataIn1 = 32'd5493
; 
32'd155669: dataIn1 = 32'd182
; 
32'd155670: dataIn1 = 32'd488
; 
32'd155671: dataIn1 = 32'd2435
; 
32'd155672: dataIn1 = 32'd4425
; 
32'd155673: dataIn1 = 32'd5394
; 
32'd155674: dataIn1 = 32'd5396
; 
32'd155675: dataIn1 = 32'd5397
; 
32'd155676: dataIn1 = 32'd5494
; 
32'd155677: dataIn1 = 32'd182
; 
32'd155678: dataIn1 = 32'd489
; 
32'd155679: dataIn1 = 32'd2435
; 
32'd155680: dataIn1 = 32'd4422
; 
32'd155681: dataIn1 = 32'd5396
; 
32'd155682: dataIn1 = 32'd5397
; 
32'd155683: dataIn1 = 32'd5399
; 
32'd155684: dataIn1 = 32'd5495
; 
32'd155685: dataIn1 = 32'd354
; 
32'd155686: dataIn1 = 32'd490
; 
32'd155687: dataIn1 = 32'd2439
; 
32'd155688: dataIn1 = 32'd4438
; 
32'd155689: dataIn1 = 32'd5398
; 
32'd155690: dataIn1 = 32'd5399
; 
32'd155691: dataIn1 = 32'd5400
; 
32'd155692: dataIn1 = 32'd5496
; 
32'd155693: dataIn1 = 32'd354
; 
32'd155694: dataIn1 = 32'd489
; 
32'd155695: dataIn1 = 32'd2439
; 
32'd155696: dataIn1 = 32'd4437
; 
32'd155697: dataIn1 = 32'd5397
; 
32'd155698: dataIn1 = 32'd5398
; 
32'd155699: dataIn1 = 32'd5399
; 
32'd155700: dataIn1 = 32'd5495
; 
32'd155701: dataIn1 = 32'd118
; 
32'd155702: dataIn1 = 32'd490
; 
32'd155703: dataIn1 = 32'd2442
; 
32'd155704: dataIn1 = 32'd4447
; 
32'd155705: dataIn1 = 32'd5398
; 
32'd155706: dataIn1 = 32'd5400
; 
32'd155707: dataIn1 = 32'd5401
; 
32'd155708: dataIn1 = 32'd5496
; 
32'd155709: dataIn1 = 32'd118
; 
32'd155710: dataIn1 = 32'd491
; 
32'd155711: dataIn1 = 32'd2442
; 
32'd155712: dataIn1 = 32'd4445
; 
32'd155713: dataIn1 = 32'd5400
; 
32'd155714: dataIn1 = 32'd5401
; 
32'd155715: dataIn1 = 32'd5403
; 
32'd155716: dataIn1 = 32'd5497
; 
32'd155717: dataIn1 = 32'd364
; 
32'd155718: dataIn1 = 32'd492
; 
32'd155719: dataIn1 = 32'd2445
; 
32'd155720: dataIn1 = 32'd4464
; 
32'd155721: dataIn1 = 32'd5402
; 
32'd155722: dataIn1 = 32'd5403
; 
32'd155723: dataIn1 = 32'd5404
; 
32'd155724: dataIn1 = 32'd5498
; 
32'd155725: dataIn1 = 32'd364
; 
32'd155726: dataIn1 = 32'd491
; 
32'd155727: dataIn1 = 32'd2445
; 
32'd155728: dataIn1 = 32'd4461
; 
32'd155729: dataIn1 = 32'd5401
; 
32'd155730: dataIn1 = 32'd5402
; 
32'd155731: dataIn1 = 32'd5403
; 
32'd155732: dataIn1 = 32'd5497
; 
32'd155733: dataIn1 = 32'd184
; 
32'd155734: dataIn1 = 32'd492
; 
32'd155735: dataIn1 = 32'd2446
; 
32'd155736: dataIn1 = 32'd4474
; 
32'd155737: dataIn1 = 32'd5402
; 
32'd155738: dataIn1 = 32'd5404
; 
32'd155739: dataIn1 = 32'd5405
; 
32'd155740: dataIn1 = 32'd5498
; 
32'd155741: dataIn1 = 32'd184
; 
32'd155742: dataIn1 = 32'd493
; 
32'd155743: dataIn1 = 32'd2446
; 
32'd155744: dataIn1 = 32'd4472
; 
32'd155745: dataIn1 = 32'd5404
; 
32'd155746: dataIn1 = 32'd5405
; 
32'd155747: dataIn1 = 32'd5406
; 
32'd155748: dataIn1 = 32'd5499
; 
32'd155749: dataIn1 = 32'd363
; 
32'd155750: dataIn1 = 32'd493
; 
32'd155751: dataIn1 = 32'd2451
; 
32'd155752: dataIn1 = 32'd4487
; 
32'd155753: dataIn1 = 32'd5405
; 
32'd155754: dataIn1 = 32'd5406
; 
32'd155755: dataIn1 = 32'd5407
; 
32'd155756: dataIn1 = 32'd5499
; 
32'd155757: dataIn1 = 32'd363
; 
32'd155758: dataIn1 = 32'd494
; 
32'd155759: dataIn1 = 32'd2451
; 
32'd155760: dataIn1 = 32'd4485
; 
32'd155761: dataIn1 = 32'd5406
; 
32'd155762: dataIn1 = 32'd5407
; 
32'd155763: dataIn1 = 32'd5409
; 
32'd155764: dataIn1 = 32'd5500
; 
32'd155765: dataIn1 = 32'd119
; 
32'd155766: dataIn1 = 32'd495
; 
32'd155767: dataIn1 = 32'd2453
; 
32'd155768: dataIn1 = 32'd4497
; 
32'd155769: dataIn1 = 32'd5408
; 
32'd155770: dataIn1 = 32'd5409
; 
32'd155771: dataIn1 = 32'd5411
; 
32'd155772: dataIn1 = 32'd5501
; 
32'd155773: dataIn1 = 32'd119
; 
32'd155774: dataIn1 = 32'd494
; 
32'd155775: dataIn1 = 32'd2453
; 
32'd155776: dataIn1 = 32'd4494
; 
32'd155777: dataIn1 = 32'd5407
; 
32'd155778: dataIn1 = 32'd5408
; 
32'd155779: dataIn1 = 32'd5409
; 
32'd155780: dataIn1 = 32'd5500
; 
32'd155781: dataIn1 = 32'd371
; 
32'd155782: dataIn1 = 32'd496
; 
32'd155783: dataIn1 = 32'd2456
; 
32'd155784: dataIn1 = 32'd4513
; 
32'd155785: dataIn1 = 32'd5410
; 
32'd155786: dataIn1 = 32'd5411
; 
32'd155787: dataIn1 = 32'd5412
; 
32'd155788: dataIn1 = 32'd5502
; 
32'd155789: dataIn1 = 32'd371
; 
32'd155790: dataIn1 = 32'd495
; 
32'd155791: dataIn1 = 32'd2456
; 
32'd155792: dataIn1 = 32'd4511
; 
32'd155793: dataIn1 = 32'd5408
; 
32'd155794: dataIn1 = 32'd5410
; 
32'd155795: dataIn1 = 32'd5411
; 
32'd155796: dataIn1 = 32'd5501
; 
32'd155797: dataIn1 = 32'd188
; 
32'd155798: dataIn1 = 32'd496
; 
32'd155799: dataIn1 = 32'd2459
; 
32'd155800: dataIn1 = 32'd4521
; 
32'd155801: dataIn1 = 32'd5410
; 
32'd155802: dataIn1 = 32'd5412
; 
32'd155803: dataIn1 = 32'd5413
; 
32'd155804: dataIn1 = 32'd5502
; 
32'd155805: dataIn1 = 32'd188
; 
32'd155806: dataIn1 = 32'd497
; 
32'd155807: dataIn1 = 32'd2459
; 
32'd155808: dataIn1 = 32'd4518
; 
32'd155809: dataIn1 = 32'd5412
; 
32'd155810: dataIn1 = 32'd5413
; 
32'd155811: dataIn1 = 32'd5415
; 
32'd155812: dataIn1 = 32'd5503
; 
32'd155813: dataIn1 = 32'd370
; 
32'd155814: dataIn1 = 32'd498
; 
32'd155815: dataIn1 = 32'd2463
; 
32'd155816: dataIn1 = 32'd4534
; 
32'd155817: dataIn1 = 32'd5414
; 
32'd155818: dataIn1 = 32'd5415
; 
32'd155819: dataIn1 = 32'd5416
; 
32'd155820: dataIn1 = 32'd5504
; 
32'd155821: dataIn1 = 32'd370
; 
32'd155822: dataIn1 = 32'd497
; 
32'd155823: dataIn1 = 32'd2463
; 
32'd155824: dataIn1 = 32'd4533
; 
32'd155825: dataIn1 = 32'd5413
; 
32'd155826: dataIn1 = 32'd5414
; 
32'd155827: dataIn1 = 32'd5415
; 
32'd155828: dataIn1 = 32'd5503
; 
32'd155829: dataIn1 = 32'd120
; 
32'd155830: dataIn1 = 32'd498
; 
32'd155831: dataIn1 = 32'd2466
; 
32'd155832: dataIn1 = 32'd4541
; 
32'd155833: dataIn1 = 32'd4543
; 
32'd155834: dataIn1 = 32'd5414
; 
32'd155835: dataIn1 = 32'd5416
; 
32'd155836: dataIn1 = 32'd5417
; 
32'd155837: dataIn1 = 32'd5504
; 
32'd155838: dataIn1 = 32'd120
; 
32'd155839: dataIn1 = 32'd499
; 
32'd155840: dataIn1 = 32'd4541
; 
32'd155841: dataIn1 = 32'd4557
; 
32'd155842: dataIn1 = 32'd5416
; 
32'd155843: dataIn1 = 32'd5417
; 
32'd155844: dataIn1 = 32'd5419
; 
32'd155845: dataIn1 = 32'd5505
; 
32'd155846: dataIn1 = 32'd380
; 
32'd155847: dataIn1 = 32'd500
; 
32'd155848: dataIn1 = 32'd4560
; 
32'd155849: dataIn1 = 32'd4570
; 
32'd155850: dataIn1 = 32'd5418
; 
32'd155851: dataIn1 = 32'd5419
; 
32'd155852: dataIn1 = 32'd5420
; 
32'd155853: dataIn1 = 32'd5506
; 
32'd155854: dataIn1 = 32'd380
; 
32'd155855: dataIn1 = 32'd2469
; 
32'd155856: dataIn1 = 32'd4557
; 
32'd155857: dataIn1 = 32'd4560
; 
32'd155858: dataIn1 = 32'd5417
; 
32'd155859: dataIn1 = 32'd5418
; 
32'd155860: dataIn1 = 32'd5419
; 
32'd155861: dataIn1 = 32'd5505
; 
32'd155862: dataIn1 = 32'd190
; 
32'd155863: dataIn1 = 32'd2470
; 
32'd155864: dataIn1 = 32'd4568
; 
32'd155865: dataIn1 = 32'd4570
; 
32'd155866: dataIn1 = 32'd5418
; 
32'd155867: dataIn1 = 32'd5420
; 
32'd155868: dataIn1 = 32'd5421
; 
32'd155869: dataIn1 = 32'd5506
; 
32'd155870: dataIn1 = 32'd190
; 
32'd155871: dataIn1 = 32'd501
; 
32'd155872: dataIn1 = 32'd4568
; 
32'd155873: dataIn1 = 32'd4583
; 
32'd155874: dataIn1 = 32'd5420
; 
32'd155875: dataIn1 = 32'd5421
; 
32'd155876: dataIn1 = 32'd5422
; 
32'd155877: dataIn1 = 32'd5507
; 
32'd155878: dataIn1 = 32'd379
; 
32'd155879: dataIn1 = 32'd2475
; 
32'd155880: dataIn1 = 32'd4581
; 
32'd155881: dataIn1 = 32'd4583
; 
32'd155882: dataIn1 = 32'd5421
; 
32'd155883: dataIn1 = 32'd5422
; 
32'd155884: dataIn1 = 32'd5423
; 
32'd155885: dataIn1 = 32'd5507
; 
32'd155886: dataIn1 = 32'd379
; 
32'd155887: dataIn1 = 32'd502
; 
32'd155888: dataIn1 = 32'd4581
; 
32'd155889: dataIn1 = 32'd4590
; 
32'd155890: dataIn1 = 32'd5422
; 
32'd155891: dataIn1 = 32'd5423
; 
32'd155892: dataIn1 = 32'd5425
; 
32'd155893: dataIn1 = 32'd5508
; 
32'd155894: dataIn1 = 32'd121
; 
32'd155895: dataIn1 = 32'd503
; 
32'd155896: dataIn1 = 32'd4593
; 
32'd155897: dataIn1 = 32'd5424
; 
32'd155898: dataIn1 = 32'd5425
; 
32'd155899: dataIn1 = 32'd121
; 
32'd155900: dataIn1 = 32'd2477
; 
32'd155901: dataIn1 = 32'd4590
; 
32'd155902: dataIn1 = 32'd4593
; 
32'd155903: dataIn1 = 32'd5423
; 
32'd155904: dataIn1 = 32'd5424
; 
32'd155905: dataIn1 = 32'd5425
; 
32'd155906: dataIn1 = 32'd5508
; 
32'd155907: dataIn1 = 32'd205
; 
32'd155908: dataIn1 = 32'd395
; 
32'd155909: dataIn1 = 32'd751
; 
32'd155910: dataIn1 = 32'd3890
; 
32'd155911: dataIn1 = 32'd4602
; 
32'd155912: dataIn1 = 32'd5426
; 
32'd155913: dataIn1 = 32'd5509
; 
32'd155914: dataIn1 = 32'd128
; 
32'd155915: dataIn1 = 32'd398
; 
32'd155916: dataIn1 = 32'd774
; 
32'd155917: dataIn1 = 32'd3891
; 
32'd155918: dataIn1 = 32'd4603
; 
32'd155919: dataIn1 = 32'd5427
; 
32'd155920: dataIn1 = 32'd5510
; 
32'd155921: dataIn1 = 32'd212
; 
32'd155922: dataIn1 = 32'd980
; 
32'd155923: dataIn1 = 32'd2049
; 
32'd155924: dataIn1 = 32'd2544
; 
32'd155925: dataIn1 = 32'd5307
; 
32'd155926: dataIn1 = 32'd5428
; 
32'd155927: dataIn1 = 32'd5429
; 
32'd155928: dataIn1 = 32'd5511
; 
32'd155929: dataIn1 = 32'd212
; 
32'd155930: dataIn1 = 32'd1042
; 
32'd155931: dataIn1 = 32'd2544
; 
32'd155932: dataIn1 = 32'd4627
; 
32'd155933: dataIn1 = 32'd5428
; 
32'd155934: dataIn1 = 32'd5429
; 
32'd155935: dataIn1 = 32'd10267
; 
32'd155936: dataIn1 = 32'd10275
; 
32'd155937: dataIn1 = 32'd2554
; 
32'd155938: dataIn1 = 32'd2619
; 
32'd155939: dataIn1 = 32'd4821
; 
32'd155940: dataIn1 = 32'd4838
; 
32'd155941: dataIn1 = 32'd5318
; 
32'd155942: dataIn1 = 32'd5430
; 
32'd155943: dataIn1 = 32'd5512
; 
32'd155944: dataIn1 = 32'd14
; 
32'd155945: dataIn1 = 32'd5431
; 
32'd155946: dataIn1 = 32'd6706
; 
32'd155947: dataIn1 = 32'd6707
; 
32'd155948: dataIn1 = 32'd6730
; 
32'd155949: dataIn1 = 32'd6734
; 
32'd155950: dataIn1 = 32'd9312
; 
32'd155951: dataIn1 = 32'd14
; 
32'd155952: dataIn1 = 32'd5432
; 
32'd155953: dataIn1 = 32'd5513
; 
32'd155954: dataIn1 = 32'd6704
; 
32'd155955: dataIn1 = 32'd6705
; 
32'd155956: dataIn1 = 32'd6733
; 
32'd155957: dataIn1 = 32'd6734
; 
32'd155958: dataIn1 = 32'd17
; 
32'd155959: dataIn1 = 32'd5433
; 
32'd155960: dataIn1 = 32'd5515
; 
32'd155961: dataIn1 = 32'd9289
; 
32'd155962: dataIn1 = 32'd9290
; 
32'd155963: dataIn1 = 32'd9328
; 
32'd155964: dataIn1 = 32'd9339
; 
32'd155965: dataIn1 = 32'd17
; 
32'd155966: dataIn1 = 32'd5434
; 
32'd155967: dataIn1 = 32'd5514
; 
32'd155968: dataIn1 = 32'd9287
; 
32'd155969: dataIn1 = 32'd9288
; 
32'd155970: dataIn1 = 32'd9327
; 
32'd155971: dataIn1 = 32'd9328
; 
32'd155972: dataIn1 = 32'd18
; 
32'd155973: dataIn1 = 32'd5435
; 
32'd155974: dataIn1 = 32'd5517
; 
32'd155975: dataIn1 = 32'd9295
; 
32'd155976: dataIn1 = 32'd9296
; 
32'd155977: dataIn1 = 32'd9330
; 
32'd155978: dataIn1 = 32'd9331
; 
32'd155979: dataIn1 = 32'd18
; 
32'd155980: dataIn1 = 32'd5436
; 
32'd155981: dataIn1 = 32'd5516
; 
32'd155982: dataIn1 = 32'd9293
; 
32'd155983: dataIn1 = 32'd9294
; 
32'd155984: dataIn1 = 32'd9324
; 
32'd155985: dataIn1 = 32'd9330
; 
32'd155986: dataIn1 = 32'd19
; 
32'd155987: dataIn1 = 32'd5437
; 
32'd155988: dataIn1 = 32'd5519
; 
32'd155989: dataIn1 = 32'd6710
; 
32'd155990: dataIn1 = 32'd6711
; 
32'd155991: dataIn1 = 32'd6736
; 
32'd155992: dataIn1 = 32'd6737
; 
32'd155993: dataIn1 = 32'd19
; 
32'd155994: dataIn1 = 32'd5438
; 
32'd155995: dataIn1 = 32'd5518
; 
32'd155996: dataIn1 = 32'd6708
; 
32'd155997: dataIn1 = 32'd6709
; 
32'd155998: dataIn1 = 32'd6735
; 
32'd155999: dataIn1 = 32'd6736
; 
32'd156000: dataIn1 = 32'd5439
; 
32'd156001: dataIn1 = 32'd5521
; 
32'd156002: dataIn1 = 32'd6715
; 
32'd156003: dataIn1 = 32'd6716
; 
32'd156004: dataIn1 = 32'd6739
; 
32'd156005: dataIn1 = 32'd6740
; 
32'd156006: dataIn1 = 32'd9755
; 
32'd156007: dataIn1 = 32'd5440
; 
32'd156008: dataIn1 = 32'd6739
; 
32'd156009: dataIn1 = 32'd9752
; 
32'd156010: dataIn1 = 32'd10127
; 
32'd156011: dataIn1 = 32'd10131
; 
32'd156012: dataIn1 = 32'd10147
; 
32'd156013: dataIn1 = 32'd10148
; 
32'd156014: dataIn1 = 32'd21
; 
32'd156015: dataIn1 = 32'd5441
; 
32'd156016: dataIn1 = 32'd5523
; 
32'd156017: dataIn1 = 32'd9301
; 
32'd156018: dataIn1 = 32'd9302
; 
32'd156019: dataIn1 = 32'd9326
; 
32'd156020: dataIn1 = 32'd9333
; 
32'd156021: dataIn1 = 32'd21
; 
32'd156022: dataIn1 = 32'd5442
; 
32'd156023: dataIn1 = 32'd5522
; 
32'd156024: dataIn1 = 32'd9299
; 
32'd156025: dataIn1 = 32'd9300
; 
32'd156026: dataIn1 = 32'd9332
; 
32'd156027: dataIn1 = 32'd9333
; 
32'd156028: dataIn1 = 32'd22
; 
32'd156029: dataIn1 = 32'd5443
; 
32'd156030: dataIn1 = 32'd5524
; 
32'd156031: dataIn1 = 32'd9307
; 
32'd156032: dataIn1 = 32'd9308
; 
32'd156033: dataIn1 = 32'd9335
; 
32'd156034: dataIn1 = 32'd9336
; 
32'd156035: dataIn1 = 32'd22
; 
32'd156036: dataIn1 = 32'd5444
; 
32'd156037: dataIn1 = 32'd6731
; 
32'd156038: dataIn1 = 32'd9305
; 
32'd156039: dataIn1 = 32'd9306
; 
32'd156040: dataIn1 = 32'd9318
; 
32'd156041: dataIn1 = 32'd9335
; 
32'd156042: dataIn1 = 32'd1138
; 
32'd156043: dataIn1 = 32'd5445
; 
32'd156044: dataIn1 = 32'd5514
; 
32'd156045: dataIn1 = 32'd9291
; 
32'd156046: dataIn1 = 32'd9292
; 
32'd156047: dataIn1 = 32'd9327
; 
32'd156048: dataIn1 = 32'd9329
; 
32'd156049: dataIn1 = 32'd1138
; 
32'd156050: dataIn1 = 32'd5446
; 
32'd156051: dataIn1 = 32'd5517
; 
32'd156052: dataIn1 = 32'd9297
; 
32'd156053: dataIn1 = 32'd9298
; 
32'd156054: dataIn1 = 32'd9329
; 
32'd156055: dataIn1 = 32'd9331
; 
32'd156056: dataIn1 = 32'd1139
; 
32'd156057: dataIn1 = 32'd5447
; 
32'd156058: dataIn1 = 32'd5516
; 
32'd156059: dataIn1 = 32'd9281
; 
32'd156060: dataIn1 = 32'd9282
; 
32'd156061: dataIn1 = 32'd9323
; 
32'd156062: dataIn1 = 32'd9324
; 
32'd156063: dataIn1 = 32'd1139
; 
32'd156064: dataIn1 = 32'd5448
; 
32'd156065: dataIn1 = 32'd5519
; 
32'd156066: dataIn1 = 32'd6721
; 
32'd156067: dataIn1 = 32'd6722
; 
32'd156068: dataIn1 = 32'd6737
; 
32'd156069: dataIn1 = 32'd9323
; 
32'd156070: dataIn1 = 32'd1140
; 
32'd156071: dataIn1 = 32'd5449
; 
32'd156072: dataIn1 = 32'd5518
; 
32'd156073: dataIn1 = 32'd6726
; 
32'd156074: dataIn1 = 32'd6727
; 
32'd156075: dataIn1 = 32'd6735
; 
32'd156076: dataIn1 = 32'd6743
; 
32'd156077: dataIn1 = 32'd1140
; 
32'd156078: dataIn1 = 32'd5450
; 
32'd156079: dataIn1 = 32'd5521
; 
32'd156080: dataIn1 = 32'd6723
; 
32'd156081: dataIn1 = 32'd6724
; 
32'd156082: dataIn1 = 32'd6740
; 
32'd156083: dataIn1 = 32'd6743
; 
32'd156084: dataIn1 = 32'd5451
; 
32'd156085: dataIn1 = 32'd6728
; 
32'd156086: dataIn1 = 32'd6729
; 
32'd156087: dataIn1 = 32'd6738
; 
32'd156088: dataIn1 = 32'd9325
; 
32'd156089: dataIn1 = 32'd9672
; 
32'd156090: dataIn1 = 32'd10224
; 
32'd156091: dataIn1 = 32'd10277
; 
32'd156092: dataIn1 = 32'd5452
; 
32'd156093: dataIn1 = 32'd5523
; 
32'd156094: dataIn1 = 32'd9283
; 
32'd156095: dataIn1 = 32'd9284
; 
32'd156096: dataIn1 = 32'd9325
; 
32'd156097: dataIn1 = 32'd9326
; 
32'd156098: dataIn1 = 32'd10281
; 
32'd156099: dataIn1 = 32'd1142
; 
32'd156100: dataIn1 = 32'd5453
; 
32'd156101: dataIn1 = 32'd5522
; 
32'd156102: dataIn1 = 32'd9303
; 
32'd156103: dataIn1 = 32'd9304
; 
32'd156104: dataIn1 = 32'd9332
; 
32'd156105: dataIn1 = 32'd9334
; 
32'd156106: dataIn1 = 32'd1142
; 
32'd156107: dataIn1 = 32'd5454
; 
32'd156108: dataIn1 = 32'd5524
; 
32'd156109: dataIn1 = 32'd9309
; 
32'd156110: dataIn1 = 32'd9310
; 
32'd156111: dataIn1 = 32'd9334
; 
32'd156112: dataIn1 = 32'd9336
; 
32'd156113: dataIn1 = 32'd65
; 
32'd156114: dataIn1 = 32'd75
; 
32'd156115: dataIn1 = 32'd2213
; 
32'd156116: dataIn1 = 32'd5312
; 
32'd156117: dataIn1 = 32'd5455
; 
32'd156118: dataIn1 = 32'd98
; 
32'd156119: dataIn1 = 32'd99
; 
32'd156120: dataIn1 = 32'd5314
; 
32'd156121: dataIn1 = 32'd5317
; 
32'd156122: dataIn1 = 32'd5456
; 
32'd156123: dataIn1 = 32'd152
; 
32'd156124: dataIn1 = 32'd276
; 
32'd156125: dataIn1 = 32'd566
; 
32'd156126: dataIn1 = 32'd3502
; 
32'd156127: dataIn1 = 32'd5319
; 
32'd156128: dataIn1 = 32'd5457
; 
32'd156129: dataIn1 = 32'd5525
; 
32'd156130: dataIn1 = 32'd153
; 
32'd156131: dataIn1 = 32'd284
; 
32'd156132: dataIn1 = 32'd5321
; 
32'd156133: dataIn1 = 32'd5324
; 
32'd156134: dataIn1 = 32'd5458
; 
32'd156135: dataIn1 = 32'd5531
; 
32'd156136: dataIn1 = 32'd5532
; 
32'd156137: dataIn1 = 32'd153
; 
32'd156138: dataIn1 = 32'd283
; 
32'd156139: dataIn1 = 32'd5325
; 
32'd156140: dataIn1 = 32'd5326
; 
32'd156141: dataIn1 = 32'd5459
; 
32'd156142: dataIn1 = 32'd5533
; 
32'd156143: dataIn1 = 32'd5534
; 
32'd156144: dataIn1 = 32'd109
; 
32'd156145: dataIn1 = 32'd283
; 
32'd156146: dataIn1 = 32'd5327
; 
32'd156147: dataIn1 = 32'd5329
; 
32'd156148: dataIn1 = 32'd5460
; 
32'd156149: dataIn1 = 32'd5535
; 
32'd156150: dataIn1 = 32'd5536
; 
32'd156151: dataIn1 = 32'd109
; 
32'd156152: dataIn1 = 32'd291
; 
32'd156153: dataIn1 = 32'd5328
; 
32'd156154: dataIn1 = 32'd5331
; 
32'd156155: dataIn1 = 32'd5461
; 
32'd156156: dataIn1 = 32'd5537
; 
32'd156157: dataIn1 = 32'd5538
; 
32'd156158: dataIn1 = 32'd158
; 
32'd156159: dataIn1 = 32'd291
; 
32'd156160: dataIn1 = 32'd5330
; 
32'd156161: dataIn1 = 32'd5332
; 
32'd156162: dataIn1 = 32'd5462
; 
32'd156163: dataIn1 = 32'd5539
; 
32'd156164: dataIn1 = 32'd5540
; 
32'd156165: dataIn1 = 32'd158
; 
32'd156166: dataIn1 = 32'd290
; 
32'd156167: dataIn1 = 32'd5333
; 
32'd156168: dataIn1 = 32'd5335
; 
32'd156169: dataIn1 = 32'd5463
; 
32'd156170: dataIn1 = 32'd5541
; 
32'd156171: dataIn1 = 32'd5542
; 
32'd156172: dataIn1 = 32'd110
; 
32'd156173: dataIn1 = 32'd290
; 
32'd156174: dataIn1 = 32'd5334
; 
32'd156175: dataIn1 = 32'd5336
; 
32'd156176: dataIn1 = 32'd5464
; 
32'd156177: dataIn1 = 32'd5543
; 
32'd156178: dataIn1 = 32'd5544
; 
32'd156179: dataIn1 = 32'd110
; 
32'd156180: dataIn1 = 32'd300
; 
32'd156181: dataIn1 = 32'd5337
; 
32'd156182: dataIn1 = 32'd5339
; 
32'd156183: dataIn1 = 32'd5465
; 
32'd156184: dataIn1 = 32'd5545
; 
32'd156185: dataIn1 = 32'd5546
; 
32'd156186: dataIn1 = 32'd160
; 
32'd156187: dataIn1 = 32'd300
; 
32'd156188: dataIn1 = 32'd5338
; 
32'd156189: dataIn1 = 32'd5340
; 
32'd156190: dataIn1 = 32'd5466
; 
32'd156191: dataIn1 = 32'd5547
; 
32'd156192: dataIn1 = 32'd5548
; 
32'd156193: dataIn1 = 32'd160
; 
32'd156194: dataIn1 = 32'd299
; 
32'd156195: dataIn1 = 32'd5341
; 
32'd156196: dataIn1 = 32'd5342
; 
32'd156197: dataIn1 = 32'd5467
; 
32'd156198: dataIn1 = 32'd5549
; 
32'd156199: dataIn1 = 32'd5550
; 
32'd156200: dataIn1 = 32'd111
; 
32'd156201: dataIn1 = 32'd299
; 
32'd156202: dataIn1 = 32'd5343
; 
32'd156203: dataIn1 = 32'd5345
; 
32'd156204: dataIn1 = 32'd5468
; 
32'd156205: dataIn1 = 32'd5551
; 
32'd156206: dataIn1 = 32'd5552
; 
32'd156207: dataIn1 = 32'd111
; 
32'd156208: dataIn1 = 32'd307
; 
32'd156209: dataIn1 = 32'd5344
; 
32'd156210: dataIn1 = 32'd5347
; 
32'd156211: dataIn1 = 32'd5469
; 
32'd156212: dataIn1 = 32'd5553
; 
32'd156213: dataIn1 = 32'd5554
; 
32'd156214: dataIn1 = 32'd164
; 
32'd156215: dataIn1 = 32'd307
; 
32'd156216: dataIn1 = 32'd5346
; 
32'd156217: dataIn1 = 32'd5348
; 
32'd156218: dataIn1 = 32'd5470
; 
32'd156219: dataIn1 = 32'd5555
; 
32'd156220: dataIn1 = 32'd5556
; 
32'd156221: dataIn1 = 32'd164
; 
32'd156222: dataIn1 = 32'd306
; 
32'd156223: dataIn1 = 32'd5349
; 
32'd156224: dataIn1 = 32'd5351
; 
32'd156225: dataIn1 = 32'd5471
; 
32'd156226: dataIn1 = 32'd5557
; 
32'd156227: dataIn1 = 32'd5558
; 
32'd156228: dataIn1 = 32'd112
; 
32'd156229: dataIn1 = 32'd306
; 
32'd156230: dataIn1 = 32'd5350
; 
32'd156231: dataIn1 = 32'd5352
; 
32'd156232: dataIn1 = 32'd5472
; 
32'd156233: dataIn1 = 32'd5559
; 
32'd156234: dataIn1 = 32'd5560
; 
32'd156235: dataIn1 = 32'd112
; 
32'd156236: dataIn1 = 32'd316
; 
32'd156237: dataIn1 = 32'd5353
; 
32'd156238: dataIn1 = 32'd5355
; 
32'd156239: dataIn1 = 32'd5473
; 
32'd156240: dataIn1 = 32'd5561
; 
32'd156241: dataIn1 = 32'd5562
; 
32'd156242: dataIn1 = 32'd166
; 
32'd156243: dataIn1 = 32'd316
; 
32'd156244: dataIn1 = 32'd5354
; 
32'd156245: dataIn1 = 32'd5356
; 
32'd156246: dataIn1 = 32'd5474
; 
32'd156247: dataIn1 = 32'd5563
; 
32'd156248: dataIn1 = 32'd5564
; 
32'd156249: dataIn1 = 32'd166
; 
32'd156250: dataIn1 = 32'd315
; 
32'd156251: dataIn1 = 32'd5357
; 
32'd156252: dataIn1 = 32'd5358
; 
32'd156253: dataIn1 = 32'd5475
; 
32'd156254: dataIn1 = 32'd5565
; 
32'd156255: dataIn1 = 32'd5566
; 
32'd156256: dataIn1 = 32'd113
; 
32'd156257: dataIn1 = 32'd315
; 
32'd156258: dataIn1 = 32'd5359
; 
32'd156259: dataIn1 = 32'd5361
; 
32'd156260: dataIn1 = 32'd5476
; 
32'd156261: dataIn1 = 32'd5567
; 
32'd156262: dataIn1 = 32'd5568
; 
32'd156263: dataIn1 = 32'd113
; 
32'd156264: dataIn1 = 32'd323
; 
32'd156265: dataIn1 = 32'd5360
; 
32'd156266: dataIn1 = 32'd5363
; 
32'd156267: dataIn1 = 32'd5477
; 
32'd156268: dataIn1 = 32'd5569
; 
32'd156269: dataIn1 = 32'd5570
; 
32'd156270: dataIn1 = 32'd170
; 
32'd156271: dataIn1 = 32'd323
; 
32'd156272: dataIn1 = 32'd5362
; 
32'd156273: dataIn1 = 32'd5364
; 
32'd156274: dataIn1 = 32'd5478
; 
32'd156275: dataIn1 = 32'd5571
; 
32'd156276: dataIn1 = 32'd5572
; 
32'd156277: dataIn1 = 32'd170
; 
32'd156278: dataIn1 = 32'd322
; 
32'd156279: dataIn1 = 32'd5365
; 
32'd156280: dataIn1 = 32'd5367
; 
32'd156281: dataIn1 = 32'd5479
; 
32'd156282: dataIn1 = 32'd5573
; 
32'd156283: dataIn1 = 32'd5574
; 
32'd156284: dataIn1 = 32'd114
; 
32'd156285: dataIn1 = 32'd322
; 
32'd156286: dataIn1 = 32'd5366
; 
32'd156287: dataIn1 = 32'd5368
; 
32'd156288: dataIn1 = 32'd5480
; 
32'd156289: dataIn1 = 32'd5575
; 
32'd156290: dataIn1 = 32'd5576
; 
32'd156291: dataIn1 = 32'd114
; 
32'd156292: dataIn1 = 32'd332
; 
32'd156293: dataIn1 = 32'd5369
; 
32'd156294: dataIn1 = 32'd5371
; 
32'd156295: dataIn1 = 32'd5481
; 
32'd156296: dataIn1 = 32'd5577
; 
32'd156297: dataIn1 = 32'd5578
; 
32'd156298: dataIn1 = 32'd172
; 
32'd156299: dataIn1 = 32'd332
; 
32'd156300: dataIn1 = 32'd5370
; 
32'd156301: dataIn1 = 32'd5372
; 
32'd156302: dataIn1 = 32'd5482
; 
32'd156303: dataIn1 = 32'd5579
; 
32'd156304: dataIn1 = 32'd5580
; 
32'd156305: dataIn1 = 32'd172
; 
32'd156306: dataIn1 = 32'd331
; 
32'd156307: dataIn1 = 32'd5373
; 
32'd156308: dataIn1 = 32'd5374
; 
32'd156309: dataIn1 = 32'd5483
; 
32'd156310: dataIn1 = 32'd5581
; 
32'd156311: dataIn1 = 32'd5582
; 
32'd156312: dataIn1 = 32'd115
; 
32'd156313: dataIn1 = 32'd331
; 
32'd156314: dataIn1 = 32'd5375
; 
32'd156315: dataIn1 = 32'd5377
; 
32'd156316: dataIn1 = 32'd5484
; 
32'd156317: dataIn1 = 32'd5583
; 
32'd156318: dataIn1 = 32'd5584
; 
32'd156319: dataIn1 = 32'd115
; 
32'd156320: dataIn1 = 32'd339
; 
32'd156321: dataIn1 = 32'd5376
; 
32'd156322: dataIn1 = 32'd5379
; 
32'd156323: dataIn1 = 32'd5485
; 
32'd156324: dataIn1 = 32'd5585
; 
32'd156325: dataIn1 = 32'd5586
; 
32'd156326: dataIn1 = 32'd176
; 
32'd156327: dataIn1 = 32'd339
; 
32'd156328: dataIn1 = 32'd5378
; 
32'd156329: dataIn1 = 32'd5380
; 
32'd156330: dataIn1 = 32'd5486
; 
32'd156331: dataIn1 = 32'd5587
; 
32'd156332: dataIn1 = 32'd5588
; 
32'd156333: dataIn1 = 32'd176
; 
32'd156334: dataIn1 = 32'd338
; 
32'd156335: dataIn1 = 32'd5381
; 
32'd156336: dataIn1 = 32'd5383
; 
32'd156337: dataIn1 = 32'd5487
; 
32'd156338: dataIn1 = 32'd5589
; 
32'd156339: dataIn1 = 32'd5590
; 
32'd156340: dataIn1 = 32'd116
; 
32'd156341: dataIn1 = 32'd338
; 
32'd156342: dataIn1 = 32'd5382
; 
32'd156343: dataIn1 = 32'd5384
; 
32'd156344: dataIn1 = 32'd5488
; 
32'd156345: dataIn1 = 32'd5591
; 
32'd156346: dataIn1 = 32'd5592
; 
32'd156347: dataIn1 = 32'd116
; 
32'd156348: dataIn1 = 32'd348
; 
32'd156349: dataIn1 = 32'd5385
; 
32'd156350: dataIn1 = 32'd5387
; 
32'd156351: dataIn1 = 32'd5489
; 
32'd156352: dataIn1 = 32'd5593
; 
32'd156353: dataIn1 = 32'd5594
; 
32'd156354: dataIn1 = 32'd178
; 
32'd156355: dataIn1 = 32'd348
; 
32'd156356: dataIn1 = 32'd5386
; 
32'd156357: dataIn1 = 32'd5388
; 
32'd156358: dataIn1 = 32'd5490
; 
32'd156359: dataIn1 = 32'd5595
; 
32'd156360: dataIn1 = 32'd5596
; 
32'd156361: dataIn1 = 32'd178
; 
32'd156362: dataIn1 = 32'd347
; 
32'd156363: dataIn1 = 32'd5389
; 
32'd156364: dataIn1 = 32'd5390
; 
32'd156365: dataIn1 = 32'd5491
; 
32'd156366: dataIn1 = 32'd5597
; 
32'd156367: dataIn1 = 32'd5598
; 
32'd156368: dataIn1 = 32'd117
; 
32'd156369: dataIn1 = 32'd347
; 
32'd156370: dataIn1 = 32'd5391
; 
32'd156371: dataIn1 = 32'd5393
; 
32'd156372: dataIn1 = 32'd5492
; 
32'd156373: dataIn1 = 32'd5599
; 
32'd156374: dataIn1 = 32'd5600
; 
32'd156375: dataIn1 = 32'd117
; 
32'd156376: dataIn1 = 32'd355
; 
32'd156377: dataIn1 = 32'd5392
; 
32'd156378: dataIn1 = 32'd5395
; 
32'd156379: dataIn1 = 32'd5493
; 
32'd156380: dataIn1 = 32'd5601
; 
32'd156381: dataIn1 = 32'd5602
; 
32'd156382: dataIn1 = 32'd182
; 
32'd156383: dataIn1 = 32'd355
; 
32'd156384: dataIn1 = 32'd5394
; 
32'd156385: dataIn1 = 32'd5396
; 
32'd156386: dataIn1 = 32'd5494
; 
32'd156387: dataIn1 = 32'd5603
; 
32'd156388: dataIn1 = 32'd5604
; 
32'd156389: dataIn1 = 32'd182
; 
32'd156390: dataIn1 = 32'd354
; 
32'd156391: dataIn1 = 32'd5397
; 
32'd156392: dataIn1 = 32'd5399
; 
32'd156393: dataIn1 = 32'd5495
; 
32'd156394: dataIn1 = 32'd5605
; 
32'd156395: dataIn1 = 32'd5606
; 
32'd156396: dataIn1 = 32'd118
; 
32'd156397: dataIn1 = 32'd354
; 
32'd156398: dataIn1 = 32'd5398
; 
32'd156399: dataIn1 = 32'd5400
; 
32'd156400: dataIn1 = 32'd5496
; 
32'd156401: dataIn1 = 32'd5607
; 
32'd156402: dataIn1 = 32'd5608
; 
32'd156403: dataIn1 = 32'd118
; 
32'd156404: dataIn1 = 32'd364
; 
32'd156405: dataIn1 = 32'd5401
; 
32'd156406: dataIn1 = 32'd5403
; 
32'd156407: dataIn1 = 32'd5497
; 
32'd156408: dataIn1 = 32'd5609
; 
32'd156409: dataIn1 = 32'd5610
; 
32'd156410: dataIn1 = 32'd184
; 
32'd156411: dataIn1 = 32'd364
; 
32'd156412: dataIn1 = 32'd5402
; 
32'd156413: dataIn1 = 32'd5404
; 
32'd156414: dataIn1 = 32'd5498
; 
32'd156415: dataIn1 = 32'd5611
; 
32'd156416: dataIn1 = 32'd5612
; 
32'd156417: dataIn1 = 32'd184
; 
32'd156418: dataIn1 = 32'd363
; 
32'd156419: dataIn1 = 32'd5405
; 
32'd156420: dataIn1 = 32'd5406
; 
32'd156421: dataIn1 = 32'd5499
; 
32'd156422: dataIn1 = 32'd5613
; 
32'd156423: dataIn1 = 32'd5614
; 
32'd156424: dataIn1 = 32'd119
; 
32'd156425: dataIn1 = 32'd363
; 
32'd156426: dataIn1 = 32'd5407
; 
32'd156427: dataIn1 = 32'd5409
; 
32'd156428: dataIn1 = 32'd5500
; 
32'd156429: dataIn1 = 32'd5615
; 
32'd156430: dataIn1 = 32'd5616
; 
32'd156431: dataIn1 = 32'd119
; 
32'd156432: dataIn1 = 32'd371
; 
32'd156433: dataIn1 = 32'd5408
; 
32'd156434: dataIn1 = 32'd5411
; 
32'd156435: dataIn1 = 32'd5501
; 
32'd156436: dataIn1 = 32'd5617
; 
32'd156437: dataIn1 = 32'd5618
; 
32'd156438: dataIn1 = 32'd188
; 
32'd156439: dataIn1 = 32'd371
; 
32'd156440: dataIn1 = 32'd5410
; 
32'd156441: dataIn1 = 32'd5412
; 
32'd156442: dataIn1 = 32'd5502
; 
32'd156443: dataIn1 = 32'd5619
; 
32'd156444: dataIn1 = 32'd5620
; 
32'd156445: dataIn1 = 32'd188
; 
32'd156446: dataIn1 = 32'd370
; 
32'd156447: dataIn1 = 32'd5413
; 
32'd156448: dataIn1 = 32'd5415
; 
32'd156449: dataIn1 = 32'd5503
; 
32'd156450: dataIn1 = 32'd5621
; 
32'd156451: dataIn1 = 32'd5622
; 
32'd156452: dataIn1 = 32'd120
; 
32'd156453: dataIn1 = 32'd370
; 
32'd156454: dataIn1 = 32'd5414
; 
32'd156455: dataIn1 = 32'd5416
; 
32'd156456: dataIn1 = 32'd5504
; 
32'd156457: dataIn1 = 32'd5623
; 
32'd156458: dataIn1 = 32'd5624
; 
32'd156459: dataIn1 = 32'd120
; 
32'd156460: dataIn1 = 32'd380
; 
32'd156461: dataIn1 = 32'd5417
; 
32'd156462: dataIn1 = 32'd5419
; 
32'd156463: dataIn1 = 32'd5505
; 
32'd156464: dataIn1 = 32'd5625
; 
32'd156465: dataIn1 = 32'd5626
; 
32'd156466: dataIn1 = 32'd190
; 
32'd156467: dataIn1 = 32'd380
; 
32'd156468: dataIn1 = 32'd5418
; 
32'd156469: dataIn1 = 32'd5420
; 
32'd156470: dataIn1 = 32'd5506
; 
32'd156471: dataIn1 = 32'd5627
; 
32'd156472: dataIn1 = 32'd5628
; 
32'd156473: dataIn1 = 32'd190
; 
32'd156474: dataIn1 = 32'd379
; 
32'd156475: dataIn1 = 32'd5421
; 
32'd156476: dataIn1 = 32'd5422
; 
32'd156477: dataIn1 = 32'd5507
; 
32'd156478: dataIn1 = 32'd5629
; 
32'd156479: dataIn1 = 32'd5630
; 
32'd156480: dataIn1 = 32'd121
; 
32'd156481: dataIn1 = 32'd379
; 
32'd156482: dataIn1 = 32'd5423
; 
32'd156483: dataIn1 = 32'd5425
; 
32'd156484: dataIn1 = 32'd5508
; 
32'd156485: dataIn1 = 32'd5631
; 
32'd156486: dataIn1 = 32'd5632
; 
32'd156487: dataIn1 = 32'd395
; 
32'd156488: dataIn1 = 32'd399
; 
32'd156489: dataIn1 = 32'd760
; 
32'd156490: dataIn1 = 32'd3890
; 
32'd156491: dataIn1 = 32'd5426
; 
32'd156492: dataIn1 = 32'd5509
; 
32'd156493: dataIn1 = 32'd5510
; 
32'd156494: dataIn1 = 32'd398
; 
32'd156495: dataIn1 = 32'd399
; 
32'd156496: dataIn1 = 32'd760
; 
32'd156497: dataIn1 = 32'd3891
; 
32'd156498: dataIn1 = 32'd5427
; 
32'd156499: dataIn1 = 32'd5509
; 
32'd156500: dataIn1 = 32'd5510
; 
32'd156501: dataIn1 = 32'd212
; 
32'd156502: dataIn1 = 32'd979
; 
32'd156503: dataIn1 = 32'd1043
; 
32'd156504: dataIn1 = 32'd2049
; 
32'd156505: dataIn1 = 32'd5428
; 
32'd156506: dataIn1 = 32'd5511
; 
32'd156507: dataIn1 = 32'd1073
; 
32'd156508: dataIn1 = 32'd2553
; 
32'd156509: dataIn1 = 32'd2554
; 
32'd156510: dataIn1 = 32'd4821
; 
32'd156511: dataIn1 = 32'd5430
; 
32'd156512: dataIn1 = 32'd5512
; 
32'd156513: dataIn1 = 32'd14
; 
32'd156514: dataIn1 = 32'd1135
; 
32'd156515: dataIn1 = 32'd2735
; 
32'd156516: dataIn1 = 32'd3434
; 
32'd156517: dataIn1 = 32'd5432
; 
32'd156518: dataIn1 = 32'd5513
; 
32'd156519: dataIn1 = 32'd6733
; 
32'd156520: dataIn1 = 32'd17
; 
32'd156521: dataIn1 = 32'd1138
; 
32'd156522: dataIn1 = 32'd2748
; 
32'd156523: dataIn1 = 32'd5434
; 
32'd156524: dataIn1 = 32'd5445
; 
32'd156525: dataIn1 = 32'd5514
; 
32'd156526: dataIn1 = 32'd9327
; 
32'd156527: dataIn1 = 32'd17
; 
32'd156528: dataIn1 = 32'd1137
; 
32'd156529: dataIn1 = 32'd2745
; 
32'd156530: dataIn1 = 32'd3419
; 
32'd156531: dataIn1 = 32'd5433
; 
32'd156532: dataIn1 = 32'd5515
; 
32'd156533: dataIn1 = 32'd9339
; 
32'd156534: dataIn1 = 32'd18
; 
32'd156535: dataIn1 = 32'd1139
; 
32'd156536: dataIn1 = 32'd2107
; 
32'd156537: dataIn1 = 32'd5436
; 
32'd156538: dataIn1 = 32'd5447
; 
32'd156539: dataIn1 = 32'd5516
; 
32'd156540: dataIn1 = 32'd9324
; 
32'd156541: dataIn1 = 32'd18
; 
32'd156542: dataIn1 = 32'd1138
; 
32'd156543: dataIn1 = 32'd2108
; 
32'd156544: dataIn1 = 32'd5435
; 
32'd156545: dataIn1 = 32'd5446
; 
32'd156546: dataIn1 = 32'd5517
; 
32'd156547: dataIn1 = 32'd9331
; 
32'd156548: dataIn1 = 32'd19
; 
32'd156549: dataIn1 = 32'd1140
; 
32'd156550: dataIn1 = 32'd2111
; 
32'd156551: dataIn1 = 32'd5438
; 
32'd156552: dataIn1 = 32'd5449
; 
32'd156553: dataIn1 = 32'd5518
; 
32'd156554: dataIn1 = 32'd6735
; 
32'd156555: dataIn1 = 32'd19
; 
32'd156556: dataIn1 = 32'd1139
; 
32'd156557: dataIn1 = 32'd2109
; 
32'd156558: dataIn1 = 32'd5437
; 
32'd156559: dataIn1 = 32'd5448
; 
32'd156560: dataIn1 = 32'd5519
; 
32'd156561: dataIn1 = 32'd6737
; 
32'd156562: dataIn1 = 32'd5520
; 
32'd156563: dataIn1 = 32'd9672
; 
32'd156564: dataIn1 = 32'd9822
; 
32'd156565: dataIn1 = 32'd9823
; 
32'd156566: dataIn1 = 32'd10132
; 
32'd156567: dataIn1 = 32'd10133
; 
32'd156568: dataIn1 = 32'd10276
; 
32'd156569: dataIn1 = 32'd20
; 
32'd156570: dataIn1 = 32'd1140
; 
32'd156571: dataIn1 = 32'd5439
; 
32'd156572: dataIn1 = 32'd5450
; 
32'd156573: dataIn1 = 32'd5521
; 
32'd156574: dataIn1 = 32'd6740
; 
32'd156575: dataIn1 = 32'd9452
; 
32'd156576: dataIn1 = 32'd9676
; 
32'd156577: dataIn1 = 32'd9755
; 
32'd156578: dataIn1 = 32'd21
; 
32'd156579: dataIn1 = 32'd1142
; 
32'd156580: dataIn1 = 32'd2117
; 
32'd156581: dataIn1 = 32'd5442
; 
32'd156582: dataIn1 = 32'd5453
; 
32'd156583: dataIn1 = 32'd5522
; 
32'd156584: dataIn1 = 32'd9332
; 
32'd156585: dataIn1 = 32'd21
; 
32'd156586: dataIn1 = 32'd1141
; 
32'd156587: dataIn1 = 32'd5441
; 
32'd156588: dataIn1 = 32'd5452
; 
32'd156589: dataIn1 = 32'd5523
; 
32'd156590: dataIn1 = 32'd9326
; 
32'd156591: dataIn1 = 32'd10154
; 
32'd156592: dataIn1 = 32'd10225
; 
32'd156593: dataIn1 = 32'd10281
; 
32'd156594: dataIn1 = 32'd22
; 
32'd156595: dataIn1 = 32'd1142
; 
32'd156596: dataIn1 = 32'd2118
; 
32'd156597: dataIn1 = 32'd5443
; 
32'd156598: dataIn1 = 32'd5454
; 
32'd156599: dataIn1 = 32'd5524
; 
32'd156600: dataIn1 = 32'd9336
; 
32'd156601: dataIn1 = 32'd275
; 
32'd156602: dataIn1 = 32'd276
; 
32'd156603: dataIn1 = 32'd566
; 
32'd156604: dataIn1 = 32'd567
; 
32'd156605: dataIn1 = 32'd5457
; 
32'd156606: dataIn1 = 32'd5525
; 
32'd156607: dataIn1 = 32'd5526
; 
32'd156608: dataIn1 = 32'd274
; 
32'd156609: dataIn1 = 32'd276
; 
32'd156610: dataIn1 = 32'd567
; 
32'd156611: dataIn1 = 32'd1720
; 
32'd156612: dataIn1 = 32'd5525
; 
32'd156613: dataIn1 = 32'd5526
; 
32'd156614: dataIn1 = 32'd5527
; 
32'd156615: dataIn1 = 32'd108
; 
32'd156616: dataIn1 = 32'd276
; 
32'd156617: dataIn1 = 32'd1720
; 
32'd156618: dataIn1 = 32'd5320
; 
32'd156619: dataIn1 = 32'd5526
; 
32'd156620: dataIn1 = 32'd5527
; 
32'd156621: dataIn1 = 32'd5528
; 
32'd156622: dataIn1 = 32'd108
; 
32'd156623: dataIn1 = 32'd448
; 
32'd156624: dataIn1 = 32'd5320
; 
32'd156625: dataIn1 = 32'd5322
; 
32'd156626: dataIn1 = 32'd5527
; 
32'd156627: dataIn1 = 32'd5528
; 
32'd156628: dataIn1 = 32'd5529
; 
32'd156629: dataIn1 = 32'd108
; 
32'd156630: dataIn1 = 32'd284
; 
32'd156631: dataIn1 = 32'd1722
; 
32'd156632: dataIn1 = 32'd5322
; 
32'd156633: dataIn1 = 32'd5528
; 
32'd156634: dataIn1 = 32'd5529
; 
32'd156635: dataIn1 = 32'd5530
; 
32'd156636: dataIn1 = 32'd278
; 
32'd156637: dataIn1 = 32'd284
; 
32'd156638: dataIn1 = 32'd582
; 
32'd156639: dataIn1 = 32'd1722
; 
32'd156640: dataIn1 = 32'd5529
; 
32'd156641: dataIn1 = 32'd5530
; 
32'd156642: dataIn1 = 32'd5531
; 
32'd156643: dataIn1 = 32'd281
; 
32'd156644: dataIn1 = 32'd284
; 
32'd156645: dataIn1 = 32'd582
; 
32'd156646: dataIn1 = 32'd5458
; 
32'd156647: dataIn1 = 32'd5530
; 
32'd156648: dataIn1 = 32'd5531
; 
32'd156649: dataIn1 = 32'd5532
; 
32'd156650: dataIn1 = 32'd153
; 
32'd156651: dataIn1 = 32'd281
; 
32'd156652: dataIn1 = 32'd575
; 
32'd156653: dataIn1 = 32'd5458
; 
32'd156654: dataIn1 = 32'd5531
; 
32'd156655: dataIn1 = 32'd5532
; 
32'd156656: dataIn1 = 32'd5533
; 
32'd156657: dataIn1 = 32'd153
; 
32'd156658: dataIn1 = 32'd280
; 
32'd156659: dataIn1 = 32'd575
; 
32'd156660: dataIn1 = 32'd5459
; 
32'd156661: dataIn1 = 32'd5532
; 
32'd156662: dataIn1 = 32'd5533
; 
32'd156663: dataIn1 = 32'd5534
; 
32'd156664: dataIn1 = 32'd280
; 
32'd156665: dataIn1 = 32'd283
; 
32'd156666: dataIn1 = 32'd581
; 
32'd156667: dataIn1 = 32'd5459
; 
32'd156668: dataIn1 = 32'd5533
; 
32'd156669: dataIn1 = 32'd5534
; 
32'd156670: dataIn1 = 32'd5535
; 
32'd156671: dataIn1 = 32'd282
; 
32'd156672: dataIn1 = 32'd283
; 
32'd156673: dataIn1 = 32'd581
; 
32'd156674: dataIn1 = 32'd5460
; 
32'd156675: dataIn1 = 32'd5534
; 
32'd156676: dataIn1 = 32'd5535
; 
32'd156677: dataIn1 = 32'd5536
; 
32'd156678: dataIn1 = 32'd109
; 
32'd156679: dataIn1 = 32'd282
; 
32'd156680: dataIn1 = 32'd598
; 
32'd156681: dataIn1 = 32'd5460
; 
32'd156682: dataIn1 = 32'd5535
; 
32'd156683: dataIn1 = 32'd5536
; 
32'd156684: dataIn1 = 32'd5537
; 
32'd156685: dataIn1 = 32'd109
; 
32'd156686: dataIn1 = 32'd292
; 
32'd156687: dataIn1 = 32'd598
; 
32'd156688: dataIn1 = 32'd5461
; 
32'd156689: dataIn1 = 32'd5536
; 
32'd156690: dataIn1 = 32'd5537
; 
32'd156691: dataIn1 = 32'd5538
; 
32'd156692: dataIn1 = 32'd291
; 
32'd156693: dataIn1 = 32'd292
; 
32'd156694: dataIn1 = 32'd594
; 
32'd156695: dataIn1 = 32'd5461
; 
32'd156696: dataIn1 = 32'd5537
; 
32'd156697: dataIn1 = 32'd5538
; 
32'd156698: dataIn1 = 32'd5539
; 
32'd156699: dataIn1 = 32'd288
; 
32'd156700: dataIn1 = 32'd291
; 
32'd156701: dataIn1 = 32'd594
; 
32'd156702: dataIn1 = 32'd5462
; 
32'd156703: dataIn1 = 32'd5538
; 
32'd156704: dataIn1 = 32'd5539
; 
32'd156705: dataIn1 = 32'd5540
; 
32'd156706: dataIn1 = 32'd158
; 
32'd156707: dataIn1 = 32'd288
; 
32'd156708: dataIn1 = 32'd588
; 
32'd156709: dataIn1 = 32'd5462
; 
32'd156710: dataIn1 = 32'd5539
; 
32'd156711: dataIn1 = 32'd5540
; 
32'd156712: dataIn1 = 32'd5541
; 
32'd156713: dataIn1 = 32'd158
; 
32'd156714: dataIn1 = 32'd287
; 
32'd156715: dataIn1 = 32'd588
; 
32'd156716: dataIn1 = 32'd5463
; 
32'd156717: dataIn1 = 32'd5540
; 
32'd156718: dataIn1 = 32'd5541
; 
32'd156719: dataIn1 = 32'd5542
; 
32'd156720: dataIn1 = 32'd287
; 
32'd156721: dataIn1 = 32'd290
; 
32'd156722: dataIn1 = 32'd593
; 
32'd156723: dataIn1 = 32'd5463
; 
32'd156724: dataIn1 = 32'd5541
; 
32'd156725: dataIn1 = 32'd5542
; 
32'd156726: dataIn1 = 32'd5543
; 
32'd156727: dataIn1 = 32'd289
; 
32'd156728: dataIn1 = 32'd290
; 
32'd156729: dataIn1 = 32'd593
; 
32'd156730: dataIn1 = 32'd5464
; 
32'd156731: dataIn1 = 32'd5542
; 
32'd156732: dataIn1 = 32'd5543
; 
32'd156733: dataIn1 = 32'd5544
; 
32'd156734: dataIn1 = 32'd110
; 
32'd156735: dataIn1 = 32'd289
; 
32'd156736: dataIn1 = 32'd599
; 
32'd156737: dataIn1 = 32'd5464
; 
32'd156738: dataIn1 = 32'd5543
; 
32'd156739: dataIn1 = 32'd5544
; 
32'd156740: dataIn1 = 32'd5545
; 
32'd156741: dataIn1 = 32'd110
; 
32'd156742: dataIn1 = 32'd294
; 
32'd156743: dataIn1 = 32'd599
; 
32'd156744: dataIn1 = 32'd5465
; 
32'd156745: dataIn1 = 32'd5544
; 
32'd156746: dataIn1 = 32'd5545
; 
32'd156747: dataIn1 = 32'd5546
; 
32'd156748: dataIn1 = 32'd294
; 
32'd156749: dataIn1 = 32'd300
; 
32'd156750: dataIn1 = 32'd610
; 
32'd156751: dataIn1 = 32'd5465
; 
32'd156752: dataIn1 = 32'd5545
; 
32'd156753: dataIn1 = 32'd5546
; 
32'd156754: dataIn1 = 32'd5547
; 
32'd156755: dataIn1 = 32'd297
; 
32'd156756: dataIn1 = 32'd300
; 
32'd156757: dataIn1 = 32'd610
; 
32'd156758: dataIn1 = 32'd5466
; 
32'd156759: dataIn1 = 32'd5546
; 
32'd156760: dataIn1 = 32'd5547
; 
32'd156761: dataIn1 = 32'd5548
; 
32'd156762: dataIn1 = 32'd160
; 
32'd156763: dataIn1 = 32'd297
; 
32'd156764: dataIn1 = 32'd603
; 
32'd156765: dataIn1 = 32'd5466
; 
32'd156766: dataIn1 = 32'd5547
; 
32'd156767: dataIn1 = 32'd5548
; 
32'd156768: dataIn1 = 32'd5549
; 
32'd156769: dataIn1 = 32'd160
; 
32'd156770: dataIn1 = 32'd296
; 
32'd156771: dataIn1 = 32'd603
; 
32'd156772: dataIn1 = 32'd5467
; 
32'd156773: dataIn1 = 32'd5548
; 
32'd156774: dataIn1 = 32'd5549
; 
32'd156775: dataIn1 = 32'd5550
; 
32'd156776: dataIn1 = 32'd296
; 
32'd156777: dataIn1 = 32'd299
; 
32'd156778: dataIn1 = 32'd609
; 
32'd156779: dataIn1 = 32'd5467
; 
32'd156780: dataIn1 = 32'd5549
; 
32'd156781: dataIn1 = 32'd5550
; 
32'd156782: dataIn1 = 32'd5551
; 
32'd156783: dataIn1 = 32'd298
; 
32'd156784: dataIn1 = 32'd299
; 
32'd156785: dataIn1 = 32'd609
; 
32'd156786: dataIn1 = 32'd5468
; 
32'd156787: dataIn1 = 32'd5550
; 
32'd156788: dataIn1 = 32'd5551
; 
32'd156789: dataIn1 = 32'd5552
; 
32'd156790: dataIn1 = 32'd111
; 
32'd156791: dataIn1 = 32'd298
; 
32'd156792: dataIn1 = 32'd622
; 
32'd156793: dataIn1 = 32'd5468
; 
32'd156794: dataIn1 = 32'd5551
; 
32'd156795: dataIn1 = 32'd5552
; 
32'd156796: dataIn1 = 32'd5553
; 
32'd156797: dataIn1 = 32'd111
; 
32'd156798: dataIn1 = 32'd308
; 
32'd156799: dataIn1 = 32'd622
; 
32'd156800: dataIn1 = 32'd5469
; 
32'd156801: dataIn1 = 32'd5552
; 
32'd156802: dataIn1 = 32'd5553
; 
32'd156803: dataIn1 = 32'd5554
; 
32'd156804: dataIn1 = 32'd307
; 
32'd156805: dataIn1 = 32'd308
; 
32'd156806: dataIn1 = 32'd618
; 
32'd156807: dataIn1 = 32'd5469
; 
32'd156808: dataIn1 = 32'd5553
; 
32'd156809: dataIn1 = 32'd5554
; 
32'd156810: dataIn1 = 32'd5555
; 
32'd156811: dataIn1 = 32'd304
; 
32'd156812: dataIn1 = 32'd307
; 
32'd156813: dataIn1 = 32'd618
; 
32'd156814: dataIn1 = 32'd5470
; 
32'd156815: dataIn1 = 32'd5554
; 
32'd156816: dataIn1 = 32'd5555
; 
32'd156817: dataIn1 = 32'd5556
; 
32'd156818: dataIn1 = 32'd164
; 
32'd156819: dataIn1 = 32'd304
; 
32'd156820: dataIn1 = 32'd612
; 
32'd156821: dataIn1 = 32'd5470
; 
32'd156822: dataIn1 = 32'd5555
; 
32'd156823: dataIn1 = 32'd5556
; 
32'd156824: dataIn1 = 32'd5557
; 
32'd156825: dataIn1 = 32'd164
; 
32'd156826: dataIn1 = 32'd303
; 
32'd156827: dataIn1 = 32'd612
; 
32'd156828: dataIn1 = 32'd5471
; 
32'd156829: dataIn1 = 32'd5556
; 
32'd156830: dataIn1 = 32'd5557
; 
32'd156831: dataIn1 = 32'd5558
; 
32'd156832: dataIn1 = 32'd303
; 
32'd156833: dataIn1 = 32'd306
; 
32'd156834: dataIn1 = 32'd617
; 
32'd156835: dataIn1 = 32'd5471
; 
32'd156836: dataIn1 = 32'd5557
; 
32'd156837: dataIn1 = 32'd5558
; 
32'd156838: dataIn1 = 32'd5559
; 
32'd156839: dataIn1 = 32'd305
; 
32'd156840: dataIn1 = 32'd306
; 
32'd156841: dataIn1 = 32'd617
; 
32'd156842: dataIn1 = 32'd5472
; 
32'd156843: dataIn1 = 32'd5558
; 
32'd156844: dataIn1 = 32'd5559
; 
32'd156845: dataIn1 = 32'd5560
; 
32'd156846: dataIn1 = 32'd112
; 
32'd156847: dataIn1 = 32'd305
; 
32'd156848: dataIn1 = 32'd623
; 
32'd156849: dataIn1 = 32'd5472
; 
32'd156850: dataIn1 = 32'd5559
; 
32'd156851: dataIn1 = 32'd5560
; 
32'd156852: dataIn1 = 32'd5561
; 
32'd156853: dataIn1 = 32'd112
; 
32'd156854: dataIn1 = 32'd310
; 
32'd156855: dataIn1 = 32'd623
; 
32'd156856: dataIn1 = 32'd5473
; 
32'd156857: dataIn1 = 32'd5560
; 
32'd156858: dataIn1 = 32'd5561
; 
32'd156859: dataIn1 = 32'd5562
; 
32'd156860: dataIn1 = 32'd310
; 
32'd156861: dataIn1 = 32'd316
; 
32'd156862: dataIn1 = 32'd634
; 
32'd156863: dataIn1 = 32'd5473
; 
32'd156864: dataIn1 = 32'd5561
; 
32'd156865: dataIn1 = 32'd5562
; 
32'd156866: dataIn1 = 32'd5563
; 
32'd156867: dataIn1 = 32'd313
; 
32'd156868: dataIn1 = 32'd316
; 
32'd156869: dataIn1 = 32'd634
; 
32'd156870: dataIn1 = 32'd5474
; 
32'd156871: dataIn1 = 32'd5562
; 
32'd156872: dataIn1 = 32'd5563
; 
32'd156873: dataIn1 = 32'd5564
; 
32'd156874: dataIn1 = 32'd166
; 
32'd156875: dataIn1 = 32'd313
; 
32'd156876: dataIn1 = 32'd627
; 
32'd156877: dataIn1 = 32'd5474
; 
32'd156878: dataIn1 = 32'd5563
; 
32'd156879: dataIn1 = 32'd5564
; 
32'd156880: dataIn1 = 32'd5565
; 
32'd156881: dataIn1 = 32'd166
; 
32'd156882: dataIn1 = 32'd312
; 
32'd156883: dataIn1 = 32'd627
; 
32'd156884: dataIn1 = 32'd5475
; 
32'd156885: dataIn1 = 32'd5564
; 
32'd156886: dataIn1 = 32'd5565
; 
32'd156887: dataIn1 = 32'd5566
; 
32'd156888: dataIn1 = 32'd312
; 
32'd156889: dataIn1 = 32'd315
; 
32'd156890: dataIn1 = 32'd633
; 
32'd156891: dataIn1 = 32'd5475
; 
32'd156892: dataIn1 = 32'd5565
; 
32'd156893: dataIn1 = 32'd5566
; 
32'd156894: dataIn1 = 32'd5567
; 
32'd156895: dataIn1 = 32'd314
; 
32'd156896: dataIn1 = 32'd315
; 
32'd156897: dataIn1 = 32'd633
; 
32'd156898: dataIn1 = 32'd5476
; 
32'd156899: dataIn1 = 32'd5566
; 
32'd156900: dataIn1 = 32'd5567
; 
32'd156901: dataIn1 = 32'd5568
; 
32'd156902: dataIn1 = 32'd113
; 
32'd156903: dataIn1 = 32'd314
; 
32'd156904: dataIn1 = 32'd646
; 
32'd156905: dataIn1 = 32'd5476
; 
32'd156906: dataIn1 = 32'd5567
; 
32'd156907: dataIn1 = 32'd5568
; 
32'd156908: dataIn1 = 32'd5569
; 
32'd156909: dataIn1 = 32'd113
; 
32'd156910: dataIn1 = 32'd324
; 
32'd156911: dataIn1 = 32'd646
; 
32'd156912: dataIn1 = 32'd5477
; 
32'd156913: dataIn1 = 32'd5568
; 
32'd156914: dataIn1 = 32'd5569
; 
32'd156915: dataIn1 = 32'd5570
; 
32'd156916: dataIn1 = 32'd323
; 
32'd156917: dataIn1 = 32'd324
; 
32'd156918: dataIn1 = 32'd642
; 
32'd156919: dataIn1 = 32'd5477
; 
32'd156920: dataIn1 = 32'd5569
; 
32'd156921: dataIn1 = 32'd5570
; 
32'd156922: dataIn1 = 32'd5571
; 
32'd156923: dataIn1 = 32'd320
; 
32'd156924: dataIn1 = 32'd323
; 
32'd156925: dataIn1 = 32'd642
; 
32'd156926: dataIn1 = 32'd5478
; 
32'd156927: dataIn1 = 32'd5570
; 
32'd156928: dataIn1 = 32'd5571
; 
32'd156929: dataIn1 = 32'd5572
; 
32'd156930: dataIn1 = 32'd170
; 
32'd156931: dataIn1 = 32'd320
; 
32'd156932: dataIn1 = 32'd636
; 
32'd156933: dataIn1 = 32'd5478
; 
32'd156934: dataIn1 = 32'd5571
; 
32'd156935: dataIn1 = 32'd5572
; 
32'd156936: dataIn1 = 32'd5573
; 
32'd156937: dataIn1 = 32'd170
; 
32'd156938: dataIn1 = 32'd319
; 
32'd156939: dataIn1 = 32'd636
; 
32'd156940: dataIn1 = 32'd5479
; 
32'd156941: dataIn1 = 32'd5572
; 
32'd156942: dataIn1 = 32'd5573
; 
32'd156943: dataIn1 = 32'd5574
; 
32'd156944: dataIn1 = 32'd319
; 
32'd156945: dataIn1 = 32'd322
; 
32'd156946: dataIn1 = 32'd641
; 
32'd156947: dataIn1 = 32'd5479
; 
32'd156948: dataIn1 = 32'd5573
; 
32'd156949: dataIn1 = 32'd5574
; 
32'd156950: dataIn1 = 32'd5575
; 
32'd156951: dataIn1 = 32'd321
; 
32'd156952: dataIn1 = 32'd322
; 
32'd156953: dataIn1 = 32'd641
; 
32'd156954: dataIn1 = 32'd5480
; 
32'd156955: dataIn1 = 32'd5574
; 
32'd156956: dataIn1 = 32'd5575
; 
32'd156957: dataIn1 = 32'd5576
; 
32'd156958: dataIn1 = 32'd114
; 
32'd156959: dataIn1 = 32'd321
; 
32'd156960: dataIn1 = 32'd647
; 
32'd156961: dataIn1 = 32'd5480
; 
32'd156962: dataIn1 = 32'd5575
; 
32'd156963: dataIn1 = 32'd5576
; 
32'd156964: dataIn1 = 32'd5577
; 
32'd156965: dataIn1 = 32'd114
; 
32'd156966: dataIn1 = 32'd326
; 
32'd156967: dataIn1 = 32'd647
; 
32'd156968: dataIn1 = 32'd5481
; 
32'd156969: dataIn1 = 32'd5576
; 
32'd156970: dataIn1 = 32'd5577
; 
32'd156971: dataIn1 = 32'd5578
; 
32'd156972: dataIn1 = 32'd326
; 
32'd156973: dataIn1 = 32'd332
; 
32'd156974: dataIn1 = 32'd658
; 
32'd156975: dataIn1 = 32'd5481
; 
32'd156976: dataIn1 = 32'd5577
; 
32'd156977: dataIn1 = 32'd5578
; 
32'd156978: dataIn1 = 32'd5579
; 
32'd156979: dataIn1 = 32'd329
; 
32'd156980: dataIn1 = 32'd332
; 
32'd156981: dataIn1 = 32'd658
; 
32'd156982: dataIn1 = 32'd5482
; 
32'd156983: dataIn1 = 32'd5578
; 
32'd156984: dataIn1 = 32'd5579
; 
32'd156985: dataIn1 = 32'd5580
; 
32'd156986: dataIn1 = 32'd172
; 
32'd156987: dataIn1 = 32'd329
; 
32'd156988: dataIn1 = 32'd651
; 
32'd156989: dataIn1 = 32'd5482
; 
32'd156990: dataIn1 = 32'd5579
; 
32'd156991: dataIn1 = 32'd5580
; 
32'd156992: dataIn1 = 32'd5581
; 
32'd156993: dataIn1 = 32'd172
; 
32'd156994: dataIn1 = 32'd328
; 
32'd156995: dataIn1 = 32'd651
; 
32'd156996: dataIn1 = 32'd5483
; 
32'd156997: dataIn1 = 32'd5580
; 
32'd156998: dataIn1 = 32'd5581
; 
32'd156999: dataIn1 = 32'd5582
; 
32'd157000: dataIn1 = 32'd328
; 
32'd157001: dataIn1 = 32'd331
; 
32'd157002: dataIn1 = 32'd657
; 
32'd157003: dataIn1 = 32'd5483
; 
32'd157004: dataIn1 = 32'd5581
; 
32'd157005: dataIn1 = 32'd5582
; 
32'd157006: dataIn1 = 32'd5583
; 
32'd157007: dataIn1 = 32'd330
; 
32'd157008: dataIn1 = 32'd331
; 
32'd157009: dataIn1 = 32'd657
; 
32'd157010: dataIn1 = 32'd5484
; 
32'd157011: dataIn1 = 32'd5582
; 
32'd157012: dataIn1 = 32'd5583
; 
32'd157013: dataIn1 = 32'd5584
; 
32'd157014: dataIn1 = 32'd115
; 
32'd157015: dataIn1 = 32'd330
; 
32'd157016: dataIn1 = 32'd670
; 
32'd157017: dataIn1 = 32'd5484
; 
32'd157018: dataIn1 = 32'd5583
; 
32'd157019: dataIn1 = 32'd5584
; 
32'd157020: dataIn1 = 32'd5585
; 
32'd157021: dataIn1 = 32'd115
; 
32'd157022: dataIn1 = 32'd340
; 
32'd157023: dataIn1 = 32'd670
; 
32'd157024: dataIn1 = 32'd5485
; 
32'd157025: dataIn1 = 32'd5584
; 
32'd157026: dataIn1 = 32'd5585
; 
32'd157027: dataIn1 = 32'd5586
; 
32'd157028: dataIn1 = 32'd339
; 
32'd157029: dataIn1 = 32'd340
; 
32'd157030: dataIn1 = 32'd666
; 
32'd157031: dataIn1 = 32'd5485
; 
32'd157032: dataIn1 = 32'd5585
; 
32'd157033: dataIn1 = 32'd5586
; 
32'd157034: dataIn1 = 32'd5587
; 
32'd157035: dataIn1 = 32'd336
; 
32'd157036: dataIn1 = 32'd339
; 
32'd157037: dataIn1 = 32'd666
; 
32'd157038: dataIn1 = 32'd5486
; 
32'd157039: dataIn1 = 32'd5586
; 
32'd157040: dataIn1 = 32'd5587
; 
32'd157041: dataIn1 = 32'd5588
; 
32'd157042: dataIn1 = 32'd176
; 
32'd157043: dataIn1 = 32'd336
; 
32'd157044: dataIn1 = 32'd660
; 
32'd157045: dataIn1 = 32'd5486
; 
32'd157046: dataIn1 = 32'd5587
; 
32'd157047: dataIn1 = 32'd5588
; 
32'd157048: dataIn1 = 32'd5589
; 
32'd157049: dataIn1 = 32'd176
; 
32'd157050: dataIn1 = 32'd335
; 
32'd157051: dataIn1 = 32'd660
; 
32'd157052: dataIn1 = 32'd5487
; 
32'd157053: dataIn1 = 32'd5588
; 
32'd157054: dataIn1 = 32'd5589
; 
32'd157055: dataIn1 = 32'd5590
; 
32'd157056: dataIn1 = 32'd335
; 
32'd157057: dataIn1 = 32'd338
; 
32'd157058: dataIn1 = 32'd665
; 
32'd157059: dataIn1 = 32'd5487
; 
32'd157060: dataIn1 = 32'd5589
; 
32'd157061: dataIn1 = 32'd5590
; 
32'd157062: dataIn1 = 32'd5591
; 
32'd157063: dataIn1 = 32'd337
; 
32'd157064: dataIn1 = 32'd338
; 
32'd157065: dataIn1 = 32'd665
; 
32'd157066: dataIn1 = 32'd5488
; 
32'd157067: dataIn1 = 32'd5590
; 
32'd157068: dataIn1 = 32'd5591
; 
32'd157069: dataIn1 = 32'd5592
; 
32'd157070: dataIn1 = 32'd116
; 
32'd157071: dataIn1 = 32'd337
; 
32'd157072: dataIn1 = 32'd671
; 
32'd157073: dataIn1 = 32'd5488
; 
32'd157074: dataIn1 = 32'd5591
; 
32'd157075: dataIn1 = 32'd5592
; 
32'd157076: dataIn1 = 32'd5593
; 
32'd157077: dataIn1 = 32'd116
; 
32'd157078: dataIn1 = 32'd342
; 
32'd157079: dataIn1 = 32'd671
; 
32'd157080: dataIn1 = 32'd5489
; 
32'd157081: dataIn1 = 32'd5592
; 
32'd157082: dataIn1 = 32'd5593
; 
32'd157083: dataIn1 = 32'd5594
; 
32'd157084: dataIn1 = 32'd342
; 
32'd157085: dataIn1 = 32'd348
; 
32'd157086: dataIn1 = 32'd682
; 
32'd157087: dataIn1 = 32'd5489
; 
32'd157088: dataIn1 = 32'd5593
; 
32'd157089: dataIn1 = 32'd5594
; 
32'd157090: dataIn1 = 32'd5595
; 
32'd157091: dataIn1 = 32'd345
; 
32'd157092: dataIn1 = 32'd348
; 
32'd157093: dataIn1 = 32'd682
; 
32'd157094: dataIn1 = 32'd5490
; 
32'd157095: dataIn1 = 32'd5594
; 
32'd157096: dataIn1 = 32'd5595
; 
32'd157097: dataIn1 = 32'd5596
; 
32'd157098: dataIn1 = 32'd178
; 
32'd157099: dataIn1 = 32'd345
; 
32'd157100: dataIn1 = 32'd675
; 
32'd157101: dataIn1 = 32'd5490
; 
32'd157102: dataIn1 = 32'd5595
; 
32'd157103: dataIn1 = 32'd5596
; 
32'd157104: dataIn1 = 32'd5597
; 
32'd157105: dataIn1 = 32'd178
; 
32'd157106: dataIn1 = 32'd344
; 
32'd157107: dataIn1 = 32'd675
; 
32'd157108: dataIn1 = 32'd5491
; 
32'd157109: dataIn1 = 32'd5596
; 
32'd157110: dataIn1 = 32'd5597
; 
32'd157111: dataIn1 = 32'd5598
; 
32'd157112: dataIn1 = 32'd344
; 
32'd157113: dataIn1 = 32'd347
; 
32'd157114: dataIn1 = 32'd681
; 
32'd157115: dataIn1 = 32'd5491
; 
32'd157116: dataIn1 = 32'd5597
; 
32'd157117: dataIn1 = 32'd5598
; 
32'd157118: dataIn1 = 32'd5599
; 
32'd157119: dataIn1 = 32'd346
; 
32'd157120: dataIn1 = 32'd347
; 
32'd157121: dataIn1 = 32'd681
; 
32'd157122: dataIn1 = 32'd5492
; 
32'd157123: dataIn1 = 32'd5598
; 
32'd157124: dataIn1 = 32'd5599
; 
32'd157125: dataIn1 = 32'd5600
; 
32'd157126: dataIn1 = 32'd117
; 
32'd157127: dataIn1 = 32'd346
; 
32'd157128: dataIn1 = 32'd694
; 
32'd157129: dataIn1 = 32'd5492
; 
32'd157130: dataIn1 = 32'd5599
; 
32'd157131: dataIn1 = 32'd5600
; 
32'd157132: dataIn1 = 32'd5601
; 
32'd157133: dataIn1 = 32'd117
; 
32'd157134: dataIn1 = 32'd356
; 
32'd157135: dataIn1 = 32'd694
; 
32'd157136: dataIn1 = 32'd5493
; 
32'd157137: dataIn1 = 32'd5600
; 
32'd157138: dataIn1 = 32'd5601
; 
32'd157139: dataIn1 = 32'd5602
; 
32'd157140: dataIn1 = 32'd355
; 
32'd157141: dataIn1 = 32'd356
; 
32'd157142: dataIn1 = 32'd690
; 
32'd157143: dataIn1 = 32'd5493
; 
32'd157144: dataIn1 = 32'd5601
; 
32'd157145: dataIn1 = 32'd5602
; 
32'd157146: dataIn1 = 32'd5603
; 
32'd157147: dataIn1 = 32'd352
; 
32'd157148: dataIn1 = 32'd355
; 
32'd157149: dataIn1 = 32'd690
; 
32'd157150: dataIn1 = 32'd5494
; 
32'd157151: dataIn1 = 32'd5602
; 
32'd157152: dataIn1 = 32'd5603
; 
32'd157153: dataIn1 = 32'd5604
; 
32'd157154: dataIn1 = 32'd182
; 
32'd157155: dataIn1 = 32'd352
; 
32'd157156: dataIn1 = 32'd684
; 
32'd157157: dataIn1 = 32'd5494
; 
32'd157158: dataIn1 = 32'd5603
; 
32'd157159: dataIn1 = 32'd5604
; 
32'd157160: dataIn1 = 32'd5605
; 
32'd157161: dataIn1 = 32'd182
; 
32'd157162: dataIn1 = 32'd351
; 
32'd157163: dataIn1 = 32'd684
; 
32'd157164: dataIn1 = 32'd5495
; 
32'd157165: dataIn1 = 32'd5604
; 
32'd157166: dataIn1 = 32'd5605
; 
32'd157167: dataIn1 = 32'd5606
; 
32'd157168: dataIn1 = 32'd351
; 
32'd157169: dataIn1 = 32'd354
; 
32'd157170: dataIn1 = 32'd689
; 
32'd157171: dataIn1 = 32'd5495
; 
32'd157172: dataIn1 = 32'd5605
; 
32'd157173: dataIn1 = 32'd5606
; 
32'd157174: dataIn1 = 32'd5607
; 
32'd157175: dataIn1 = 32'd353
; 
32'd157176: dataIn1 = 32'd354
; 
32'd157177: dataIn1 = 32'd689
; 
32'd157178: dataIn1 = 32'd5496
; 
32'd157179: dataIn1 = 32'd5606
; 
32'd157180: dataIn1 = 32'd5607
; 
32'd157181: dataIn1 = 32'd5608
; 
32'd157182: dataIn1 = 32'd118
; 
32'd157183: dataIn1 = 32'd353
; 
32'd157184: dataIn1 = 32'd695
; 
32'd157185: dataIn1 = 32'd5496
; 
32'd157186: dataIn1 = 32'd5607
; 
32'd157187: dataIn1 = 32'd5608
; 
32'd157188: dataIn1 = 32'd5609
; 
32'd157189: dataIn1 = 32'd118
; 
32'd157190: dataIn1 = 32'd358
; 
32'd157191: dataIn1 = 32'd695
; 
32'd157192: dataIn1 = 32'd5497
; 
32'd157193: dataIn1 = 32'd5608
; 
32'd157194: dataIn1 = 32'd5609
; 
32'd157195: dataIn1 = 32'd5610
; 
32'd157196: dataIn1 = 32'd358
; 
32'd157197: dataIn1 = 32'd364
; 
32'd157198: dataIn1 = 32'd706
; 
32'd157199: dataIn1 = 32'd5497
; 
32'd157200: dataIn1 = 32'd5609
; 
32'd157201: dataIn1 = 32'd5610
; 
32'd157202: dataIn1 = 32'd5611
; 
32'd157203: dataIn1 = 32'd361
; 
32'd157204: dataIn1 = 32'd364
; 
32'd157205: dataIn1 = 32'd706
; 
32'd157206: dataIn1 = 32'd5498
; 
32'd157207: dataIn1 = 32'd5610
; 
32'd157208: dataIn1 = 32'd5611
; 
32'd157209: dataIn1 = 32'd5612
; 
32'd157210: dataIn1 = 32'd184
; 
32'd157211: dataIn1 = 32'd361
; 
32'd157212: dataIn1 = 32'd699
; 
32'd157213: dataIn1 = 32'd5498
; 
32'd157214: dataIn1 = 32'd5611
; 
32'd157215: dataIn1 = 32'd5612
; 
32'd157216: dataIn1 = 32'd5613
; 
32'd157217: dataIn1 = 32'd184
; 
32'd157218: dataIn1 = 32'd360
; 
32'd157219: dataIn1 = 32'd699
; 
32'd157220: dataIn1 = 32'd5499
; 
32'd157221: dataIn1 = 32'd5612
; 
32'd157222: dataIn1 = 32'd5613
; 
32'd157223: dataIn1 = 32'd5614
; 
32'd157224: dataIn1 = 32'd360
; 
32'd157225: dataIn1 = 32'd363
; 
32'd157226: dataIn1 = 32'd705
; 
32'd157227: dataIn1 = 32'd5499
; 
32'd157228: dataIn1 = 32'd5613
; 
32'd157229: dataIn1 = 32'd5614
; 
32'd157230: dataIn1 = 32'd5615
; 
32'd157231: dataIn1 = 32'd362
; 
32'd157232: dataIn1 = 32'd363
; 
32'd157233: dataIn1 = 32'd705
; 
32'd157234: dataIn1 = 32'd5500
; 
32'd157235: dataIn1 = 32'd5614
; 
32'd157236: dataIn1 = 32'd5615
; 
32'd157237: dataIn1 = 32'd5616
; 
32'd157238: dataIn1 = 32'd119
; 
32'd157239: dataIn1 = 32'd362
; 
32'd157240: dataIn1 = 32'd718
; 
32'd157241: dataIn1 = 32'd5500
; 
32'd157242: dataIn1 = 32'd5615
; 
32'd157243: dataIn1 = 32'd5616
; 
32'd157244: dataIn1 = 32'd5617
; 
32'd157245: dataIn1 = 32'd119
; 
32'd157246: dataIn1 = 32'd372
; 
32'd157247: dataIn1 = 32'd718
; 
32'd157248: dataIn1 = 32'd5501
; 
32'd157249: dataIn1 = 32'd5616
; 
32'd157250: dataIn1 = 32'd5617
; 
32'd157251: dataIn1 = 32'd5618
; 
32'd157252: dataIn1 = 32'd371
; 
32'd157253: dataIn1 = 32'd372
; 
32'd157254: dataIn1 = 32'd714
; 
32'd157255: dataIn1 = 32'd5501
; 
32'd157256: dataIn1 = 32'd5617
; 
32'd157257: dataIn1 = 32'd5618
; 
32'd157258: dataIn1 = 32'd5619
; 
32'd157259: dataIn1 = 32'd368
; 
32'd157260: dataIn1 = 32'd371
; 
32'd157261: dataIn1 = 32'd714
; 
32'd157262: dataIn1 = 32'd5502
; 
32'd157263: dataIn1 = 32'd5618
; 
32'd157264: dataIn1 = 32'd5619
; 
32'd157265: dataIn1 = 32'd5620
; 
32'd157266: dataIn1 = 32'd188
; 
32'd157267: dataIn1 = 32'd368
; 
32'd157268: dataIn1 = 32'd708
; 
32'd157269: dataIn1 = 32'd5502
; 
32'd157270: dataIn1 = 32'd5619
; 
32'd157271: dataIn1 = 32'd5620
; 
32'd157272: dataIn1 = 32'd5621
; 
32'd157273: dataIn1 = 32'd188
; 
32'd157274: dataIn1 = 32'd367
; 
32'd157275: dataIn1 = 32'd708
; 
32'd157276: dataIn1 = 32'd5503
; 
32'd157277: dataIn1 = 32'd5620
; 
32'd157278: dataIn1 = 32'd5621
; 
32'd157279: dataIn1 = 32'd5622
; 
32'd157280: dataIn1 = 32'd367
; 
32'd157281: dataIn1 = 32'd370
; 
32'd157282: dataIn1 = 32'd713
; 
32'd157283: dataIn1 = 32'd5503
; 
32'd157284: dataIn1 = 32'd5621
; 
32'd157285: dataIn1 = 32'd5622
; 
32'd157286: dataIn1 = 32'd5623
; 
32'd157287: dataIn1 = 32'd369
; 
32'd157288: dataIn1 = 32'd370
; 
32'd157289: dataIn1 = 32'd713
; 
32'd157290: dataIn1 = 32'd5504
; 
32'd157291: dataIn1 = 32'd5622
; 
32'd157292: dataIn1 = 32'd5623
; 
32'd157293: dataIn1 = 32'd5624
; 
32'd157294: dataIn1 = 32'd120
; 
32'd157295: dataIn1 = 32'd369
; 
32'd157296: dataIn1 = 32'd719
; 
32'd157297: dataIn1 = 32'd5504
; 
32'd157298: dataIn1 = 32'd5623
; 
32'd157299: dataIn1 = 32'd5624
; 
32'd157300: dataIn1 = 32'd5625
; 
32'd157301: dataIn1 = 32'd120
; 
32'd157302: dataIn1 = 32'd374
; 
32'd157303: dataIn1 = 32'd719
; 
32'd157304: dataIn1 = 32'd5505
; 
32'd157305: dataIn1 = 32'd5624
; 
32'd157306: dataIn1 = 32'd5625
; 
32'd157307: dataIn1 = 32'd5626
; 
32'd157308: dataIn1 = 32'd374
; 
32'd157309: dataIn1 = 32'd380
; 
32'd157310: dataIn1 = 32'd730
; 
32'd157311: dataIn1 = 32'd5505
; 
32'd157312: dataIn1 = 32'd5625
; 
32'd157313: dataIn1 = 32'd5626
; 
32'd157314: dataIn1 = 32'd5627
; 
32'd157315: dataIn1 = 32'd377
; 
32'd157316: dataIn1 = 32'd380
; 
32'd157317: dataIn1 = 32'd730
; 
32'd157318: dataIn1 = 32'd5506
; 
32'd157319: dataIn1 = 32'd5626
; 
32'd157320: dataIn1 = 32'd5627
; 
32'd157321: dataIn1 = 32'd5628
; 
32'd157322: dataIn1 = 32'd190
; 
32'd157323: dataIn1 = 32'd377
; 
32'd157324: dataIn1 = 32'd723
; 
32'd157325: dataIn1 = 32'd5506
; 
32'd157326: dataIn1 = 32'd5627
; 
32'd157327: dataIn1 = 32'd5628
; 
32'd157328: dataIn1 = 32'd5629
; 
32'd157329: dataIn1 = 32'd190
; 
32'd157330: dataIn1 = 32'd376
; 
32'd157331: dataIn1 = 32'd723
; 
32'd157332: dataIn1 = 32'd5507
; 
32'd157333: dataIn1 = 32'd5628
; 
32'd157334: dataIn1 = 32'd5629
; 
32'd157335: dataIn1 = 32'd5630
; 
32'd157336: dataIn1 = 32'd376
; 
32'd157337: dataIn1 = 32'd379
; 
32'd157338: dataIn1 = 32'd729
; 
32'd157339: dataIn1 = 32'd5507
; 
32'd157340: dataIn1 = 32'd5629
; 
32'd157341: dataIn1 = 32'd5630
; 
32'd157342: dataIn1 = 32'd5631
; 
32'd157343: dataIn1 = 32'd378
; 
32'd157344: dataIn1 = 32'd379
; 
32'd157345: dataIn1 = 32'd729
; 
32'd157346: dataIn1 = 32'd5508
; 
32'd157347: dataIn1 = 32'd5630
; 
32'd157348: dataIn1 = 32'd5631
; 
32'd157349: dataIn1 = 32'd5632
; 
32'd157350: dataIn1 = 32'd121
; 
32'd157351: dataIn1 = 32'd378
; 
32'd157352: dataIn1 = 32'd5508
; 
32'd157353: dataIn1 = 32'd5631
; 
32'd157354: dataIn1 = 32'd5632
; 
32'd157355: dataIn1 = 32'd451
; 
32'd157356: dataIn1 = 32'd2739
; 
32'd157357: dataIn1 = 32'd5273
; 
32'd157358: dataIn1 = 32'd5323
; 
32'd157359: dataIn1 = 32'd5633
; 
32'd157360: dataIn1 = 32'd5634
; 
32'd157361: dataIn1 = 32'd6691
; 
32'd157362: dataIn1 = 32'd2738
; 
32'd157363: dataIn1 = 32'd2739
; 
32'd157364: dataIn1 = 32'd2740
; 
32'd157365: dataIn1 = 32'd5273
; 
32'd157366: dataIn1 = 32'd5633
; 
32'd157367: dataIn1 = 32'd5634
; 
32'd157368: dataIn1 = 32'd5635
; 
32'd157369: dataIn1 = 32'd9343
; 
32'd157370: dataIn1 = 32'd9344
; 
32'd157371: dataIn1 = 32'd9352
; 
32'd157372: dataIn1 = 32'd9359
; 
32'd157373: dataIn1 = 32'd9366
; 
32'd157374: dataIn1 = 32'd9367
; 
32'd157375: dataIn1 = 32'd5636
; 
32'd157376: dataIn1 = 32'd6806
; 
32'd157377: dataIn1 = 32'd9345
; 
32'd157378: dataIn1 = 32'd9346
; 
32'd157379: dataIn1 = 32'd9360
; 
32'd157380: dataIn1 = 32'd9383
; 
32'd157381: dataIn1 = 32'd5637
; 
32'd157382: dataIn1 = 32'd6821
; 
32'd157383: dataIn1 = 32'd9347
; 
32'd157384: dataIn1 = 32'd9348
; 
32'd157385: dataIn1 = 32'd9355
; 
32'd157386: dataIn1 = 32'd9390
; 
32'd157387: dataIn1 = 32'd5638
; 
32'd157388: dataIn1 = 32'd9370
; 
32'd157389: dataIn1 = 32'd9371
; 
32'd157390: dataIn1 = 32'd9376
; 
32'd157391: dataIn1 = 32'd9810
; 
32'd157392: dataIn1 = 32'd5639
; 
32'd157393: dataIn1 = 32'd6816
; 
32'd157394: dataIn1 = 32'd6817
; 
32'd157395: dataIn1 = 32'd6819
; 
32'd157396: dataIn1 = 32'd6820
; 
32'd157397: dataIn1 = 32'd9263
; 
32'd157398: dataIn1 = 32'd5640
; 
32'd157399: dataIn1 = 32'd6827
; 
32'd157400: dataIn1 = 32'd9387
; 
32'd157401: dataIn1 = 32'd9388
; 
32'd157402: dataIn1 = 32'd5641
; 
32'd157403: dataIn1 = 32'd6821
; 
32'd157404: dataIn1 = 32'd6823
; 
32'd157405: dataIn1 = 32'd6824
; 
32'd157406: dataIn1 = 32'd6826
; 
32'd157407: dataIn1 = 32'd9264
; 
32'd157408: dataIn1 = 32'd5642
; 
32'd157409: dataIn1 = 32'd9394
; 
32'd157410: dataIn1 = 32'd9395
; 
32'd157411: dataIn1 = 32'd9403
; 
32'd157412: dataIn1 = 32'd9410
; 
32'd157413: dataIn1 = 32'd9417
; 
32'd157414: dataIn1 = 32'd9418
; 
32'd157415: dataIn1 = 32'd5643
; 
32'd157416: dataIn1 = 32'd6842
; 
32'd157417: dataIn1 = 32'd9396
; 
32'd157418: dataIn1 = 32'd9397
; 
32'd157419: dataIn1 = 32'd9411
; 
32'd157420: dataIn1 = 32'd9440
; 
32'd157421: dataIn1 = 32'd5644
; 
32'd157422: dataIn1 = 32'd6831
; 
32'd157423: dataIn1 = 32'd9398
; 
32'd157424: dataIn1 = 32'd9399
; 
32'd157425: dataIn1 = 32'd9406
; 
32'd157426: dataIn1 = 32'd9445
; 
32'd157427: dataIn1 = 32'd5645
; 
32'd157428: dataIn1 = 32'd9419
; 
32'd157429: dataIn1 = 32'd9420
; 
32'd157430: dataIn1 = 32'd9426
; 
32'd157431: dataIn1 = 32'd9433
; 
32'd157432: dataIn1 = 32'd5646
; 
32'd157433: dataIn1 = 32'd9438
; 
32'd157434: dataIn1 = 32'd9439
; 
32'd157435: dataIn1 = 32'd10291
; 
32'd157436: dataIn1 = 32'd2105
; 
32'd157437: dataIn1 = 32'd5647
; 
32'd157438: dataIn1 = 32'd6842
; 
32'd157439: dataIn1 = 32'd6843
; 
32'd157440: dataIn1 = 32'd6845
; 
32'd157441: dataIn1 = 32'd9266
; 
32'd157442: dataIn1 = 32'd5648
; 
32'd157443: dataIn1 = 32'd6847
; 
32'd157444: dataIn1 = 32'd6849
; 
32'd157445: dataIn1 = 32'd6850
; 
32'd157446: dataIn1 = 32'd9257
; 
32'd157447: dataIn1 = 32'd9269
; 
32'd157448: dataIn1 = 32'd2296
; 
32'd157449: dataIn1 = 32'd3872
; 
32'd157450: dataIn1 = 32'd3873
; 
32'd157451: dataIn1 = 32'd5649
; 
32'd157452: dataIn1 = 32'd5650
; 
32'd157453: dataIn1 = 32'd5651
; 
32'd157454: dataIn1 = 32'd3871
; 
32'd157455: dataIn1 = 32'd3873
; 
32'd157456: dataIn1 = 32'd5649
; 
32'd157457: dataIn1 = 32'd5650
; 
32'd157458: dataIn1 = 32'd5651
; 
32'd157459: dataIn1 = 32'd5652
; 
32'd157460: dataIn1 = 32'd5653
; 
32'd157461: dataIn1 = 32'd3871
; 
32'd157462: dataIn1 = 32'd3872
; 
32'd157463: dataIn1 = 32'd5649
; 
32'd157464: dataIn1 = 32'd5650
; 
32'd157465: dataIn1 = 32'd5651
; 
32'd157466: dataIn1 = 32'd5654
; 
32'd157467: dataIn1 = 32'd5655
; 
32'd157468: dataIn1 = 32'd2297
; 
32'd157469: dataIn1 = 32'd3873
; 
32'd157470: dataIn1 = 32'd5650
; 
32'd157471: dataIn1 = 32'd5652
; 
32'd157472: dataIn1 = 32'd5653
; 
32'd157473: dataIn1 = 32'd5663
; 
32'd157474: dataIn1 = 32'd5664
; 
32'd157475: dataIn1 = 32'd2297
; 
32'd157476: dataIn1 = 32'd3871
; 
32'd157477: dataIn1 = 32'd5650
; 
32'd157478: dataIn1 = 32'd5652
; 
32'd157479: dataIn1 = 32'd5653
; 
32'd157480: dataIn1 = 32'd5657
; 
32'd157481: dataIn1 = 32'd5659
; 
32'd157482: dataIn1 = 32'd2298
; 
32'd157483: dataIn1 = 32'd3872
; 
32'd157484: dataIn1 = 32'd5651
; 
32'd157485: dataIn1 = 32'd5654
; 
32'd157486: dataIn1 = 32'd5655
; 
32'd157487: dataIn1 = 32'd5661
; 
32'd157488: dataIn1 = 32'd5662
; 
32'd157489: dataIn1 = 32'd2298
; 
32'd157490: dataIn1 = 32'd3871
; 
32'd157491: dataIn1 = 32'd5651
; 
32'd157492: dataIn1 = 32'd5654
; 
32'd157493: dataIn1 = 32'd5655
; 
32'd157494: dataIn1 = 32'd5658
; 
32'd157495: dataIn1 = 32'd5660
; 
32'd157496: dataIn1 = 32'd205
; 
32'd157497: dataIn1 = 32'd3874
; 
32'd157498: dataIn1 = 32'd3875
; 
32'd157499: dataIn1 = 32'd5656
; 
32'd157500: dataIn1 = 32'd5657
; 
32'd157501: dataIn1 = 32'd5658
; 
32'd157502: dataIn1 = 32'd3871
; 
32'd157503: dataIn1 = 32'd3875
; 
32'd157504: dataIn1 = 32'd5653
; 
32'd157505: dataIn1 = 32'd5656
; 
32'd157506: dataIn1 = 32'd5657
; 
32'd157507: dataIn1 = 32'd5658
; 
32'd157508: dataIn1 = 32'd5659
; 
32'd157509: dataIn1 = 32'd3871
; 
32'd157510: dataIn1 = 32'd3874
; 
32'd157511: dataIn1 = 32'd5655
; 
32'd157512: dataIn1 = 32'd5656
; 
32'd157513: dataIn1 = 32'd5657
; 
32'd157514: dataIn1 = 32'd5658
; 
32'd157515: dataIn1 = 32'd5660
; 
32'd157516: dataIn1 = 32'd2297
; 
32'd157517: dataIn1 = 32'd3875
; 
32'd157518: dataIn1 = 32'd5653
; 
32'd157519: dataIn1 = 32'd5657
; 
32'd157520: dataIn1 = 32'd5659
; 
32'd157521: dataIn1 = 32'd5670
; 
32'd157522: dataIn1 = 32'd5671
; 
32'd157523: dataIn1 = 32'd2298
; 
32'd157524: dataIn1 = 32'd3874
; 
32'd157525: dataIn1 = 32'd5655
; 
32'd157526: dataIn1 = 32'd5658
; 
32'd157527: dataIn1 = 32'd5660
; 
32'd157528: dataIn1 = 32'd5685
; 
32'd157529: dataIn1 = 32'd5686
; 
32'd157530: dataIn1 = 32'd2298
; 
32'd157531: dataIn1 = 32'd3876
; 
32'd157532: dataIn1 = 32'd5654
; 
32'd157533: dataIn1 = 32'd5661
; 
32'd157534: dataIn1 = 32'd5662
; 
32'd157535: dataIn1 = 32'd5684
; 
32'd157536: dataIn1 = 32'd5687
; 
32'd157537: dataIn1 = 32'd3872
; 
32'd157538: dataIn1 = 32'd3876
; 
32'd157539: dataIn1 = 32'd3877
; 
32'd157540: dataIn1 = 32'd5654
; 
32'd157541: dataIn1 = 32'd5661
; 
32'd157542: dataIn1 = 32'd5662
; 
32'd157543: dataIn1 = 32'd3873
; 
32'd157544: dataIn1 = 32'd3878
; 
32'd157545: dataIn1 = 32'd3879
; 
32'd157546: dataIn1 = 32'd5652
; 
32'd157547: dataIn1 = 32'd5663
; 
32'd157548: dataIn1 = 32'd5664
; 
32'd157549: dataIn1 = 32'd2297
; 
32'd157550: dataIn1 = 32'd3878
; 
32'd157551: dataIn1 = 32'd5652
; 
32'd157552: dataIn1 = 32'd5663
; 
32'd157553: dataIn1 = 32'd5664
; 
32'd157554: dataIn1 = 32'd5668
; 
32'd157555: dataIn1 = 32'd5673
; 
32'd157556: dataIn1 = 32'd3880
; 
32'd157557: dataIn1 = 32'd3883
; 
32'd157558: dataIn1 = 32'd3884
; 
32'd157559: dataIn1 = 32'd5665
; 
32'd157560: dataIn1 = 32'd5666
; 
32'd157561: dataIn1 = 32'd5667
; 
32'd157562: dataIn1 = 32'd127
; 
32'd157563: dataIn1 = 32'd3884
; 
32'd157564: dataIn1 = 32'd5665
; 
32'd157565: dataIn1 = 32'd5666
; 
32'd157566: dataIn1 = 32'd5667
; 
32'd157567: dataIn1 = 32'd5784
; 
32'd157568: dataIn1 = 32'd5787
; 
32'd157569: dataIn1 = 32'd127
; 
32'd157570: dataIn1 = 32'd3883
; 
32'd157571: dataIn1 = 32'd5665
; 
32'd157572: dataIn1 = 32'd5666
; 
32'd157573: dataIn1 = 32'd5667
; 
32'd157574: dataIn1 = 32'd5941
; 
32'd157575: dataIn1 = 32'd5944
; 
32'd157576: dataIn1 = 32'd2297
; 
32'd157577: dataIn1 = 32'd3889
; 
32'd157578: dataIn1 = 32'd5664
; 
32'd157579: dataIn1 = 32'd5668
; 
32'd157580: dataIn1 = 32'd5669
; 
32'd157581: dataIn1 = 32'd5670
; 
32'd157582: dataIn1 = 32'd5673
; 
32'd157583: dataIn1 = 32'd3887
; 
32'd157584: dataIn1 = 32'd3888
; 
32'd157585: dataIn1 = 32'd3889
; 
32'd157586: dataIn1 = 32'd5668
; 
32'd157587: dataIn1 = 32'd5669
; 
32'd157588: dataIn1 = 32'd5670
; 
32'd157589: dataIn1 = 32'd2297
; 
32'd157590: dataIn1 = 32'd3887
; 
32'd157591: dataIn1 = 32'd5659
; 
32'd157592: dataIn1 = 32'd5668
; 
32'd157593: dataIn1 = 32'd5669
; 
32'd157594: dataIn1 = 32'd5670
; 
32'd157595: dataIn1 = 32'd5671
; 
32'd157596: dataIn1 = 32'd3875
; 
32'd157597: dataIn1 = 32'd3887
; 
32'd157598: dataIn1 = 32'd3890
; 
32'd157599: dataIn1 = 32'd5659
; 
32'd157600: dataIn1 = 32'd5670
; 
32'd157601: dataIn1 = 32'd5671
; 
32'd157602: dataIn1 = 32'd3889
; 
32'd157603: dataIn1 = 32'd3893
; 
32'd157604: dataIn1 = 32'd5672
; 
32'd157605: dataIn1 = 32'd5673
; 
32'd157606: dataIn1 = 32'd5674
; 
32'd157607: dataIn1 = 32'd5675
; 
32'd157608: dataIn1 = 32'd5676
; 
32'd157609: dataIn1 = 32'd3878
; 
32'd157610: dataIn1 = 32'd3889
; 
32'd157611: dataIn1 = 32'd5664
; 
32'd157612: dataIn1 = 32'd5668
; 
32'd157613: dataIn1 = 32'd5672
; 
32'd157614: dataIn1 = 32'd5673
; 
32'd157615: dataIn1 = 32'd5674
; 
32'd157616: dataIn1 = 32'd445
; 
32'd157617: dataIn1 = 32'd3878
; 
32'd157618: dataIn1 = 32'd3893
; 
32'd157619: dataIn1 = 32'd5672
; 
32'd157620: dataIn1 = 32'd5673
; 
32'd157621: dataIn1 = 32'd5674
; 
32'd157622: dataIn1 = 32'd2301
; 
32'd157623: dataIn1 = 32'd3888
; 
32'd157624: dataIn1 = 32'd3889
; 
32'd157625: dataIn1 = 32'd5672
; 
32'd157626: dataIn1 = 32'd5675
; 
32'd157627: dataIn1 = 32'd5676
; 
32'd157628: dataIn1 = 32'd2301
; 
32'd157629: dataIn1 = 32'd3893
; 
32'd157630: dataIn1 = 32'd5672
; 
32'd157631: dataIn1 = 32'd5675
; 
32'd157632: dataIn1 = 32'd5676
; 
32'd157633: dataIn1 = 32'd5799
; 
32'd157634: dataIn1 = 32'd5804
; 
32'd157635: dataIn1 = 32'd3895
; 
32'd157636: dataIn1 = 32'd3896
; 
32'd157637: dataIn1 = 32'd5677
; 
32'd157638: dataIn1 = 32'd5678
; 
32'd157639: dataIn1 = 32'd5679
; 
32'd157640: dataIn1 = 32'd5680
; 
32'd157641: dataIn1 = 32'd5681
; 
32'd157642: dataIn1 = 32'd3894
; 
32'd157643: dataIn1 = 32'd3896
; 
32'd157644: dataIn1 = 32'd5677
; 
32'd157645: dataIn1 = 32'd5678
; 
32'd157646: dataIn1 = 32'd5679
; 
32'd157647: dataIn1 = 32'd5682
; 
32'd157648: dataIn1 = 32'd5683
; 
32'd157649: dataIn1 = 32'd3894
; 
32'd157650: dataIn1 = 32'd3895
; 
32'd157651: dataIn1 = 32'd5677
; 
32'd157652: dataIn1 = 32'd5678
; 
32'd157653: dataIn1 = 32'd5679
; 
32'd157654: dataIn1 = 32'd5684
; 
32'd157655: dataIn1 = 32'd5685
; 
32'd157656: dataIn1 = 32'd2302
; 
32'd157657: dataIn1 = 32'd3896
; 
32'd157658: dataIn1 = 32'd5677
; 
32'd157659: dataIn1 = 32'd5680
; 
32'd157660: dataIn1 = 32'd5681
; 
32'd157661: dataIn1 = 32'd5688
; 
32'd157662: dataIn1 = 32'd5691
; 
32'd157663: dataIn1 = 32'd2302
; 
32'd157664: dataIn1 = 32'd3895
; 
32'd157665: dataIn1 = 32'd3898
; 
32'd157666: dataIn1 = 32'd5677
; 
32'd157667: dataIn1 = 32'd5680
; 
32'd157668: dataIn1 = 32'd5681
; 
32'd157669: dataIn1 = 32'd400
; 
32'd157670: dataIn1 = 32'd3896
; 
32'd157671: dataIn1 = 32'd5678
; 
32'd157672: dataIn1 = 32'd5682
; 
32'd157673: dataIn1 = 32'd5683
; 
32'd157674: dataIn1 = 32'd5689
; 
32'd157675: dataIn1 = 32'd5692
; 
32'd157676: dataIn1 = 32'd400
; 
32'd157677: dataIn1 = 32'd3894
; 
32'd157678: dataIn1 = 32'd3897
; 
32'd157679: dataIn1 = 32'd5678
; 
32'd157680: dataIn1 = 32'd5682
; 
32'd157681: dataIn1 = 32'd5683
; 
32'd157682: dataIn1 = 32'd2298
; 
32'd157683: dataIn1 = 32'd3895
; 
32'd157684: dataIn1 = 32'd5661
; 
32'd157685: dataIn1 = 32'd5679
; 
32'd157686: dataIn1 = 32'd5684
; 
32'd157687: dataIn1 = 32'd5685
; 
32'd157688: dataIn1 = 32'd5687
; 
32'd157689: dataIn1 = 32'd2298
; 
32'd157690: dataIn1 = 32'd3894
; 
32'd157691: dataIn1 = 32'd5660
; 
32'd157692: dataIn1 = 32'd5679
; 
32'd157693: dataIn1 = 32'd5684
; 
32'd157694: dataIn1 = 32'd5685
; 
32'd157695: dataIn1 = 32'd5686
; 
32'd157696: dataIn1 = 32'd3874
; 
32'd157697: dataIn1 = 32'd3894
; 
32'd157698: dataIn1 = 32'd3897
; 
32'd157699: dataIn1 = 32'd5660
; 
32'd157700: dataIn1 = 32'd5685
; 
32'd157701: dataIn1 = 32'd5686
; 
32'd157702: dataIn1 = 32'd3876
; 
32'd157703: dataIn1 = 32'd3895
; 
32'd157704: dataIn1 = 32'd3898
; 
32'd157705: dataIn1 = 32'd5661
; 
32'd157706: dataIn1 = 32'd5684
; 
32'd157707: dataIn1 = 32'd5687
; 
32'd157708: dataIn1 = 32'd3896
; 
32'd157709: dataIn1 = 32'd3899
; 
32'd157710: dataIn1 = 32'd5680
; 
32'd157711: dataIn1 = 32'd5688
; 
32'd157712: dataIn1 = 32'd5689
; 
32'd157713: dataIn1 = 32'd5690
; 
32'd157714: dataIn1 = 32'd5691
; 
32'd157715: dataIn1 = 32'd2288
; 
32'd157716: dataIn1 = 32'd3896
; 
32'd157717: dataIn1 = 32'd5682
; 
32'd157718: dataIn1 = 32'd5688
; 
32'd157719: dataIn1 = 32'd5689
; 
32'd157720: dataIn1 = 32'd5690
; 
32'd157721: dataIn1 = 32'd5692
; 
32'd157722: dataIn1 = 32'd2288
; 
32'd157723: dataIn1 = 32'd3866
; 
32'd157724: dataIn1 = 32'd3899
; 
32'd157725: dataIn1 = 32'd5688
; 
32'd157726: dataIn1 = 32'd5689
; 
32'd157727: dataIn1 = 32'd5690
; 
32'd157728: dataIn1 = 32'd5951
; 
32'd157729: dataIn1 = 32'd2302
; 
32'd157730: dataIn1 = 32'd3899
; 
32'd157731: dataIn1 = 32'd5680
; 
32'd157732: dataIn1 = 32'd5688
; 
32'd157733: dataIn1 = 32'd5691
; 
32'd157734: dataIn1 = 32'd5947
; 
32'd157735: dataIn1 = 32'd5950
; 
32'd157736: dataIn1 = 32'd400
; 
32'd157737: dataIn1 = 32'd2288
; 
32'd157738: dataIn1 = 32'd2289
; 
32'd157739: dataIn1 = 32'd5682
; 
32'd157740: dataIn1 = 32'd5689
; 
32'd157741: dataIn1 = 32'd5692
; 
32'd157742: dataIn1 = 32'd3901
; 
32'd157743: dataIn1 = 32'd3902
; 
32'd157744: dataIn1 = 32'd5693
; 
32'd157745: dataIn1 = 32'd5694
; 
32'd157746: dataIn1 = 32'd5695
; 
32'd157747: dataIn1 = 32'd5696
; 
32'd157748: dataIn1 = 32'd5697
; 
32'd157749: dataIn1 = 32'd2304
; 
32'd157750: dataIn1 = 32'd3900
; 
32'd157751: dataIn1 = 32'd3902
; 
32'd157752: dataIn1 = 32'd5693
; 
32'd157753: dataIn1 = 32'd5694
; 
32'd157754: dataIn1 = 32'd5695
; 
32'd157755: dataIn1 = 32'd3900
; 
32'd157756: dataIn1 = 32'd3901
; 
32'd157757: dataIn1 = 32'd5693
; 
32'd157758: dataIn1 = 32'd5694
; 
32'd157759: dataIn1 = 32'd5695
; 
32'd157760: dataIn1 = 32'd5698
; 
32'd157761: dataIn1 = 32'd5699
; 
32'd157762: dataIn1 = 32'd2303
; 
32'd157763: dataIn1 = 32'd3902
; 
32'd157764: dataIn1 = 32'd5693
; 
32'd157765: dataIn1 = 32'd5696
; 
32'd157766: dataIn1 = 32'd5697
; 
32'd157767: dataIn1 = 32'd5707
; 
32'd157768: dataIn1 = 32'd5708
; 
32'd157769: dataIn1 = 32'd2303
; 
32'd157770: dataIn1 = 32'd3901
; 
32'd157771: dataIn1 = 32'd5693
; 
32'd157772: dataIn1 = 32'd5696
; 
32'd157773: dataIn1 = 32'd5697
; 
32'd157774: dataIn1 = 32'd5702
; 
32'd157775: dataIn1 = 32'd5705
; 
32'd157776: dataIn1 = 32'd2305
; 
32'd157777: dataIn1 = 32'd3901
; 
32'd157778: dataIn1 = 32'd5695
; 
32'd157779: dataIn1 = 32'd5698
; 
32'd157780: dataIn1 = 32'd5699
; 
32'd157781: dataIn1 = 32'd5704
; 
32'd157782: dataIn1 = 32'd5706
; 
32'd157783: dataIn1 = 32'd2305
; 
32'd157784: dataIn1 = 32'd3900
; 
32'd157785: dataIn1 = 32'd5695
; 
32'd157786: dataIn1 = 32'd5698
; 
32'd157787: dataIn1 = 32'd5699
; 
32'd157788: dataIn1 = 32'd5700
; 
32'd157789: dataIn1 = 32'd5701
; 
32'd157790: dataIn1 = 32'd2305
; 
32'd157791: dataIn1 = 32'd3903
; 
32'd157792: dataIn1 = 32'd5699
; 
32'd157793: dataIn1 = 32'd5700
; 
32'd157794: dataIn1 = 32'd5701
; 
32'd157795: dataIn1 = 32'd5751
; 
32'd157796: dataIn1 = 32'd5754
; 
32'd157797: dataIn1 = 32'd3900
; 
32'd157798: dataIn1 = 32'd3903
; 
32'd157799: dataIn1 = 32'd3904
; 
32'd157800: dataIn1 = 32'd5699
; 
32'd157801: dataIn1 = 32'd5700
; 
32'd157802: dataIn1 = 32'd5701
; 
32'd157803: dataIn1 = 32'd3901
; 
32'd157804: dataIn1 = 32'd3906
; 
32'd157805: dataIn1 = 32'd5697
; 
32'd157806: dataIn1 = 32'd5702
; 
32'd157807: dataIn1 = 32'd5703
; 
32'd157808: dataIn1 = 32'd5704
; 
32'd157809: dataIn1 = 32'd5705
; 
32'd157810: dataIn1 = 32'd206
; 
32'd157811: dataIn1 = 32'd3905
; 
32'd157812: dataIn1 = 32'd3906
; 
32'd157813: dataIn1 = 32'd5702
; 
32'd157814: dataIn1 = 32'd5703
; 
32'd157815: dataIn1 = 32'd5704
; 
32'd157816: dataIn1 = 32'd3901
; 
32'd157817: dataIn1 = 32'd3905
; 
32'd157818: dataIn1 = 32'd5698
; 
32'd157819: dataIn1 = 32'd5702
; 
32'd157820: dataIn1 = 32'd5703
; 
32'd157821: dataIn1 = 32'd5704
; 
32'd157822: dataIn1 = 32'd5706
; 
32'd157823: dataIn1 = 32'd2303
; 
32'd157824: dataIn1 = 32'd3906
; 
32'd157825: dataIn1 = 32'd5697
; 
32'd157826: dataIn1 = 32'd5702
; 
32'd157827: dataIn1 = 32'd5705
; 
32'd157828: dataIn1 = 32'd5713
; 
32'd157829: dataIn1 = 32'd5725
; 
32'd157830: dataIn1 = 32'd2305
; 
32'd157831: dataIn1 = 32'd3905
; 
32'd157832: dataIn1 = 32'd5698
; 
32'd157833: dataIn1 = 32'd5704
; 
32'd157834: dataIn1 = 32'd5706
; 
32'd157835: dataIn1 = 32'd5750
; 
32'd157836: dataIn1 = 32'd5756
; 
32'd157837: dataIn1 = 32'd3902
; 
32'd157838: dataIn1 = 32'd3907
; 
32'd157839: dataIn1 = 32'd3908
; 
32'd157840: dataIn1 = 32'd5696
; 
32'd157841: dataIn1 = 32'd5707
; 
32'd157842: dataIn1 = 32'd5708
; 
32'd157843: dataIn1 = 32'd2303
; 
32'd157844: dataIn1 = 32'd3908
; 
32'd157845: dataIn1 = 32'd5696
; 
32'd157846: dataIn1 = 32'd5707
; 
32'd157847: dataIn1 = 32'd5708
; 
32'd157848: dataIn1 = 32'd5712
; 
32'd157849: dataIn1 = 32'd5726
; 
32'd157850: dataIn1 = 32'd3910
; 
32'd157851: dataIn1 = 32'd3911
; 
32'd157852: dataIn1 = 32'd5709
; 
32'd157853: dataIn1 = 32'd5710
; 
32'd157854: dataIn1 = 32'd5711
; 
32'd157855: dataIn1 = 32'd5712
; 
32'd157856: dataIn1 = 32'd5713
; 
32'd157857: dataIn1 = 32'd3909
; 
32'd157858: dataIn1 = 32'd3911
; 
32'd157859: dataIn1 = 32'd5709
; 
32'd157860: dataIn1 = 32'd5710
; 
32'd157861: dataIn1 = 32'd5711
; 
32'd157862: dataIn1 = 32'd5714
; 
32'd157863: dataIn1 = 32'd5715
; 
32'd157864: dataIn1 = 32'd3909
; 
32'd157865: dataIn1 = 32'd3910
; 
32'd157866: dataIn1 = 32'd5709
; 
32'd157867: dataIn1 = 32'd5710
; 
32'd157868: dataIn1 = 32'd5711
; 
32'd157869: dataIn1 = 32'd5716
; 
32'd157870: dataIn1 = 32'd5717
; 
32'd157871: dataIn1 = 32'd2303
; 
32'd157872: dataIn1 = 32'd3911
; 
32'd157873: dataIn1 = 32'd5708
; 
32'd157874: dataIn1 = 32'd5709
; 
32'd157875: dataIn1 = 32'd5712
; 
32'd157876: dataIn1 = 32'd5713
; 
32'd157877: dataIn1 = 32'd5726
; 
32'd157878: dataIn1 = 32'd2303
; 
32'd157879: dataIn1 = 32'd3910
; 
32'd157880: dataIn1 = 32'd5705
; 
32'd157881: dataIn1 = 32'd5709
; 
32'd157882: dataIn1 = 32'd5712
; 
32'd157883: dataIn1 = 32'd5713
; 
32'd157884: dataIn1 = 32'd5725
; 
32'd157885: dataIn1 = 32'd2306
; 
32'd157886: dataIn1 = 32'd3911
; 
32'd157887: dataIn1 = 32'd3913
; 
32'd157888: dataIn1 = 32'd5710
; 
32'd157889: dataIn1 = 32'd5714
; 
32'd157890: dataIn1 = 32'd5715
; 
32'd157891: dataIn1 = 32'd2306
; 
32'd157892: dataIn1 = 32'd3909
; 
32'd157893: dataIn1 = 32'd5710
; 
32'd157894: dataIn1 = 32'd5714
; 
32'd157895: dataIn1 = 32'd5715
; 
32'd157896: dataIn1 = 32'd5719
; 
32'd157897: dataIn1 = 32'd5723
; 
32'd157898: dataIn1 = 32'd974
; 
32'd157899: dataIn1 = 32'd2527
; 
32'd157900: dataIn1 = 32'd3910
; 
32'd157901: dataIn1 = 32'd5711
; 
32'd157902: dataIn1 = 32'd5716
; 
32'd157903: dataIn1 = 32'd5717
; 
32'd157904: dataIn1 = 32'd974
; 
32'd157905: dataIn1 = 32'd3909
; 
32'd157906: dataIn1 = 32'd5711
; 
32'd157907: dataIn1 = 32'd5716
; 
32'd157908: dataIn1 = 32'd5717
; 
32'd157909: dataIn1 = 32'd5720
; 
32'd157910: dataIn1 = 32'd5724
; 
32'd157911: dataIn1 = 32'd2525
; 
32'd157912: dataIn1 = 32'd3912
; 
32'd157913: dataIn1 = 32'd5718
; 
32'd157914: dataIn1 = 32'd5719
; 
32'd157915: dataIn1 = 32'd5720
; 
32'd157916: dataIn1 = 32'd5721
; 
32'd157917: dataIn1 = 32'd5722
; 
32'd157918: dataIn1 = 32'd3909
; 
32'd157919: dataIn1 = 32'd3912
; 
32'd157920: dataIn1 = 32'd5715
; 
32'd157921: dataIn1 = 32'd5718
; 
32'd157922: dataIn1 = 32'd5719
; 
32'd157923: dataIn1 = 32'd5720
; 
32'd157924: dataIn1 = 32'd5723
; 
32'd157925: dataIn1 = 32'd2525
; 
32'd157926: dataIn1 = 32'd3909
; 
32'd157927: dataIn1 = 32'd5717
; 
32'd157928: dataIn1 = 32'd5718
; 
32'd157929: dataIn1 = 32'd5719
; 
32'd157930: dataIn1 = 32'd5720
; 
32'd157931: dataIn1 = 32'd5724
; 
32'd157932: dataIn1 = 32'd129
; 
32'd157933: dataIn1 = 32'd3912
; 
32'd157934: dataIn1 = 32'd5718
; 
32'd157935: dataIn1 = 32'd5721
; 
32'd157936: dataIn1 = 32'd5722
; 
32'd157937: dataIn1 = 32'd5936
; 
32'd157938: dataIn1 = 32'd6063
; 
32'd157939: dataIn1 = 32'd129
; 
32'd157940: dataIn1 = 32'd2525
; 
32'd157941: dataIn1 = 32'd2526
; 
32'd157942: dataIn1 = 32'd5718
; 
32'd157943: dataIn1 = 32'd5721
; 
32'd157944: dataIn1 = 32'd5722
; 
32'd157945: dataIn1 = 32'd2306
; 
32'd157946: dataIn1 = 32'd3912
; 
32'd157947: dataIn1 = 32'd5715
; 
32'd157948: dataIn1 = 32'd5719
; 
32'd157949: dataIn1 = 32'd5723
; 
32'd157950: dataIn1 = 32'd6062
; 
32'd157951: dataIn1 = 32'd6064
; 
32'd157952: dataIn1 = 32'd974
; 
32'd157953: dataIn1 = 32'd2523
; 
32'd157954: dataIn1 = 32'd2525
; 
32'd157955: dataIn1 = 32'd5717
; 
32'd157956: dataIn1 = 32'd5720
; 
32'd157957: dataIn1 = 32'd5724
; 
32'd157958: dataIn1 = 32'd2527
; 
32'd157959: dataIn1 = 32'd3906
; 
32'd157960: dataIn1 = 32'd3910
; 
32'd157961: dataIn1 = 32'd5705
; 
32'd157962: dataIn1 = 32'd5713
; 
32'd157963: dataIn1 = 32'd5725
; 
32'd157964: dataIn1 = 32'd3908
; 
32'd157965: dataIn1 = 32'd3911
; 
32'd157966: dataIn1 = 32'd3913
; 
32'd157967: dataIn1 = 32'd5708
; 
32'd157968: dataIn1 = 32'd5712
; 
32'd157969: dataIn1 = 32'd5726
; 
32'd157970: dataIn1 = 32'd3915
; 
32'd157971: dataIn1 = 32'd3916
; 
32'd157972: dataIn1 = 32'd5727
; 
32'd157973: dataIn1 = 32'd5728
; 
32'd157974: dataIn1 = 32'd5729
; 
32'd157975: dataIn1 = 32'd5730
; 
32'd157976: dataIn1 = 32'd5731
; 
32'd157977: dataIn1 = 32'd2304
; 
32'd157978: dataIn1 = 32'd3914
; 
32'd157979: dataIn1 = 32'd3916
; 
32'd157980: dataIn1 = 32'd5727
; 
32'd157981: dataIn1 = 32'd5728
; 
32'd157982: dataIn1 = 32'd5729
; 
32'd157983: dataIn1 = 32'd3914
; 
32'd157984: dataIn1 = 32'd3915
; 
32'd157985: dataIn1 = 32'd5727
; 
32'd157986: dataIn1 = 32'd5728
; 
32'd157987: dataIn1 = 32'd5729
; 
32'd157988: dataIn1 = 32'd5732
; 
32'd157989: dataIn1 = 32'd5733
; 
32'd157990: dataIn1 = 32'd2307
; 
32'd157991: dataIn1 = 32'd3916
; 
32'd157992: dataIn1 = 32'd5727
; 
32'd157993: dataIn1 = 32'd5730
; 
32'd157994: dataIn1 = 32'd5731
; 
32'd157995: dataIn1 = 32'd5743
; 
32'd157996: dataIn1 = 32'd5744
; 
32'd157997: dataIn1 = 32'd2307
; 
32'd157998: dataIn1 = 32'd3915
; 
32'd157999: dataIn1 = 32'd5727
; 
32'd158000: dataIn1 = 32'd5730
; 
32'd158001: dataIn1 = 32'd5731
; 
32'd158002: dataIn1 = 32'd5736
; 
32'd158003: dataIn1 = 32'd5739
; 
32'd158004: dataIn1 = 32'd2308
; 
32'd158005: dataIn1 = 32'd3915
; 
32'd158006: dataIn1 = 32'd5729
; 
32'd158007: dataIn1 = 32'd5732
; 
32'd158008: dataIn1 = 32'd5733
; 
32'd158009: dataIn1 = 32'd5738
; 
32'd158010: dataIn1 = 32'd5742
; 
32'd158011: dataIn1 = 32'd2308
; 
32'd158012: dataIn1 = 32'd3914
; 
32'd158013: dataIn1 = 32'd5729
; 
32'd158014: dataIn1 = 32'd5732
; 
32'd158015: dataIn1 = 32'd5733
; 
32'd158016: dataIn1 = 32'd5734
; 
32'd158017: dataIn1 = 32'd5735
; 
32'd158018: dataIn1 = 32'd2308
; 
32'd158019: dataIn1 = 32'd3917
; 
32'd158020: dataIn1 = 32'd5733
; 
32'd158021: dataIn1 = 32'd5734
; 
32'd158022: dataIn1 = 32'd5735
; 
32'd158023: dataIn1 = 32'd5811
; 
32'd158024: dataIn1 = 32'd5815
; 
32'd158025: dataIn1 = 32'd3904
; 
32'd158026: dataIn1 = 32'd3914
; 
32'd158027: dataIn1 = 32'd3917
; 
32'd158028: dataIn1 = 32'd5733
; 
32'd158029: dataIn1 = 32'd5734
; 
32'd158030: dataIn1 = 32'd5735
; 
32'd158031: dataIn1 = 32'd3915
; 
32'd158032: dataIn1 = 32'd3919
; 
32'd158033: dataIn1 = 32'd5731
; 
32'd158034: dataIn1 = 32'd5736
; 
32'd158035: dataIn1 = 32'd5737
; 
32'd158036: dataIn1 = 32'd5738
; 
32'd158037: dataIn1 = 32'd5739
; 
32'd158038: dataIn1 = 32'd3918
; 
32'd158039: dataIn1 = 32'd3919
; 
32'd158040: dataIn1 = 32'd5736
; 
32'd158041: dataIn1 = 32'd5737
; 
32'd158042: dataIn1 = 32'd5738
; 
32'd158043: dataIn1 = 32'd5740
; 
32'd158044: dataIn1 = 32'd5741
; 
32'd158045: dataIn1 = 32'd3915
; 
32'd158046: dataIn1 = 32'd3918
; 
32'd158047: dataIn1 = 32'd5732
; 
32'd158048: dataIn1 = 32'd5736
; 
32'd158049: dataIn1 = 32'd5737
; 
32'd158050: dataIn1 = 32'd5738
; 
32'd158051: dataIn1 = 32'd5742
; 
32'd158052: dataIn1 = 32'd2307
; 
32'd158053: dataIn1 = 32'd3919
; 
32'd158054: dataIn1 = 32'd5731
; 
32'd158055: dataIn1 = 32'd5736
; 
32'd158056: dataIn1 = 32'd5739
; 
32'd158057: dataIn1 = 32'd6049
; 
32'd158058: dataIn1 = 32'd6054
; 
32'd158059: dataIn1 = 32'd5
; 
32'd158060: dataIn1 = 32'd3919
; 
32'd158061: dataIn1 = 32'd5737
; 
32'd158062: dataIn1 = 32'd5740
; 
32'd158063: dataIn1 = 32'd5741
; 
32'd158064: dataIn1 = 32'd6053
; 
32'd158065: dataIn1 = 32'd6055
; 
32'd158066: dataIn1 = 32'd5
; 
32'd158067: dataIn1 = 32'd3918
; 
32'd158068: dataIn1 = 32'd5737
; 
32'd158069: dataIn1 = 32'd5740
; 
32'd158070: dataIn1 = 32'd5741
; 
32'd158071: dataIn1 = 32'd5824
; 
32'd158072: dataIn1 = 32'd5826
; 
32'd158073: dataIn1 = 32'd2308
; 
32'd158074: dataIn1 = 32'd3918
; 
32'd158075: dataIn1 = 32'd5732
; 
32'd158076: dataIn1 = 32'd5738
; 
32'd158077: dataIn1 = 32'd5742
; 
32'd158078: dataIn1 = 32'd5810
; 
32'd158079: dataIn1 = 32'd5823
; 
32'd158080: dataIn1 = 32'd3907
; 
32'd158081: dataIn1 = 32'd3916
; 
32'd158082: dataIn1 = 32'd3920
; 
32'd158083: dataIn1 = 32'd5730
; 
32'd158084: dataIn1 = 32'd5743
; 
32'd158085: dataIn1 = 32'd5744
; 
32'd158086: dataIn1 = 32'd2307
; 
32'd158087: dataIn1 = 32'd3920
; 
32'd158088: dataIn1 = 32'd5730
; 
32'd158089: dataIn1 = 32'd5743
; 
32'd158090: dataIn1 = 32'd5744
; 
32'd158091: dataIn1 = 32'd6050
; 
32'd158092: dataIn1 = 32'd6696
; 
32'd158093: dataIn1 = 32'd404
; 
32'd158094: dataIn1 = 32'd3922
; 
32'd158095: dataIn1 = 32'd3923
; 
32'd158096: dataIn1 = 32'd5745
; 
32'd158097: dataIn1 = 32'd5746
; 
32'd158098: dataIn1 = 32'd5747
; 
32'd158099: dataIn1 = 32'd3921
; 
32'd158100: dataIn1 = 32'd3923
; 
32'd158101: dataIn1 = 32'd5745
; 
32'd158102: dataIn1 = 32'd5746
; 
32'd158103: dataIn1 = 32'd5747
; 
32'd158104: dataIn1 = 32'd5748
; 
32'd158105: dataIn1 = 32'd5749
; 
32'd158106: dataIn1 = 32'd3921
; 
32'd158107: dataIn1 = 32'd3922
; 
32'd158108: dataIn1 = 32'd5745
; 
32'd158109: dataIn1 = 32'd5746
; 
32'd158110: dataIn1 = 32'd5747
; 
32'd158111: dataIn1 = 32'd5750
; 
32'd158112: dataIn1 = 32'd5751
; 
32'd158113: dataIn1 = 32'd2309
; 
32'd158114: dataIn1 = 32'd3923
; 
32'd158115: dataIn1 = 32'd3925
; 
32'd158116: dataIn1 = 32'd5746
; 
32'd158117: dataIn1 = 32'd5748
; 
32'd158118: dataIn1 = 32'd5749
; 
32'd158119: dataIn1 = 32'd2309
; 
32'd158120: dataIn1 = 32'd3921
; 
32'd158121: dataIn1 = 32'd5746
; 
32'd158122: dataIn1 = 32'd5748
; 
32'd158123: dataIn1 = 32'd5749
; 
32'd158124: dataIn1 = 32'd5753
; 
32'd158125: dataIn1 = 32'd5755
; 
32'd158126: dataIn1 = 32'd2305
; 
32'd158127: dataIn1 = 32'd3922
; 
32'd158128: dataIn1 = 32'd5706
; 
32'd158129: dataIn1 = 32'd5747
; 
32'd158130: dataIn1 = 32'd5750
; 
32'd158131: dataIn1 = 32'd5751
; 
32'd158132: dataIn1 = 32'd5756
; 
32'd158133: dataIn1 = 32'd2305
; 
32'd158134: dataIn1 = 32'd3921
; 
32'd158135: dataIn1 = 32'd5700
; 
32'd158136: dataIn1 = 32'd5747
; 
32'd158137: dataIn1 = 32'd5750
; 
32'd158138: dataIn1 = 32'd5751
; 
32'd158139: dataIn1 = 32'd5754
; 
32'd158140: dataIn1 = 32'd446
; 
32'd158141: dataIn1 = 32'd3903
; 
32'd158142: dataIn1 = 32'd3924
; 
32'd158143: dataIn1 = 32'd5752
; 
32'd158144: dataIn1 = 32'd5753
; 
32'd158145: dataIn1 = 32'd5754
; 
32'd158146: dataIn1 = 32'd3921
; 
32'd158147: dataIn1 = 32'd3924
; 
32'd158148: dataIn1 = 32'd5749
; 
32'd158149: dataIn1 = 32'd5752
; 
32'd158150: dataIn1 = 32'd5753
; 
32'd158151: dataIn1 = 32'd5754
; 
32'd158152: dataIn1 = 32'd5755
; 
32'd158153: dataIn1 = 32'd3903
; 
32'd158154: dataIn1 = 32'd3921
; 
32'd158155: dataIn1 = 32'd5700
; 
32'd158156: dataIn1 = 32'd5751
; 
32'd158157: dataIn1 = 32'd5752
; 
32'd158158: dataIn1 = 32'd5753
; 
32'd158159: dataIn1 = 32'd5754
; 
32'd158160: dataIn1 = 32'd2309
; 
32'd158161: dataIn1 = 32'd3924
; 
32'd158162: dataIn1 = 32'd5749
; 
32'd158163: dataIn1 = 32'd5753
; 
32'd158164: dataIn1 = 32'd5755
; 
32'd158165: dataIn1 = 32'd5802
; 
32'd158166: dataIn1 = 32'd5803
; 
32'd158167: dataIn1 = 32'd2293
; 
32'd158168: dataIn1 = 32'd3905
; 
32'd158169: dataIn1 = 32'd3922
; 
32'd158170: dataIn1 = 32'd5706
; 
32'd158171: dataIn1 = 32'd5750
; 
32'd158172: dataIn1 = 32'd5756
; 
32'd158173: dataIn1 = 32'd3935
; 
32'd158174: dataIn1 = 32'd3936
; 
32'd158175: dataIn1 = 32'd5757
; 
32'd158176: dataIn1 = 32'd5758
; 
32'd158177: dataIn1 = 32'd5759
; 
32'd158178: dataIn1 = 32'd5760
; 
32'd158179: dataIn1 = 32'd5761
; 
32'd158180: dataIn1 = 32'd2313
; 
32'd158181: dataIn1 = 32'd3934
; 
32'd158182: dataIn1 = 32'd3936
; 
32'd158183: dataIn1 = 32'd5757
; 
32'd158184: dataIn1 = 32'd5758
; 
32'd158185: dataIn1 = 32'd5759
; 
32'd158186: dataIn1 = 32'd3934
; 
32'd158187: dataIn1 = 32'd3935
; 
32'd158188: dataIn1 = 32'd5757
; 
32'd158189: dataIn1 = 32'd5758
; 
32'd158190: dataIn1 = 32'd5759
; 
32'd158191: dataIn1 = 32'd5762
; 
32'd158192: dataIn1 = 32'd5763
; 
32'd158193: dataIn1 = 32'd2312
; 
32'd158194: dataIn1 = 32'd3936
; 
32'd158195: dataIn1 = 32'd5757
; 
32'd158196: dataIn1 = 32'd5760
; 
32'd158197: dataIn1 = 32'd5761
; 
32'd158198: dataIn1 = 32'd5773
; 
32'd158199: dataIn1 = 32'd5774
; 
32'd158200: dataIn1 = 32'd2312
; 
32'd158201: dataIn1 = 32'd3935
; 
32'd158202: dataIn1 = 32'd5757
; 
32'd158203: dataIn1 = 32'd5760
; 
32'd158204: dataIn1 = 32'd5761
; 
32'd158205: dataIn1 = 32'd5766
; 
32'd158206: dataIn1 = 32'd5769
; 
32'd158207: dataIn1 = 32'd2314
; 
32'd158208: dataIn1 = 32'd3935
; 
32'd158209: dataIn1 = 32'd5759
; 
32'd158210: dataIn1 = 32'd5762
; 
32'd158211: dataIn1 = 32'd5763
; 
32'd158212: dataIn1 = 32'd5768
; 
32'd158213: dataIn1 = 32'd5772
; 
32'd158214: dataIn1 = 32'd2314
; 
32'd158215: dataIn1 = 32'd3934
; 
32'd158216: dataIn1 = 32'd5759
; 
32'd158217: dataIn1 = 32'd5762
; 
32'd158218: dataIn1 = 32'd5763
; 
32'd158219: dataIn1 = 32'd5764
; 
32'd158220: dataIn1 = 32'd5765
; 
32'd158221: dataIn1 = 32'd2314
; 
32'd158222: dataIn1 = 32'd3937
; 
32'd158223: dataIn1 = 32'd5763
; 
32'd158224: dataIn1 = 32'd5764
; 
32'd158225: dataIn1 = 32'd5765
; 
32'd158226: dataIn1 = 32'd5813
; 
32'd158227: dataIn1 = 32'd5816
; 
32'd158228: dataIn1 = 32'd3934
; 
32'd158229: dataIn1 = 32'd3937
; 
32'd158230: dataIn1 = 32'd3938
; 
32'd158231: dataIn1 = 32'd5763
; 
32'd158232: dataIn1 = 32'd5764
; 
32'd158233: dataIn1 = 32'd5765
; 
32'd158234: dataIn1 = 32'd3935
; 
32'd158235: dataIn1 = 32'd3940
; 
32'd158236: dataIn1 = 32'd5761
; 
32'd158237: dataIn1 = 32'd5766
; 
32'd158238: dataIn1 = 32'd5767
; 
32'd158239: dataIn1 = 32'd5768
; 
32'd158240: dataIn1 = 32'd5769
; 
32'd158241: dataIn1 = 32'd3939
; 
32'd158242: dataIn1 = 32'd3940
; 
32'd158243: dataIn1 = 32'd5766
; 
32'd158244: dataIn1 = 32'd5767
; 
32'd158245: dataIn1 = 32'd5768
; 
32'd158246: dataIn1 = 32'd5770
; 
32'd158247: dataIn1 = 32'd5771
; 
32'd158248: dataIn1 = 32'd3935
; 
32'd158249: dataIn1 = 32'd3939
; 
32'd158250: dataIn1 = 32'd5762
; 
32'd158251: dataIn1 = 32'd5766
; 
32'd158252: dataIn1 = 32'd5767
; 
32'd158253: dataIn1 = 32'd5768
; 
32'd158254: dataIn1 = 32'd5772
; 
32'd158255: dataIn1 = 32'd2312
; 
32'd158256: dataIn1 = 32'd3940
; 
32'd158257: dataIn1 = 32'd5761
; 
32'd158258: dataIn1 = 32'd5766
; 
32'd158259: dataIn1 = 32'd5769
; 
32'd158260: dataIn1 = 32'd5779
; 
32'd158261: dataIn1 = 32'd5790
; 
32'd158262: dataIn1 = 32'd449
; 
32'd158263: dataIn1 = 32'd3940
; 
32'd158264: dataIn1 = 32'd5767
; 
32'd158265: dataIn1 = 32'd5770
; 
32'd158266: dataIn1 = 32'd5771
; 
32'd158267: dataIn1 = 32'd5791
; 
32'd158268: dataIn1 = 32'd5793
; 
32'd158269: dataIn1 = 32'd449
; 
32'd158270: dataIn1 = 32'd3939
; 
32'd158271: dataIn1 = 32'd5767
; 
32'd158272: dataIn1 = 32'd5770
; 
32'd158273: dataIn1 = 32'd5771
; 
32'd158274: dataIn1 = 32'd5818
; 
32'd158275: dataIn1 = 32'd5821
; 
32'd158276: dataIn1 = 32'd2314
; 
32'd158277: dataIn1 = 32'd3939
; 
32'd158278: dataIn1 = 32'd5762
; 
32'd158279: dataIn1 = 32'd5768
; 
32'd158280: dataIn1 = 32'd5772
; 
32'd158281: dataIn1 = 32'd5812
; 
32'd158282: dataIn1 = 32'd5819
; 
32'd158283: dataIn1 = 32'd3936
; 
32'd158284: dataIn1 = 32'd3941
; 
32'd158285: dataIn1 = 32'd3942
; 
32'd158286: dataIn1 = 32'd5760
; 
32'd158287: dataIn1 = 32'd5773
; 
32'd158288: dataIn1 = 32'd5774
; 
32'd158289: dataIn1 = 32'd2312
; 
32'd158290: dataIn1 = 32'd3942
; 
32'd158291: dataIn1 = 32'd5760
; 
32'd158292: dataIn1 = 32'd5773
; 
32'd158293: dataIn1 = 32'd5774
; 
32'd158294: dataIn1 = 32'd5778
; 
32'd158295: dataIn1 = 32'd5795
; 
32'd158296: dataIn1 = 32'd3944
; 
32'd158297: dataIn1 = 32'd3945
; 
32'd158298: dataIn1 = 32'd5775
; 
32'd158299: dataIn1 = 32'd5776
; 
32'd158300: dataIn1 = 32'd5777
; 
32'd158301: dataIn1 = 32'd5778
; 
32'd158302: dataIn1 = 32'd5779
; 
32'd158303: dataIn1 = 32'd3943
; 
32'd158304: dataIn1 = 32'd3945
; 
32'd158305: dataIn1 = 32'd5775
; 
32'd158306: dataIn1 = 32'd5776
; 
32'd158307: dataIn1 = 32'd5777
; 
32'd158308: dataIn1 = 32'd5780
; 
32'd158309: dataIn1 = 32'd5781
; 
32'd158310: dataIn1 = 32'd3943
; 
32'd158311: dataIn1 = 32'd3944
; 
32'd158312: dataIn1 = 32'd5775
; 
32'd158313: dataIn1 = 32'd5776
; 
32'd158314: dataIn1 = 32'd5777
; 
32'd158315: dataIn1 = 32'd5782
; 
32'd158316: dataIn1 = 32'd5783
; 
32'd158317: dataIn1 = 32'd2312
; 
32'd158318: dataIn1 = 32'd3945
; 
32'd158319: dataIn1 = 32'd5774
; 
32'd158320: dataIn1 = 32'd5775
; 
32'd158321: dataIn1 = 32'd5778
; 
32'd158322: dataIn1 = 32'd5779
; 
32'd158323: dataIn1 = 32'd5795
; 
32'd158324: dataIn1 = 32'd2312
; 
32'd158325: dataIn1 = 32'd3944
; 
32'd158326: dataIn1 = 32'd5769
; 
32'd158327: dataIn1 = 32'd5775
; 
32'd158328: dataIn1 = 32'd5778
; 
32'd158329: dataIn1 = 32'd5779
; 
32'd158330: dataIn1 = 32'd5790
; 
32'd158331: dataIn1 = 32'd2299
; 
32'd158332: dataIn1 = 32'd3886
; 
32'd158333: dataIn1 = 32'd3945
; 
32'd158334: dataIn1 = 32'd5776
; 
32'd158335: dataIn1 = 32'd5780
; 
32'd158336: dataIn1 = 32'd5781
; 
32'd158337: dataIn1 = 32'd2299
; 
32'd158338: dataIn1 = 32'd3943
; 
32'd158339: dataIn1 = 32'd5776
; 
32'd158340: dataIn1 = 32'd5780
; 
32'd158341: dataIn1 = 32'd5781
; 
32'd158342: dataIn1 = 32'd5785
; 
32'd158343: dataIn1 = 32'd5788
; 
32'd158344: dataIn1 = 32'd2315
; 
32'd158345: dataIn1 = 32'd3944
; 
32'd158346: dataIn1 = 32'd5777
; 
32'd158347: dataIn1 = 32'd5782
; 
32'd158348: dataIn1 = 32'd5783
; 
32'd158349: dataIn1 = 32'd5792
; 
32'd158350: dataIn1 = 32'd5794
; 
32'd158351: dataIn1 = 32'd2315
; 
32'd158352: dataIn1 = 32'd3943
; 
32'd158353: dataIn1 = 32'd5777
; 
32'd158354: dataIn1 = 32'd5782
; 
32'd158355: dataIn1 = 32'd5783
; 
32'd158356: dataIn1 = 32'd5786
; 
32'd158357: dataIn1 = 32'd5789
; 
32'd158358: dataIn1 = 32'd3884
; 
32'd158359: dataIn1 = 32'd3946
; 
32'd158360: dataIn1 = 32'd5666
; 
32'd158361: dataIn1 = 32'd5784
; 
32'd158362: dataIn1 = 32'd5785
; 
32'd158363: dataIn1 = 32'd5786
; 
32'd158364: dataIn1 = 32'd5787
; 
32'd158365: dataIn1 = 32'd3884
; 
32'd158366: dataIn1 = 32'd3943
; 
32'd158367: dataIn1 = 32'd5781
; 
32'd158368: dataIn1 = 32'd5784
; 
32'd158369: dataIn1 = 32'd5785
; 
32'd158370: dataIn1 = 32'd5786
; 
32'd158371: dataIn1 = 32'd5788
; 
32'd158372: dataIn1 = 32'd3943
; 
32'd158373: dataIn1 = 32'd3946
; 
32'd158374: dataIn1 = 32'd5783
; 
32'd158375: dataIn1 = 32'd5784
; 
32'd158376: dataIn1 = 32'd5785
; 
32'd158377: dataIn1 = 32'd5786
; 
32'd158378: dataIn1 = 32'd5789
; 
32'd158379: dataIn1 = 32'd127
; 
32'd158380: dataIn1 = 32'd3946
; 
32'd158381: dataIn1 = 32'd5666
; 
32'd158382: dataIn1 = 32'd5784
; 
32'd158383: dataIn1 = 32'd5787
; 
32'd158384: dataIn1 = 32'd6892
; 
32'd158385: dataIn1 = 32'd7030
; 
32'd158386: dataIn1 = 32'd2299
; 
32'd158387: dataIn1 = 32'd3880
; 
32'd158388: dataIn1 = 32'd3884
; 
32'd158389: dataIn1 = 32'd5781
; 
32'd158390: dataIn1 = 32'd5785
; 
32'd158391: dataIn1 = 32'd5788
; 
32'd158392: dataIn1 = 32'd2315
; 
32'd158393: dataIn1 = 32'd3946
; 
32'd158394: dataIn1 = 32'd5783
; 
32'd158395: dataIn1 = 32'd5786
; 
32'd158396: dataIn1 = 32'd5789
; 
32'd158397: dataIn1 = 32'd7024
; 
32'd158398: dataIn1 = 32'd7031
; 
32'd158399: dataIn1 = 32'd3940
; 
32'd158400: dataIn1 = 32'd3944
; 
32'd158401: dataIn1 = 32'd5769
; 
32'd158402: dataIn1 = 32'd5779
; 
32'd158403: dataIn1 = 32'd5790
; 
32'd158404: dataIn1 = 32'd5791
; 
32'd158405: dataIn1 = 32'd5792
; 
32'd158406: dataIn1 = 32'd3940
; 
32'd158407: dataIn1 = 32'd3947
; 
32'd158408: dataIn1 = 32'd5770
; 
32'd158409: dataIn1 = 32'd5790
; 
32'd158410: dataIn1 = 32'd5791
; 
32'd158411: dataIn1 = 32'd5792
; 
32'd158412: dataIn1 = 32'd5793
; 
32'd158413: dataIn1 = 32'd3944
; 
32'd158414: dataIn1 = 32'd3947
; 
32'd158415: dataIn1 = 32'd5782
; 
32'd158416: dataIn1 = 32'd5790
; 
32'd158417: dataIn1 = 32'd5791
; 
32'd158418: dataIn1 = 32'd5792
; 
32'd158419: dataIn1 = 32'd5794
; 
32'd158420: dataIn1 = 32'd449
; 
32'd158421: dataIn1 = 32'd3947
; 
32'd158422: dataIn1 = 32'd5770
; 
32'd158423: dataIn1 = 32'd5791
; 
32'd158424: dataIn1 = 32'd5793
; 
32'd158425: dataIn1 = 32'd7001
; 
32'd158426: dataIn1 = 32'd7026
; 
32'd158427: dataIn1 = 32'd2315
; 
32'd158428: dataIn1 = 32'd3947
; 
32'd158429: dataIn1 = 32'd5782
; 
32'd158430: dataIn1 = 32'd5792
; 
32'd158431: dataIn1 = 32'd5794
; 
32'd158432: dataIn1 = 32'd7025
; 
32'd158433: dataIn1 = 32'd7028
; 
32'd158434: dataIn1 = 32'd3886
; 
32'd158435: dataIn1 = 32'd3942
; 
32'd158436: dataIn1 = 32'd3945
; 
32'd158437: dataIn1 = 32'd5774
; 
32'd158438: dataIn1 = 32'd5778
; 
32'd158439: dataIn1 = 32'd5795
; 
32'd158440: dataIn1 = 32'd3949
; 
32'd158441: dataIn1 = 32'd3950
; 
32'd158442: dataIn1 = 32'd5796
; 
32'd158443: dataIn1 = 32'd5797
; 
32'd158444: dataIn1 = 32'd5798
; 
32'd158445: dataIn1 = 32'd5799
; 
32'd158446: dataIn1 = 32'd5800
; 
32'd158447: dataIn1 = 32'd2313
; 
32'd158448: dataIn1 = 32'd3948
; 
32'd158449: dataIn1 = 32'd3950
; 
32'd158450: dataIn1 = 32'd5796
; 
32'd158451: dataIn1 = 32'd5797
; 
32'd158452: dataIn1 = 32'd5798
; 
32'd158453: dataIn1 = 32'd3948
; 
32'd158454: dataIn1 = 32'd3949
; 
32'd158455: dataIn1 = 32'd5796
; 
32'd158456: dataIn1 = 32'd5797
; 
32'd158457: dataIn1 = 32'd5798
; 
32'd158458: dataIn1 = 32'd5801
; 
32'd158459: dataIn1 = 32'd5802
; 
32'd158460: dataIn1 = 32'd2301
; 
32'd158461: dataIn1 = 32'd3950
; 
32'd158462: dataIn1 = 32'd5676
; 
32'd158463: dataIn1 = 32'd5796
; 
32'd158464: dataIn1 = 32'd5799
; 
32'd158465: dataIn1 = 32'd5800
; 
32'd158466: dataIn1 = 32'd5804
; 
32'd158467: dataIn1 = 32'd2301
; 
32'd158468: dataIn1 = 32'd3892
; 
32'd158469: dataIn1 = 32'd3949
; 
32'd158470: dataIn1 = 32'd5796
; 
32'd158471: dataIn1 = 32'd5799
; 
32'd158472: dataIn1 = 32'd5800
; 
32'd158473: dataIn1 = 32'd2309
; 
32'd158474: dataIn1 = 32'd3925
; 
32'd158475: dataIn1 = 32'd3949
; 
32'd158476: dataIn1 = 32'd5798
; 
32'd158477: dataIn1 = 32'd5801
; 
32'd158478: dataIn1 = 32'd5802
; 
32'd158479: dataIn1 = 32'd2309
; 
32'd158480: dataIn1 = 32'd3948
; 
32'd158481: dataIn1 = 32'd5755
; 
32'd158482: dataIn1 = 32'd5798
; 
32'd158483: dataIn1 = 32'd5801
; 
32'd158484: dataIn1 = 32'd5802
; 
32'd158485: dataIn1 = 32'd5803
; 
32'd158486: dataIn1 = 32'd3924
; 
32'd158487: dataIn1 = 32'd3938
; 
32'd158488: dataIn1 = 32'd3948
; 
32'd158489: dataIn1 = 32'd5755
; 
32'd158490: dataIn1 = 32'd5802
; 
32'd158491: dataIn1 = 32'd5803
; 
32'd158492: dataIn1 = 32'd3893
; 
32'd158493: dataIn1 = 32'd3941
; 
32'd158494: dataIn1 = 32'd3950
; 
32'd158495: dataIn1 = 32'd5676
; 
32'd158496: dataIn1 = 32'd5799
; 
32'd158497: dataIn1 = 32'd5804
; 
32'd158498: dataIn1 = 32'd3952
; 
32'd158499: dataIn1 = 32'd3953
; 
32'd158500: dataIn1 = 32'd5805
; 
32'd158501: dataIn1 = 32'd5806
; 
32'd158502: dataIn1 = 32'd5807
; 
32'd158503: dataIn1 = 32'd5808
; 
32'd158504: dataIn1 = 32'd5809
; 
32'd158505: dataIn1 = 32'd3951
; 
32'd158506: dataIn1 = 32'd3953
; 
32'd158507: dataIn1 = 32'd5805
; 
32'd158508: dataIn1 = 32'd5806
; 
32'd158509: dataIn1 = 32'd5807
; 
32'd158510: dataIn1 = 32'd5810
; 
32'd158511: dataIn1 = 32'd5811
; 
32'd158512: dataIn1 = 32'd3951
; 
32'd158513: dataIn1 = 32'd3952
; 
32'd158514: dataIn1 = 32'd5805
; 
32'd158515: dataIn1 = 32'd5806
; 
32'd158516: dataIn1 = 32'd5807
; 
32'd158517: dataIn1 = 32'd5812
; 
32'd158518: dataIn1 = 32'd5813
; 
32'd158519: dataIn1 = 32'd2316
; 
32'd158520: dataIn1 = 32'd3953
; 
32'd158521: dataIn1 = 32'd5805
; 
32'd158522: dataIn1 = 32'd5808
; 
32'd158523: dataIn1 = 32'd5809
; 
32'd158524: dataIn1 = 32'd5822
; 
32'd158525: dataIn1 = 32'd5825
; 
32'd158526: dataIn1 = 32'd2316
; 
32'd158527: dataIn1 = 32'd3952
; 
32'd158528: dataIn1 = 32'd5805
; 
32'd158529: dataIn1 = 32'd5808
; 
32'd158530: dataIn1 = 32'd5809
; 
32'd158531: dataIn1 = 32'd5817
; 
32'd158532: dataIn1 = 32'd5820
; 
32'd158533: dataIn1 = 32'd2308
; 
32'd158534: dataIn1 = 32'd3953
; 
32'd158535: dataIn1 = 32'd5742
; 
32'd158536: dataIn1 = 32'd5806
; 
32'd158537: dataIn1 = 32'd5810
; 
32'd158538: dataIn1 = 32'd5811
; 
32'd158539: dataIn1 = 32'd5823
; 
32'd158540: dataIn1 = 32'd2308
; 
32'd158541: dataIn1 = 32'd3951
; 
32'd158542: dataIn1 = 32'd5734
; 
32'd158543: dataIn1 = 32'd5806
; 
32'd158544: dataIn1 = 32'd5810
; 
32'd158545: dataIn1 = 32'd5811
; 
32'd158546: dataIn1 = 32'd5815
; 
32'd158547: dataIn1 = 32'd2314
; 
32'd158548: dataIn1 = 32'd3952
; 
32'd158549: dataIn1 = 32'd5772
; 
32'd158550: dataIn1 = 32'd5807
; 
32'd158551: dataIn1 = 32'd5812
; 
32'd158552: dataIn1 = 32'd5813
; 
32'd158553: dataIn1 = 32'd5819
; 
32'd158554: dataIn1 = 32'd2314
; 
32'd158555: dataIn1 = 32'd3951
; 
32'd158556: dataIn1 = 32'd5764
; 
32'd158557: dataIn1 = 32'd5807
; 
32'd158558: dataIn1 = 32'd5812
; 
32'd158559: dataIn1 = 32'd5813
; 
32'd158560: dataIn1 = 32'd5816
; 
32'd158561: dataIn1 = 32'd446
; 
32'd158562: dataIn1 = 32'd3917
; 
32'd158563: dataIn1 = 32'd3937
; 
32'd158564: dataIn1 = 32'd5814
; 
32'd158565: dataIn1 = 32'd5815
; 
32'd158566: dataIn1 = 32'd5816
; 
32'd158567: dataIn1 = 32'd3917
; 
32'd158568: dataIn1 = 32'd3951
; 
32'd158569: dataIn1 = 32'd5734
; 
32'd158570: dataIn1 = 32'd5811
; 
32'd158571: dataIn1 = 32'd5814
; 
32'd158572: dataIn1 = 32'd5815
; 
32'd158573: dataIn1 = 32'd5816
; 
32'd158574: dataIn1 = 32'd3937
; 
32'd158575: dataIn1 = 32'd3951
; 
32'd158576: dataIn1 = 32'd5764
; 
32'd158577: dataIn1 = 32'd5813
; 
32'd158578: dataIn1 = 32'd5814
; 
32'd158579: dataIn1 = 32'd5815
; 
32'd158580: dataIn1 = 32'd5816
; 
32'd158581: dataIn1 = 32'd3952
; 
32'd158582: dataIn1 = 32'd3954
; 
32'd158583: dataIn1 = 32'd5809
; 
32'd158584: dataIn1 = 32'd5817
; 
32'd158585: dataIn1 = 32'd5818
; 
32'd158586: dataIn1 = 32'd5819
; 
32'd158587: dataIn1 = 32'd5820
; 
32'd158588: dataIn1 = 32'd3939
; 
32'd158589: dataIn1 = 32'd3954
; 
32'd158590: dataIn1 = 32'd5771
; 
32'd158591: dataIn1 = 32'd5817
; 
32'd158592: dataIn1 = 32'd5818
; 
32'd158593: dataIn1 = 32'd5819
; 
32'd158594: dataIn1 = 32'd5821
; 
32'd158595: dataIn1 = 32'd3939
; 
32'd158596: dataIn1 = 32'd3952
; 
32'd158597: dataIn1 = 32'd5772
; 
32'd158598: dataIn1 = 32'd5812
; 
32'd158599: dataIn1 = 32'd5817
; 
32'd158600: dataIn1 = 32'd5818
; 
32'd158601: dataIn1 = 32'd5819
; 
32'd158602: dataIn1 = 32'd2316
; 
32'd158603: dataIn1 = 32'd3954
; 
32'd158604: dataIn1 = 32'd5809
; 
32'd158605: dataIn1 = 32'd5817
; 
32'd158606: dataIn1 = 32'd5820
; 
32'd158607: dataIn1 = 32'd7041
; 
32'd158608: dataIn1 = 32'd7045
; 
32'd158609: dataIn1 = 32'd449
; 
32'd158610: dataIn1 = 32'd3954
; 
32'd158611: dataIn1 = 32'd5771
; 
32'd158612: dataIn1 = 32'd5818
; 
32'd158613: dataIn1 = 32'd5821
; 
32'd158614: dataIn1 = 32'd7002
; 
32'd158615: dataIn1 = 32'd7044
; 
32'd158616: dataIn1 = 32'd3953
; 
32'd158617: dataIn1 = 32'd3955
; 
32'd158618: dataIn1 = 32'd5808
; 
32'd158619: dataIn1 = 32'd5822
; 
32'd158620: dataIn1 = 32'd5823
; 
32'd158621: dataIn1 = 32'd5824
; 
32'd158622: dataIn1 = 32'd5825
; 
32'd158623: dataIn1 = 32'd3918
; 
32'd158624: dataIn1 = 32'd3953
; 
32'd158625: dataIn1 = 32'd5742
; 
32'd158626: dataIn1 = 32'd5810
; 
32'd158627: dataIn1 = 32'd5822
; 
32'd158628: dataIn1 = 32'd5823
; 
32'd158629: dataIn1 = 32'd5824
; 
32'd158630: dataIn1 = 32'd3918
; 
32'd158631: dataIn1 = 32'd3955
; 
32'd158632: dataIn1 = 32'd5741
; 
32'd158633: dataIn1 = 32'd5822
; 
32'd158634: dataIn1 = 32'd5823
; 
32'd158635: dataIn1 = 32'd5824
; 
32'd158636: dataIn1 = 32'd5826
; 
32'd158637: dataIn1 = 32'd2316
; 
32'd158638: dataIn1 = 32'd3955
; 
32'd158639: dataIn1 = 32'd5808
; 
32'd158640: dataIn1 = 32'd5822
; 
32'd158641: dataIn1 = 32'd5825
; 
32'd158642: dataIn1 = 32'd7040
; 
32'd158643: dataIn1 = 32'd7052
; 
32'd158644: dataIn1 = 32'd5
; 
32'd158645: dataIn1 = 32'd3955
; 
32'd158646: dataIn1 = 32'd5741
; 
32'd158647: dataIn1 = 32'd5824
; 
32'd158648: dataIn1 = 32'd5826
; 
32'd158649: dataIn1 = 32'd7053
; 
32'd158650: dataIn1 = 32'd8925
; 
32'd158651: dataIn1 = 32'd5827
; 
32'd158652: dataIn1 = 32'd6852
; 
32'd158653: dataIn1 = 32'd6853
; 
32'd158654: dataIn1 = 32'd6857
; 
32'd158655: dataIn1 = 32'd6859
; 
32'd158656: dataIn1 = 32'd6861
; 
32'd158657: dataIn1 = 32'd6862
; 
32'd158658: dataIn1 = 32'd5828
; 
32'd158659: dataIn1 = 32'd6851
; 
32'd158660: dataIn1 = 32'd6853
; 
32'd158661: dataIn1 = 32'd6855
; 
32'd158662: dataIn1 = 32'd6858
; 
32'd158663: dataIn1 = 32'd9270
; 
32'd158664: dataIn1 = 32'd9271
; 
32'd158665: dataIn1 = 32'd5829
; 
32'd158666: dataIn1 = 32'd6851
; 
32'd158667: dataIn1 = 32'd6852
; 
32'd158668: dataIn1 = 32'd6854
; 
32'd158669: dataIn1 = 32'd6856
; 
32'd158670: dataIn1 = 32'd6867
; 
32'd158671: dataIn1 = 32'd6868
; 
32'd158672: dataIn1 = 32'd5830
; 
32'd158673: dataIn1 = 32'd6860
; 
32'd158674: dataIn1 = 32'd6862
; 
32'd158675: dataIn1 = 32'd6864
; 
32'd158676: dataIn1 = 32'd6866
; 
32'd158677: dataIn1 = 32'd6900
; 
32'd158678: dataIn1 = 32'd6902
; 
32'd158679: dataIn1 = 32'd5831
; 
32'd158680: dataIn1 = 32'd6860
; 
32'd158681: dataIn1 = 32'd6861
; 
32'd158682: dataIn1 = 32'd6863
; 
32'd158683: dataIn1 = 32'd6865
; 
32'd158684: dataIn1 = 32'd6883
; 
32'd158685: dataIn1 = 32'd6884
; 
32'd158686: dataIn1 = 32'd5832
; 
32'd158687: dataIn1 = 32'd6868
; 
32'd158688: dataIn1 = 32'd6869
; 
32'd158689: dataIn1 = 32'd6871
; 
32'd158690: dataIn1 = 32'd6873
; 
32'd158691: dataIn1 = 32'd6896
; 
32'd158692: dataIn1 = 32'd6897
; 
32'd158693: dataIn1 = 32'd5833
; 
32'd158694: dataIn1 = 32'd5834
; 
32'd158695: dataIn1 = 32'd5835
; 
32'd158696: dataIn1 = 32'd6867
; 
32'd158697: dataIn1 = 32'd6869
; 
32'd158698: dataIn1 = 32'd6870
; 
32'd158699: dataIn1 = 32'd6872
; 
32'd158700: dataIn1 = 32'd2321
; 
32'd158701: dataIn1 = 32'd3966
; 
32'd158702: dataIn1 = 32'd5833
; 
32'd158703: dataIn1 = 32'd5834
; 
32'd158704: dataIn1 = 32'd5835
; 
32'd158705: dataIn1 = 32'd5879
; 
32'd158706: dataIn1 = 32'd5880
; 
32'd158707: dataIn1 = 32'd6872
; 
32'd158708: dataIn1 = 32'd7015
; 
32'd158709: dataIn1 = 32'd3963
; 
32'd158710: dataIn1 = 32'd3966
; 
32'd158711: dataIn1 = 32'd3967
; 
32'd158712: dataIn1 = 32'd5833
; 
32'd158713: dataIn1 = 32'd5834
; 
32'd158714: dataIn1 = 32'd5835
; 
32'd158715: dataIn1 = 32'd6870
; 
32'd158716: dataIn1 = 32'd5836
; 
32'd158717: dataIn1 = 32'd6875
; 
32'd158718: dataIn1 = 32'd6876
; 
32'd158719: dataIn1 = 32'd6880
; 
32'd158720: dataIn1 = 32'd6882
; 
32'd158721: dataIn1 = 32'd6884
; 
32'd158722: dataIn1 = 32'd6885
; 
32'd158723: dataIn1 = 32'd5837
; 
32'd158724: dataIn1 = 32'd6874
; 
32'd158725: dataIn1 = 32'd6876
; 
32'd158726: dataIn1 = 32'd6878
; 
32'd158727: dataIn1 = 32'd6881
; 
32'd158728: dataIn1 = 32'd6888
; 
32'd158729: dataIn1 = 32'd6890
; 
32'd158730: dataIn1 = 32'd5838
; 
32'd158731: dataIn1 = 32'd6874
; 
32'd158732: dataIn1 = 32'd6875
; 
32'd158733: dataIn1 = 32'd6877
; 
32'd158734: dataIn1 = 32'd6879
; 
32'd158735: dataIn1 = 32'd6895
; 
32'd158736: dataIn1 = 32'd6896
; 
32'd158737: dataIn1 = 32'd5839
; 
32'd158738: dataIn1 = 32'd6883
; 
32'd158739: dataIn1 = 32'd6885
; 
32'd158740: dataIn1 = 32'd6886
; 
32'd158741: dataIn1 = 32'd6887
; 
32'd158742: dataIn1 = 32'd6961
; 
32'd158743: dataIn1 = 32'd6963
; 
32'd158744: dataIn1 = 32'd5840
; 
32'd158745: dataIn1 = 32'd6889
; 
32'd158746: dataIn1 = 32'd6890
; 
32'd158747: dataIn1 = 32'd6893
; 
32'd158748: dataIn1 = 32'd6894
; 
32'd158749: dataIn1 = 32'd6965
; 
32'd158750: dataIn1 = 32'd6966
; 
32'd158751: dataIn1 = 32'd5841
; 
32'd158752: dataIn1 = 32'd6888
; 
32'd158753: dataIn1 = 32'd6889
; 
32'd158754: dataIn1 = 32'd6891
; 
32'd158755: dataIn1 = 32'd6892
; 
32'd158756: dataIn1 = 32'd7029
; 
32'd158757: dataIn1 = 32'd7030
; 
32'd158758: dataIn1 = 32'd5842
; 
32'd158759: dataIn1 = 32'd6895
; 
32'd158760: dataIn1 = 32'd6897
; 
32'd158761: dataIn1 = 32'd6898
; 
32'd158762: dataIn1 = 32'd6899
; 
32'd158763: dataIn1 = 32'd7032
; 
32'd158764: dataIn1 = 32'd7034
; 
32'd158765: dataIn1 = 32'd5843
; 
32'd158766: dataIn1 = 32'd5844
; 
32'd158767: dataIn1 = 32'd5845
; 
32'd158768: dataIn1 = 32'd6901
; 
32'd158769: dataIn1 = 32'd6902
; 
32'd158770: dataIn1 = 32'd6905
; 
32'd158771: dataIn1 = 32'd6906
; 
32'd158772: dataIn1 = 32'd3965
; 
32'd158773: dataIn1 = 32'd3970
; 
32'd158774: dataIn1 = 32'd5843
; 
32'd158775: dataIn1 = 32'd5844
; 
32'd158776: dataIn1 = 32'd5845
; 
32'd158777: dataIn1 = 32'd6906
; 
32'd158778: dataIn1 = 32'd9270
; 
32'd158779: dataIn1 = 32'd9319
; 
32'd158780: dataIn1 = 32'd3970
; 
32'd158781: dataIn1 = 32'd3971
; 
32'd158782: dataIn1 = 32'd5843
; 
32'd158783: dataIn1 = 32'd5844
; 
32'd158784: dataIn1 = 32'd5845
; 
32'd158785: dataIn1 = 32'd5847
; 
32'd158786: dataIn1 = 32'd5848
; 
32'd158787: dataIn1 = 32'd6905
; 
32'd158788: dataIn1 = 32'd5846
; 
32'd158789: dataIn1 = 32'd6900
; 
32'd158790: dataIn1 = 32'd6901
; 
32'd158791: dataIn1 = 32'd6903
; 
32'd158792: dataIn1 = 32'd6904
; 
32'd158793: dataIn1 = 32'd6981
; 
32'd158794: dataIn1 = 32'd6982
; 
32'd158795: dataIn1 = 32'd452
; 
32'd158796: dataIn1 = 32'd3971
; 
32'd158797: dataIn1 = 32'd5845
; 
32'd158798: dataIn1 = 32'd5847
; 
32'd158799: dataIn1 = 32'd5848
; 
32'd158800: dataIn1 = 32'd5868
; 
32'd158801: dataIn1 = 32'd5870
; 
32'd158802: dataIn1 = 32'd6977
; 
32'd158803: dataIn1 = 32'd452
; 
32'd158804: dataIn1 = 32'd3970
; 
32'd158805: dataIn1 = 32'd3980
; 
32'd158806: dataIn1 = 32'd5845
; 
32'd158807: dataIn1 = 32'd5847
; 
32'd158808: dataIn1 = 32'd5848
; 
32'd158809: dataIn1 = 32'd5849
; 
32'd158810: dataIn1 = 32'd6908
; 
32'd158811: dataIn1 = 32'd6909
; 
32'd158812: dataIn1 = 32'd6913
; 
32'd158813: dataIn1 = 32'd6915
; 
32'd158814: dataIn1 = 32'd6917
; 
32'd158815: dataIn1 = 32'd6918
; 
32'd158816: dataIn1 = 32'd5850
; 
32'd158817: dataIn1 = 32'd6907
; 
32'd158818: dataIn1 = 32'd6909
; 
32'd158819: dataIn1 = 32'd6911
; 
32'd158820: dataIn1 = 32'd6914
; 
32'd158821: dataIn1 = 32'd6923
; 
32'd158822: dataIn1 = 32'd6925
; 
32'd158823: dataIn1 = 32'd5851
; 
32'd158824: dataIn1 = 32'd6907
; 
32'd158825: dataIn1 = 32'd6908
; 
32'd158826: dataIn1 = 32'd6910
; 
32'd158827: dataIn1 = 32'd6912
; 
32'd158828: dataIn1 = 32'd6930
; 
32'd158829: dataIn1 = 32'd6931
; 
32'd158830: dataIn1 = 32'd5852
; 
32'd158831: dataIn1 = 32'd6916
; 
32'd158832: dataIn1 = 32'd6918
; 
32'd158833: dataIn1 = 32'd6920
; 
32'd158834: dataIn1 = 32'd6922
; 
32'd158835: dataIn1 = 32'd6981
; 
32'd158836: dataIn1 = 32'd6983
; 
32'd158837: dataIn1 = 32'd5853
; 
32'd158838: dataIn1 = 32'd6916
; 
32'd158839: dataIn1 = 32'd6917
; 
32'd158840: dataIn1 = 32'd6919
; 
32'd158841: dataIn1 = 32'd6921
; 
32'd158842: dataIn1 = 32'd6961
; 
32'd158843: dataIn1 = 32'd6962
; 
32'd158844: dataIn1 = 32'd5854
; 
32'd158845: dataIn1 = 32'd6924
; 
32'd158846: dataIn1 = 32'd6925
; 
32'd158847: dataIn1 = 32'd6928
; 
32'd158848: dataIn1 = 32'd6929
; 
32'd158849: dataIn1 = 32'd6985
; 
32'd158850: dataIn1 = 32'd6986
; 
32'd158851: dataIn1 = 32'd5855
; 
32'd158852: dataIn1 = 32'd6923
; 
32'd158853: dataIn1 = 32'd6924
; 
32'd158854: dataIn1 = 32'd6926
; 
32'd158855: dataIn1 = 32'd6927
; 
32'd158856: dataIn1 = 32'd6946
; 
32'd158857: dataIn1 = 32'd6947
; 
32'd158858: dataIn1 = 32'd5856
; 
32'd158859: dataIn1 = 32'd6931
; 
32'd158860: dataIn1 = 32'd6932
; 
32'd158861: dataIn1 = 32'd6934
; 
32'd158862: dataIn1 = 32'd6936
; 
32'd158863: dataIn1 = 32'd6968
; 
32'd158864: dataIn1 = 32'd6969
; 
32'd158865: dataIn1 = 32'd4837
; 
32'd158866: dataIn1 = 32'd5857
; 
32'd158867: dataIn1 = 32'd6930
; 
32'd158868: dataIn1 = 32'd6932
; 
32'd158869: dataIn1 = 32'd6933
; 
32'd158870: dataIn1 = 32'd6935
; 
32'd158871: dataIn1 = 32'd6951
; 
32'd158872: dataIn1 = 32'd2621
; 
32'd158873: dataIn1 = 32'd4836
; 
32'd158874: dataIn1 = 32'd5858
; 
32'd158875: dataIn1 = 32'd6938
; 
32'd158876: dataIn1 = 32'd6939
; 
32'd158877: dataIn1 = 32'd6943
; 
32'd158878: dataIn1 = 32'd6945
; 
32'd158879: dataIn1 = 32'd5859
; 
32'd158880: dataIn1 = 32'd6937
; 
32'd158881: dataIn1 = 32'd6939
; 
32'd158882: dataIn1 = 32'd6941
; 
32'd158883: dataIn1 = 32'd6942
; 
32'd158884: dataIn1 = 32'd6946
; 
32'd158885: dataIn1 = 32'd6948
; 
32'd158886: dataIn1 = 32'd2621
; 
32'd158887: dataIn1 = 32'd4837
; 
32'd158888: dataIn1 = 32'd5860
; 
32'd158889: dataIn1 = 32'd6937
; 
32'd158890: dataIn1 = 32'd6938
; 
32'd158891: dataIn1 = 32'd6940
; 
32'd158892: dataIn1 = 32'd6951
; 
32'd158893: dataIn1 = 32'd4
; 
32'd158894: dataIn1 = 32'd4836
; 
32'd158895: dataIn1 = 32'd5861
; 
32'd158896: dataIn1 = 32'd6944
; 
32'd158897: dataIn1 = 32'd6945
; 
32'd158898: dataIn1 = 32'd8902
; 
32'd158899: dataIn1 = 32'd8903
; 
32'd158900: dataIn1 = 32'd5862
; 
32'd158901: dataIn1 = 32'd6947
; 
32'd158902: dataIn1 = 32'd6948
; 
32'd158903: dataIn1 = 32'd6949
; 
32'd158904: dataIn1 = 32'd6950
; 
32'd158905: dataIn1 = 32'd8909
; 
32'd158906: dataIn1 = 32'd8910
; 
32'd158907: dataIn1 = 32'd5863
; 
32'd158908: dataIn1 = 32'd6953
; 
32'd158909: dataIn1 = 32'd6954
; 
32'd158910: dataIn1 = 32'd6958
; 
32'd158911: dataIn1 = 32'd6960
; 
32'd158912: dataIn1 = 32'd6962
; 
32'd158913: dataIn1 = 32'd6963
; 
32'd158914: dataIn1 = 32'd5864
; 
32'd158915: dataIn1 = 32'd6952
; 
32'd158916: dataIn1 = 32'd6954
; 
32'd158917: dataIn1 = 32'd6956
; 
32'd158918: dataIn1 = 32'd6959
; 
32'd158919: dataIn1 = 32'd6964
; 
32'd158920: dataIn1 = 32'd6966
; 
32'd158921: dataIn1 = 32'd5865
; 
32'd158922: dataIn1 = 32'd6952
; 
32'd158923: dataIn1 = 32'd6953
; 
32'd158924: dataIn1 = 32'd6955
; 
32'd158925: dataIn1 = 32'd6957
; 
32'd158926: dataIn1 = 32'd6967
; 
32'd158927: dataIn1 = 32'd6968
; 
32'd158928: dataIn1 = 32'd5866
; 
32'd158929: dataIn1 = 32'd6973
; 
32'd158930: dataIn1 = 32'd6974
; 
32'd158931: dataIn1 = 32'd6978
; 
32'd158932: dataIn1 = 32'd6980
; 
32'd158933: dataIn1 = 32'd6982
; 
32'd158934: dataIn1 = 32'd6983
; 
32'd158935: dataIn1 = 32'd5867
; 
32'd158936: dataIn1 = 32'd6972
; 
32'd158937: dataIn1 = 32'd6974
; 
32'd158938: dataIn1 = 32'd6976
; 
32'd158939: dataIn1 = 32'd6979
; 
32'd158940: dataIn1 = 32'd6984
; 
32'd158941: dataIn1 = 32'd6986
; 
32'd158942: dataIn1 = 32'd5847
; 
32'd158943: dataIn1 = 32'd5868
; 
32'd158944: dataIn1 = 32'd5870
; 
32'd158945: dataIn1 = 32'd6972
; 
32'd158946: dataIn1 = 32'd6973
; 
32'd158947: dataIn1 = 32'd6975
; 
32'd158948: dataIn1 = 32'd6977
; 
32'd158949: dataIn1 = 32'd5869
; 
32'd158950: dataIn1 = 32'd6984
; 
32'd158951: dataIn1 = 32'd6985
; 
32'd158952: dataIn1 = 32'd6987
; 
32'd158953: dataIn1 = 32'd6988
; 
32'd158954: dataIn1 = 32'd8911
; 
32'd158955: dataIn1 = 32'd8913
; 
32'd158956: dataIn1 = 32'd452
; 
32'd158957: dataIn1 = 32'd3976
; 
32'd158958: dataIn1 = 32'd5847
; 
32'd158959: dataIn1 = 32'd5868
; 
32'd158960: dataIn1 = 32'd5870
; 
32'd158961: dataIn1 = 32'd6586
; 
32'd158962: dataIn1 = 32'd6589
; 
32'd158963: dataIn1 = 32'd6975
; 
32'd158964: dataIn1 = 32'd5871
; 
32'd158965: dataIn1 = 32'd6990
; 
32'd158966: dataIn1 = 32'd6991
; 
32'd158967: dataIn1 = 32'd6995
; 
32'd158968: dataIn1 = 32'd6997
; 
32'd158969: dataIn1 = 32'd6999
; 
32'd158970: dataIn1 = 32'd7000
; 
32'd158971: dataIn1 = 32'd5872
; 
32'd158972: dataIn1 = 32'd6989
; 
32'd158973: dataIn1 = 32'd6991
; 
32'd158974: dataIn1 = 32'd6993
; 
32'd158975: dataIn1 = 32'd6996
; 
32'd158976: dataIn1 = 32'd7005
; 
32'd158977: dataIn1 = 32'd7007
; 
32'd158978: dataIn1 = 32'd5873
; 
32'd158979: dataIn1 = 32'd6989
; 
32'd158980: dataIn1 = 32'd6990
; 
32'd158981: dataIn1 = 32'd6992
; 
32'd158982: dataIn1 = 32'd6994
; 
32'd158983: dataIn1 = 32'd7010
; 
32'd158984: dataIn1 = 32'd7011
; 
32'd158985: dataIn1 = 32'd5874
; 
32'd158986: dataIn1 = 32'd6998
; 
32'd158987: dataIn1 = 32'd7000
; 
32'd158988: dataIn1 = 32'd7002
; 
32'd158989: dataIn1 = 32'd7004
; 
32'd158990: dataIn1 = 32'd7044
; 
32'd158991: dataIn1 = 32'd7046
; 
32'd158992: dataIn1 = 32'd5875
; 
32'd158993: dataIn1 = 32'd6998
; 
32'd158994: dataIn1 = 32'd6999
; 
32'd158995: dataIn1 = 32'd7001
; 
32'd158996: dataIn1 = 32'd7003
; 
32'd158997: dataIn1 = 32'd7026
; 
32'd158998: dataIn1 = 32'd7027
; 
32'd158999: dataIn1 = 32'd2325
; 
32'd159000: dataIn1 = 32'd5876
; 
32'd159001: dataIn1 = 32'd7006
; 
32'd159002: dataIn1 = 32'd7007
; 
32'd159003: dataIn1 = 32'd7009
; 
32'd159004: dataIn1 = 32'd7048
; 
32'd159005: dataIn1 = 32'd7049
; 
32'd159006: dataIn1 = 32'd2325
; 
32'd159007: dataIn1 = 32'd5877
; 
32'd159008: dataIn1 = 32'd7005
; 
32'd159009: dataIn1 = 32'd7006
; 
32'd159010: dataIn1 = 32'd7008
; 
32'd159011: dataIn1 = 32'd9272
; 
32'd159012: dataIn1 = 32'd9273
; 
32'd159013: dataIn1 = 32'd5878
; 
32'd159014: dataIn1 = 32'd7011
; 
32'd159015: dataIn1 = 32'd7012
; 
32'd159016: dataIn1 = 32'd7014
; 
32'd159017: dataIn1 = 32'd7016
; 
32'd159018: dataIn1 = 32'd7033
; 
32'd159019: dataIn1 = 32'd7034
; 
32'd159020: dataIn1 = 32'd5834
; 
32'd159021: dataIn1 = 32'd5879
; 
32'd159022: dataIn1 = 32'd5880
; 
32'd159023: dataIn1 = 32'd7010
; 
32'd159024: dataIn1 = 32'd7012
; 
32'd159025: dataIn1 = 32'd7013
; 
32'd159026: dataIn1 = 32'd7015
; 
32'd159027: dataIn1 = 32'd3966
; 
32'd159028: dataIn1 = 32'd3981
; 
32'd159029: dataIn1 = 32'd5834
; 
32'd159030: dataIn1 = 32'd5879
; 
32'd159031: dataIn1 = 32'd5880
; 
32'd159032: dataIn1 = 32'd7013
; 
32'd159033: dataIn1 = 32'd9273
; 
32'd159034: dataIn1 = 32'd9320
; 
32'd159035: dataIn1 = 32'd5881
; 
32'd159036: dataIn1 = 32'd7018
; 
32'd159037: dataIn1 = 32'd7019
; 
32'd159038: dataIn1 = 32'd7023
; 
32'd159039: dataIn1 = 32'd7025
; 
32'd159040: dataIn1 = 32'd7027
; 
32'd159041: dataIn1 = 32'd7028
; 
32'd159042: dataIn1 = 32'd5882
; 
32'd159043: dataIn1 = 32'd7017
; 
32'd159044: dataIn1 = 32'd7019
; 
32'd159045: dataIn1 = 32'd7021
; 
32'd159046: dataIn1 = 32'd7024
; 
32'd159047: dataIn1 = 32'd7029
; 
32'd159048: dataIn1 = 32'd7031
; 
32'd159049: dataIn1 = 32'd5883
; 
32'd159050: dataIn1 = 32'd7017
; 
32'd159051: dataIn1 = 32'd7018
; 
32'd159052: dataIn1 = 32'd7020
; 
32'd159053: dataIn1 = 32'd7022
; 
32'd159054: dataIn1 = 32'd7032
; 
32'd159055: dataIn1 = 32'd7033
; 
32'd159056: dataIn1 = 32'd5884
; 
32'd159057: dataIn1 = 32'd7036
; 
32'd159058: dataIn1 = 32'd7037
; 
32'd159059: dataIn1 = 32'd7041
; 
32'd159060: dataIn1 = 32'd7043
; 
32'd159061: dataIn1 = 32'd7045
; 
32'd159062: dataIn1 = 32'd7046
; 
32'd159063: dataIn1 = 32'd5885
; 
32'd159064: dataIn1 = 32'd7035
; 
32'd159065: dataIn1 = 32'd7037
; 
32'd159066: dataIn1 = 32'd7039
; 
32'd159067: dataIn1 = 32'd7042
; 
32'd159068: dataIn1 = 32'd7047
; 
32'd159069: dataIn1 = 32'd7049
; 
32'd159070: dataIn1 = 32'd5886
; 
32'd159071: dataIn1 = 32'd7035
; 
32'd159072: dataIn1 = 32'd7036
; 
32'd159073: dataIn1 = 32'd7038
; 
32'd159074: dataIn1 = 32'd7040
; 
32'd159075: dataIn1 = 32'd7051
; 
32'd159076: dataIn1 = 32'd7052
; 
32'd159077: dataIn1 = 32'd2325
; 
32'd159078: dataIn1 = 32'd5887
; 
32'd159079: dataIn1 = 32'd6598
; 
32'd159080: dataIn1 = 32'd7047
; 
32'd159081: dataIn1 = 32'd7048
; 
32'd159082: dataIn1 = 32'd7050
; 
32'd159083: dataIn1 = 32'd9779
; 
32'd159084: dataIn1 = 32'd5888
; 
32'd159085: dataIn1 = 32'd7051
; 
32'd159086: dataIn1 = 32'd7053
; 
32'd159087: dataIn1 = 32'd7054
; 
32'd159088: dataIn1 = 32'd8921
; 
32'd159089: dataIn1 = 32'd8923
; 
32'd159090: dataIn1 = 32'd8925
; 
32'd159091: dataIn1 = 32'd4647
; 
32'd159092: dataIn1 = 32'd4650
; 
32'd159093: dataIn1 = 32'd4651
; 
32'd159094: dataIn1 = 32'd5889
; 
32'd159095: dataIn1 = 32'd5890
; 
32'd159096: dataIn1 = 32'd5891
; 
32'd159097: dataIn1 = 32'd209
; 
32'd159098: dataIn1 = 32'd4651
; 
32'd159099: dataIn1 = 32'd5889
; 
32'd159100: dataIn1 = 32'd5890
; 
32'd159101: dataIn1 = 32'd5891
; 
32'd159102: dataIn1 = 32'd5917
; 
32'd159103: dataIn1 = 32'd5920
; 
32'd159104: dataIn1 = 32'd209
; 
32'd159105: dataIn1 = 32'd4650
; 
32'd159106: dataIn1 = 32'd5889
; 
32'd159107: dataIn1 = 32'd5890
; 
32'd159108: dataIn1 = 32'd5891
; 
32'd159109: dataIn1 = 32'd5927
; 
32'd159110: dataIn1 = 32'd5930
; 
32'd159111: dataIn1 = 32'd2558
; 
32'd159112: dataIn1 = 32'd4657
; 
32'd159113: dataIn1 = 32'd4658
; 
32'd159114: dataIn1 = 32'd5892
; 
32'd159115: dataIn1 = 32'd5893
; 
32'd159116: dataIn1 = 32'd5894
; 
32'd159117: dataIn1 = 32'd4656
; 
32'd159118: dataIn1 = 32'd4658
; 
32'd159119: dataIn1 = 32'd5892
; 
32'd159120: dataIn1 = 32'd5893
; 
32'd159121: dataIn1 = 32'd5894
; 
32'd159122: dataIn1 = 32'd5895
; 
32'd159123: dataIn1 = 32'd5896
; 
32'd159124: dataIn1 = 32'd4656
; 
32'd159125: dataIn1 = 32'd4657
; 
32'd159126: dataIn1 = 32'd5892
; 
32'd159127: dataIn1 = 32'd5893
; 
32'd159128: dataIn1 = 32'd5894
; 
32'd159129: dataIn1 = 32'd5897
; 
32'd159130: dataIn1 = 32'd5898
; 
32'd159131: dataIn1 = 32'd2561
; 
32'd159132: dataIn1 = 32'd4658
; 
32'd159133: dataIn1 = 32'd5893
; 
32'd159134: dataIn1 = 32'd5895
; 
32'd159135: dataIn1 = 32'd5896
; 
32'd159136: dataIn1 = 32'd5912
; 
32'd159137: dataIn1 = 32'd5913
; 
32'd159138: dataIn1 = 32'd2561
; 
32'd159139: dataIn1 = 32'd4656
; 
32'd159140: dataIn1 = 32'd5893
; 
32'd159141: dataIn1 = 32'd5895
; 
32'd159142: dataIn1 = 32'd5896
; 
32'd159143: dataIn1 = 32'd5900
; 
32'd159144: dataIn1 = 32'd5904
; 
32'd159145: dataIn1 = 32'd2562
; 
32'd159146: dataIn1 = 32'd4657
; 
32'd159147: dataIn1 = 32'd5894
; 
32'd159148: dataIn1 = 32'd5897
; 
32'd159149: dataIn1 = 32'd5898
; 
32'd159150: dataIn1 = 32'd5908
; 
32'd159151: dataIn1 = 32'd5911
; 
32'd159152: dataIn1 = 32'd2562
; 
32'd159153: dataIn1 = 32'd4656
; 
32'd159154: dataIn1 = 32'd5894
; 
32'd159155: dataIn1 = 32'd5897
; 
32'd159156: dataIn1 = 32'd5898
; 
32'd159157: dataIn1 = 32'd5901
; 
32'd159158: dataIn1 = 32'd5905
; 
32'd159159: dataIn1 = 32'd4659
; 
32'd159160: dataIn1 = 32'd4660
; 
32'd159161: dataIn1 = 32'd5899
; 
32'd159162: dataIn1 = 32'd5900
; 
32'd159163: dataIn1 = 32'd5901
; 
32'd159164: dataIn1 = 32'd5902
; 
32'd159165: dataIn1 = 32'd5903
; 
32'd159166: dataIn1 = 32'd4656
; 
32'd159167: dataIn1 = 32'd4660
; 
32'd159168: dataIn1 = 32'd5896
; 
32'd159169: dataIn1 = 32'd5899
; 
32'd159170: dataIn1 = 32'd5900
; 
32'd159171: dataIn1 = 32'd5901
; 
32'd159172: dataIn1 = 32'd5904
; 
32'd159173: dataIn1 = 32'd4656
; 
32'd159174: dataIn1 = 32'd4659
; 
32'd159175: dataIn1 = 32'd5898
; 
32'd159176: dataIn1 = 32'd5899
; 
32'd159177: dataIn1 = 32'd5900
; 
32'd159178: dataIn1 = 32'd5901
; 
32'd159179: dataIn1 = 32'd5905
; 
32'd159180: dataIn1 = 32'd130
; 
32'd159181: dataIn1 = 32'd4660
; 
32'd159182: dataIn1 = 32'd5899
; 
32'd159183: dataIn1 = 32'd5902
; 
32'd159184: dataIn1 = 32'd5903
; 
32'd159185: dataIn1 = 32'd5969
; 
32'd159186: dataIn1 = 32'd5972
; 
32'd159187: dataIn1 = 32'd130
; 
32'd159188: dataIn1 = 32'd4659
; 
32'd159189: dataIn1 = 32'd5899
; 
32'd159190: dataIn1 = 32'd5902
; 
32'd159191: dataIn1 = 32'd5903
; 
32'd159192: dataIn1 = 32'd6030
; 
32'd159193: dataIn1 = 32'd6033
; 
32'd159194: dataIn1 = 32'd2561
; 
32'd159195: dataIn1 = 32'd4660
; 
32'd159196: dataIn1 = 32'd5896
; 
32'd159197: dataIn1 = 32'd5900
; 
32'd159198: dataIn1 = 32'd5904
; 
32'd159199: dataIn1 = 32'd5966
; 
32'd159200: dataIn1 = 32'd5970
; 
32'd159201: dataIn1 = 32'd2562
; 
32'd159202: dataIn1 = 32'd4659
; 
32'd159203: dataIn1 = 32'd5898
; 
32'd159204: dataIn1 = 32'd5901
; 
32'd159205: dataIn1 = 32'd5905
; 
32'd159206: dataIn1 = 32'd6029
; 
32'd159207: dataIn1 = 32'd6032
; 
32'd159208: dataIn1 = 32'd2558
; 
32'd159209: dataIn1 = 32'd4653
; 
32'd159210: dataIn1 = 32'd4657
; 
32'd159211: dataIn1 = 32'd5906
; 
32'd159212: dataIn1 = 32'd5907
; 
32'd159213: dataIn1 = 32'd5908
; 
32'd159214: dataIn1 = 32'd4653
; 
32'd159215: dataIn1 = 32'd4661
; 
32'd159216: dataIn1 = 32'd5906
; 
32'd159217: dataIn1 = 32'd5907
; 
32'd159218: dataIn1 = 32'd5908
; 
32'd159219: dataIn1 = 32'd5909
; 
32'd159220: dataIn1 = 32'd5910
; 
32'd159221: dataIn1 = 32'd4657
; 
32'd159222: dataIn1 = 32'd4661
; 
32'd159223: dataIn1 = 32'd5897
; 
32'd159224: dataIn1 = 32'd5906
; 
32'd159225: dataIn1 = 32'd5907
; 
32'd159226: dataIn1 = 32'd5908
; 
32'd159227: dataIn1 = 32'd5911
; 
32'd159228: dataIn1 = 32'd1074
; 
32'd159229: dataIn1 = 32'd4652
; 
32'd159230: dataIn1 = 32'd4653
; 
32'd159231: dataIn1 = 32'd5907
; 
32'd159232: dataIn1 = 32'd5909
; 
32'd159233: dataIn1 = 32'd5910
; 
32'd159234: dataIn1 = 32'd1074
; 
32'd159235: dataIn1 = 32'd4661
; 
32'd159236: dataIn1 = 32'd5907
; 
32'd159237: dataIn1 = 32'd5909
; 
32'd159238: dataIn1 = 32'd5910
; 
32'd159239: dataIn1 = 32'd6036
; 
32'd159240: dataIn1 = 32'd6697
; 
32'd159241: dataIn1 = 32'd2562
; 
32'd159242: dataIn1 = 32'd4661
; 
32'd159243: dataIn1 = 32'd5897
; 
32'd159244: dataIn1 = 32'd5908
; 
32'd159245: dataIn1 = 32'd5911
; 
32'd159246: dataIn1 = 32'd6028
; 
32'd159247: dataIn1 = 32'd6037
; 
32'd159248: dataIn1 = 32'd4655
; 
32'd159249: dataIn1 = 32'd4658
; 
32'd159250: dataIn1 = 32'd4662
; 
32'd159251: dataIn1 = 32'd5895
; 
32'd159252: dataIn1 = 32'd5912
; 
32'd159253: dataIn1 = 32'd5913
; 
32'd159254: dataIn1 = 32'd2561
; 
32'd159255: dataIn1 = 32'd4662
; 
32'd159256: dataIn1 = 32'd5895
; 
32'd159257: dataIn1 = 32'd5912
; 
32'd159258: dataIn1 = 32'd5913
; 
32'd159259: dataIn1 = 32'd5965
; 
32'd159260: dataIn1 = 32'd5979
; 
32'd159261: dataIn1 = 32'd1041
; 
32'd159262: dataIn1 = 32'd4622
; 
32'd159263: dataIn1 = 32'd4664
; 
32'd159264: dataIn1 = 32'd5914
; 
32'd159265: dataIn1 = 32'd5915
; 
32'd159266: dataIn1 = 32'd5916
; 
32'd159267: dataIn1 = 32'd5923
; 
32'd159268: dataIn1 = 32'd1041
; 
32'd159269: dataIn1 = 32'd4616
; 
32'd159270: dataIn1 = 32'd4663
; 
32'd159271: dataIn1 = 32'd5914
; 
32'd159272: dataIn1 = 32'd5915
; 
32'd159273: dataIn1 = 32'd5916
; 
32'd159274: dataIn1 = 32'd5919
; 
32'd159275: dataIn1 = 32'd4663
; 
32'd159276: dataIn1 = 32'd4664
; 
32'd159277: dataIn1 = 32'd4665
; 
32'd159278: dataIn1 = 32'd5914
; 
32'd159279: dataIn1 = 32'd5915
; 
32'd159280: dataIn1 = 32'd5916
; 
32'd159281: dataIn1 = 32'd2542
; 
32'd159282: dataIn1 = 32'd4651
; 
32'd159283: dataIn1 = 32'd5890
; 
32'd159284: dataIn1 = 32'd5917
; 
32'd159285: dataIn1 = 32'd5918
; 
32'd159286: dataIn1 = 32'd5919
; 
32'd159287: dataIn1 = 32'd5920
; 
32'd159288: dataIn1 = 32'd2559
; 
32'd159289: dataIn1 = 32'd4651
; 
32'd159290: dataIn1 = 32'd4663
; 
32'd159291: dataIn1 = 32'd5917
; 
32'd159292: dataIn1 = 32'd5918
; 
32'd159293: dataIn1 = 32'd5919
; 
32'd159294: dataIn1 = 32'd2542
; 
32'd159295: dataIn1 = 32'd4616
; 
32'd159296: dataIn1 = 32'd4663
; 
32'd159297: dataIn1 = 32'd5915
; 
32'd159298: dataIn1 = 32'd5917
; 
32'd159299: dataIn1 = 32'd5918
; 
32'd159300: dataIn1 = 32'd5919
; 
32'd159301: dataIn1 = 32'd209
; 
32'd159302: dataIn1 = 32'd2530
; 
32'd159303: dataIn1 = 32'd2542
; 
32'd159304: dataIn1 = 32'd5890
; 
32'd159305: dataIn1 = 32'd5917
; 
32'd159306: dataIn1 = 32'd5920
; 
32'd159307: dataIn1 = 32'd2563
; 
32'd159308: dataIn1 = 32'd4664
; 
32'd159309: dataIn1 = 32'd4666
; 
32'd159310: dataIn1 = 32'd5921
; 
32'd159311: dataIn1 = 32'd5922
; 
32'd159312: dataIn1 = 32'd5923
; 
32'd159313: dataIn1 = 32'd2543
; 
32'd159314: dataIn1 = 32'd4621
; 
32'd159315: dataIn1 = 32'd4666
; 
32'd159316: dataIn1 = 32'd5921
; 
32'd159317: dataIn1 = 32'd5922
; 
32'd159318: dataIn1 = 32'd5923
; 
32'd159319: dataIn1 = 32'd5980
; 
32'd159320: dataIn1 = 32'd2543
; 
32'd159321: dataIn1 = 32'd4622
; 
32'd159322: dataIn1 = 32'd4664
; 
32'd159323: dataIn1 = 32'd5914
; 
32'd159324: dataIn1 = 32'd5921
; 
32'd159325: dataIn1 = 32'd5922
; 
32'd159326: dataIn1 = 32'd5923
; 
32'd159327: dataIn1 = 32'd1040
; 
32'd159328: dataIn1 = 32'd4670
; 
32'd159329: dataIn1 = 32'd5924
; 
32'd159330: dataIn1 = 32'd5925
; 
32'd159331: dataIn1 = 32'd5926
; 
32'd159332: dataIn1 = 32'd5933
; 
32'd159333: dataIn1 = 32'd5935
; 
32'd159334: dataIn1 = 32'd4668
; 
32'd159335: dataIn1 = 32'd4669
; 
32'd159336: dataIn1 = 32'd4670
; 
32'd159337: dataIn1 = 32'd5924
; 
32'd159338: dataIn1 = 32'd5925
; 
32'd159339: dataIn1 = 32'd5926
; 
32'd159340: dataIn1 = 32'd1040
; 
32'd159341: dataIn1 = 32'd4668
; 
32'd159342: dataIn1 = 32'd5924
; 
32'd159343: dataIn1 = 32'd5925
; 
32'd159344: dataIn1 = 32'd5926
; 
32'd159345: dataIn1 = 32'd5928
; 
32'd159346: dataIn1 = 32'd5931
; 
32'd159347: dataIn1 = 32'd2538
; 
32'd159348: dataIn1 = 32'd4650
; 
32'd159349: dataIn1 = 32'd5891
; 
32'd159350: dataIn1 = 32'd5927
; 
32'd159351: dataIn1 = 32'd5928
; 
32'd159352: dataIn1 = 32'd5929
; 
32'd159353: dataIn1 = 32'd5930
; 
32'd159354: dataIn1 = 32'd2538
; 
32'd159355: dataIn1 = 32'd4668
; 
32'd159356: dataIn1 = 32'd5926
; 
32'd159357: dataIn1 = 32'd5927
; 
32'd159358: dataIn1 = 32'd5928
; 
32'd159359: dataIn1 = 32'd5929
; 
32'd159360: dataIn1 = 32'd5931
; 
32'd159361: dataIn1 = 32'd2560
; 
32'd159362: dataIn1 = 32'd4650
; 
32'd159363: dataIn1 = 32'd4668
; 
32'd159364: dataIn1 = 32'd5927
; 
32'd159365: dataIn1 = 32'd5928
; 
32'd159366: dataIn1 = 32'd5929
; 
32'd159367: dataIn1 = 32'd209
; 
32'd159368: dataIn1 = 32'd2529
; 
32'd159369: dataIn1 = 32'd2538
; 
32'd159370: dataIn1 = 32'd5891
; 
32'd159371: dataIn1 = 32'd5927
; 
32'd159372: dataIn1 = 32'd5930
; 
32'd159373: dataIn1 = 32'd1040
; 
32'd159374: dataIn1 = 32'd2536
; 
32'd159375: dataIn1 = 32'd2538
; 
32'd159376: dataIn1 = 32'd5926
; 
32'd159377: dataIn1 = 32'd5928
; 
32'd159378: dataIn1 = 32'd5931
; 
32'd159379: dataIn1 = 32'd2564
; 
32'd159380: dataIn1 = 32'd4670
; 
32'd159381: dataIn1 = 32'd4672
; 
32'd159382: dataIn1 = 32'd5932
; 
32'd159383: dataIn1 = 32'd5933
; 
32'd159384: dataIn1 = 32'd5934
; 
32'd159385: dataIn1 = 32'd2539
; 
32'd159386: dataIn1 = 32'd4670
; 
32'd159387: dataIn1 = 32'd5924
; 
32'd159388: dataIn1 = 32'd5932
; 
32'd159389: dataIn1 = 32'd5933
; 
32'd159390: dataIn1 = 32'd5934
; 
32'd159391: dataIn1 = 32'd5935
; 
32'd159392: dataIn1 = 32'd2539
; 
32'd159393: dataIn1 = 32'd4672
; 
32'd159394: dataIn1 = 32'd5932
; 
32'd159395: dataIn1 = 32'd5933
; 
32'd159396: dataIn1 = 32'd5934
; 
32'd159397: dataIn1 = 32'd5936
; 
32'd159398: dataIn1 = 32'd5937
; 
32'd159399: dataIn1 = 32'd1040
; 
32'd159400: dataIn1 = 32'd2537
; 
32'd159401: dataIn1 = 32'd2539
; 
32'd159402: dataIn1 = 32'd5924
; 
32'd159403: dataIn1 = 32'd5933
; 
32'd159404: dataIn1 = 32'd5935
; 
32'd159405: dataIn1 = 32'd129
; 
32'd159406: dataIn1 = 32'd4672
; 
32'd159407: dataIn1 = 32'd5721
; 
32'd159408: dataIn1 = 32'd5934
; 
32'd159409: dataIn1 = 32'd5936
; 
32'd159410: dataIn1 = 32'd5937
; 
32'd159411: dataIn1 = 32'd6063
; 
32'd159412: dataIn1 = 32'd129
; 
32'd159413: dataIn1 = 32'd2528
; 
32'd159414: dataIn1 = 32'd2539
; 
32'd159415: dataIn1 = 32'd5934
; 
32'd159416: dataIn1 = 32'd5936
; 
32'd159417: dataIn1 = 32'd5937
; 
32'd159418: dataIn1 = 32'd6
; 
32'd159419: dataIn1 = 32'd4679
; 
32'd159420: dataIn1 = 32'd5938
; 
32'd159421: dataIn1 = 32'd5939
; 
32'd159422: dataIn1 = 32'd5940
; 
32'd159423: dataIn1 = 32'd6065
; 
32'd159424: dataIn1 = 32'd6066
; 
32'd159425: dataIn1 = 32'd4674
; 
32'd159426: dataIn1 = 32'd4678
; 
32'd159427: dataIn1 = 32'd4679
; 
32'd159428: dataIn1 = 32'd5938
; 
32'd159429: dataIn1 = 32'd5939
; 
32'd159430: dataIn1 = 32'd5940
; 
32'd159431: dataIn1 = 32'd6
; 
32'd159432: dataIn1 = 32'd4678
; 
32'd159433: dataIn1 = 32'd5938
; 
32'd159434: dataIn1 = 32'd5939
; 
32'd159435: dataIn1 = 32'd5940
; 
32'd159436: dataIn1 = 32'd5993
; 
32'd159437: dataIn1 = 32'd5995
; 
32'd159438: dataIn1 = 32'd3883
; 
32'd159439: dataIn1 = 32'd4830
; 
32'd159440: dataIn1 = 32'd5667
; 
32'd159441: dataIn1 = 32'd5941
; 
32'd159442: dataIn1 = 32'd5942
; 
32'd159443: dataIn1 = 32'd5943
; 
32'd159444: dataIn1 = 32'd5944
; 
32'd159445: dataIn1 = 32'd4827
; 
32'd159446: dataIn1 = 32'd4830
; 
32'd159447: dataIn1 = 32'd5941
; 
32'd159448: dataIn1 = 32'd5942
; 
32'd159449: dataIn1 = 32'd5943
; 
32'd159450: dataIn1 = 32'd5945
; 
32'd159451: dataIn1 = 32'd5946
; 
32'd159452: dataIn1 = 32'd2300
; 
32'd159453: dataIn1 = 32'd3883
; 
32'd159454: dataIn1 = 32'd4827
; 
32'd159455: dataIn1 = 32'd5941
; 
32'd159456: dataIn1 = 32'd5942
; 
32'd159457: dataIn1 = 32'd5943
; 
32'd159458: dataIn1 = 32'd127
; 
32'd159459: dataIn1 = 32'd4830
; 
32'd159460: dataIn1 = 32'd5667
; 
32'd159461: dataIn1 = 32'd5941
; 
32'd159462: dataIn1 = 32'd5944
; 
32'd159463: dataIn1 = 32'd6893
; 
32'd159464: dataIn1 = 32'd6965
; 
32'd159465: dataIn1 = 32'd2620
; 
32'd159466: dataIn1 = 32'd4830
; 
32'd159467: dataIn1 = 32'd5942
; 
32'd159468: dataIn1 = 32'd5945
; 
32'd159469: dataIn1 = 32'd5946
; 
32'd159470: dataIn1 = 32'd6956
; 
32'd159471: dataIn1 = 32'd6964
; 
32'd159472: dataIn1 = 32'd2620
; 
32'd159473: dataIn1 = 32'd4827
; 
32'd159474: dataIn1 = 32'd4829
; 
32'd159475: dataIn1 = 32'd5942
; 
32'd159476: dataIn1 = 32'd5945
; 
32'd159477: dataIn1 = 32'd5946
; 
32'd159478: dataIn1 = 32'd3899
; 
32'd159479: dataIn1 = 32'd4838
; 
32'd159480: dataIn1 = 32'd5691
; 
32'd159481: dataIn1 = 32'd5947
; 
32'd159482: dataIn1 = 32'd5948
; 
32'd159483: dataIn1 = 32'd5949
; 
32'd159484: dataIn1 = 32'd5950
; 
32'd159485: dataIn1 = 32'd2554
; 
32'd159486: dataIn1 = 32'd4643
; 
32'd159487: dataIn1 = 32'd4838
; 
32'd159488: dataIn1 = 32'd5947
; 
32'd159489: dataIn1 = 32'd5948
; 
32'd159490: dataIn1 = 32'd5949
; 
32'd159491: dataIn1 = 32'd3899
; 
32'd159492: dataIn1 = 32'd4643
; 
32'd159493: dataIn1 = 32'd5947
; 
32'd159494: dataIn1 = 32'd5948
; 
32'd159495: dataIn1 = 32'd5949
; 
32'd159496: dataIn1 = 32'd5951
; 
32'd159497: dataIn1 = 32'd5952
; 
32'd159498: dataIn1 = 32'd2302
; 
32'd159499: dataIn1 = 32'd4838
; 
32'd159500: dataIn1 = 32'd5318
; 
32'd159501: dataIn1 = 32'd5691
; 
32'd159502: dataIn1 = 32'd5947
; 
32'd159503: dataIn1 = 32'd5950
; 
32'd159504: dataIn1 = 32'd126
; 
32'd159505: dataIn1 = 32'd3866
; 
32'd159506: dataIn1 = 32'd3899
; 
32'd159507: dataIn1 = 32'd5690
; 
32'd159508: dataIn1 = 32'd5949
; 
32'd159509: dataIn1 = 32'd5951
; 
32'd159510: dataIn1 = 32'd5952
; 
32'd159511: dataIn1 = 32'd126
; 
32'd159512: dataIn1 = 32'd4610
; 
32'd159513: dataIn1 = 32'd4643
; 
32'd159514: dataIn1 = 32'd5949
; 
32'd159515: dataIn1 = 32'd5951
; 
32'd159516: dataIn1 = 32'd5952
; 
32'd159517: dataIn1 = 32'd6698
; 
32'd159518: dataIn1 = 32'd4840
; 
32'd159519: dataIn1 = 32'd4845
; 
32'd159520: dataIn1 = 32'd5953
; 
32'd159521: dataIn1 = 32'd5954
; 
32'd159522: dataIn1 = 32'd5955
; 
32'd159523: dataIn1 = 32'd5956
; 
32'd159524: dataIn1 = 32'd5957
; 
32'd159525: dataIn1 = 32'd4844
; 
32'd159526: dataIn1 = 32'd4845
; 
32'd159527: dataIn1 = 32'd5953
; 
32'd159528: dataIn1 = 32'd5954
; 
32'd159529: dataIn1 = 32'd5955
; 
32'd159530: dataIn1 = 32'd5958
; 
32'd159531: dataIn1 = 32'd5959
; 
32'd159532: dataIn1 = 32'd2624
; 
32'd159533: dataIn1 = 32'd4840
; 
32'd159534: dataIn1 = 32'd4844
; 
32'd159535: dataIn1 = 32'd5953
; 
32'd159536: dataIn1 = 32'd5954
; 
32'd159537: dataIn1 = 32'd5955
; 
32'd159538: dataIn1 = 32'd2622
; 
32'd159539: dataIn1 = 32'd4845
; 
32'd159540: dataIn1 = 32'd5953
; 
32'd159541: dataIn1 = 32'd5956
; 
32'd159542: dataIn1 = 32'd5957
; 
32'd159543: dataIn1 = 32'd5964
; 
32'd159544: dataIn1 = 32'd5974
; 
32'd159545: dataIn1 = 32'd2622
; 
32'd159546: dataIn1 = 32'd4840
; 
32'd159547: dataIn1 = 32'd4841
; 
32'd159548: dataIn1 = 32'd5953
; 
32'd159549: dataIn1 = 32'd5956
; 
32'd159550: dataIn1 = 32'd5957
; 
32'd159551: dataIn1 = 32'd1105
; 
32'd159552: dataIn1 = 32'd4845
; 
32'd159553: dataIn1 = 32'd5954
; 
32'd159554: dataIn1 = 32'd5958
; 
32'd159555: dataIn1 = 32'd5959
; 
32'd159556: dataIn1 = 32'd5975
; 
32'd159557: dataIn1 = 32'd5977
; 
32'd159558: dataIn1 = 32'd1105
; 
32'd159559: dataIn1 = 32'd4844
; 
32'd159560: dataIn1 = 32'd5954
; 
32'd159561: dataIn1 = 32'd5958
; 
32'd159562: dataIn1 = 32'd5959
; 
32'd159563: dataIn1 = 32'd5987
; 
32'd159564: dataIn1 = 32'd5990
; 
32'd159565: dataIn1 = 32'd4849
; 
32'd159566: dataIn1 = 32'd4850
; 
32'd159567: dataIn1 = 32'd5960
; 
32'd159568: dataIn1 = 32'd5961
; 
32'd159569: dataIn1 = 32'd5962
; 
32'd159570: dataIn1 = 32'd5963
; 
32'd159571: dataIn1 = 32'd5964
; 
32'd159572: dataIn1 = 32'd4848
; 
32'd159573: dataIn1 = 32'd4850
; 
32'd159574: dataIn1 = 32'd5960
; 
32'd159575: dataIn1 = 32'd5961
; 
32'd159576: dataIn1 = 32'd5962
; 
32'd159577: dataIn1 = 32'd5965
; 
32'd159578: dataIn1 = 32'd5966
; 
32'd159579: dataIn1 = 32'd4848
; 
32'd159580: dataIn1 = 32'd4849
; 
32'd159581: dataIn1 = 32'd5960
; 
32'd159582: dataIn1 = 32'd5961
; 
32'd159583: dataIn1 = 32'd5962
; 
32'd159584: dataIn1 = 32'd5967
; 
32'd159585: dataIn1 = 32'd5968
; 
32'd159586: dataIn1 = 32'd2622
; 
32'd159587: dataIn1 = 32'd4847
; 
32'd159588: dataIn1 = 32'd4850
; 
32'd159589: dataIn1 = 32'd5960
; 
32'd159590: dataIn1 = 32'd5963
; 
32'd159591: dataIn1 = 32'd5964
; 
32'd159592: dataIn1 = 32'd2622
; 
32'd159593: dataIn1 = 32'd4849
; 
32'd159594: dataIn1 = 32'd5956
; 
32'd159595: dataIn1 = 32'd5960
; 
32'd159596: dataIn1 = 32'd5963
; 
32'd159597: dataIn1 = 32'd5964
; 
32'd159598: dataIn1 = 32'd5974
; 
32'd159599: dataIn1 = 32'd2561
; 
32'd159600: dataIn1 = 32'd4850
; 
32'd159601: dataIn1 = 32'd5913
; 
32'd159602: dataIn1 = 32'd5961
; 
32'd159603: dataIn1 = 32'd5965
; 
32'd159604: dataIn1 = 32'd5966
; 
32'd159605: dataIn1 = 32'd5979
; 
32'd159606: dataIn1 = 32'd2561
; 
32'd159607: dataIn1 = 32'd4848
; 
32'd159608: dataIn1 = 32'd5904
; 
32'd159609: dataIn1 = 32'd5961
; 
32'd159610: dataIn1 = 32'd5965
; 
32'd159611: dataIn1 = 32'd5966
; 
32'd159612: dataIn1 = 32'd5970
; 
32'd159613: dataIn1 = 32'd2625
; 
32'd159614: dataIn1 = 32'd4849
; 
32'd159615: dataIn1 = 32'd5962
; 
32'd159616: dataIn1 = 32'd5967
; 
32'd159617: dataIn1 = 32'd5968
; 
32'd159618: dataIn1 = 32'd5976
; 
32'd159619: dataIn1 = 32'd5978
; 
32'd159620: dataIn1 = 32'd2625
; 
32'd159621: dataIn1 = 32'd4848
; 
32'd159622: dataIn1 = 32'd5962
; 
32'd159623: dataIn1 = 32'd5967
; 
32'd159624: dataIn1 = 32'd5968
; 
32'd159625: dataIn1 = 32'd5971
; 
32'd159626: dataIn1 = 32'd5973
; 
32'd159627: dataIn1 = 32'd4660
; 
32'd159628: dataIn1 = 32'd4851
; 
32'd159629: dataIn1 = 32'd5902
; 
32'd159630: dataIn1 = 32'd5969
; 
32'd159631: dataIn1 = 32'd5970
; 
32'd159632: dataIn1 = 32'd5971
; 
32'd159633: dataIn1 = 32'd5972
; 
32'd159634: dataIn1 = 32'd4660
; 
32'd159635: dataIn1 = 32'd4848
; 
32'd159636: dataIn1 = 32'd5904
; 
32'd159637: dataIn1 = 32'd5966
; 
32'd159638: dataIn1 = 32'd5969
; 
32'd159639: dataIn1 = 32'd5970
; 
32'd159640: dataIn1 = 32'd5971
; 
32'd159641: dataIn1 = 32'd4848
; 
32'd159642: dataIn1 = 32'd4851
; 
32'd159643: dataIn1 = 32'd5968
; 
32'd159644: dataIn1 = 32'd5969
; 
32'd159645: dataIn1 = 32'd5970
; 
32'd159646: dataIn1 = 32'd5971
; 
32'd159647: dataIn1 = 32'd5973
; 
32'd159648: dataIn1 = 32'd130
; 
32'd159649: dataIn1 = 32'd4851
; 
32'd159650: dataIn1 = 32'd5902
; 
32'd159651: dataIn1 = 32'd5969
; 
32'd159652: dataIn1 = 32'd5972
; 
32'd159653: dataIn1 = 32'd7237
; 
32'd159654: dataIn1 = 32'd7330
; 
32'd159655: dataIn1 = 32'd2625
; 
32'd159656: dataIn1 = 32'd4851
; 
32'd159657: dataIn1 = 32'd5968
; 
32'd159658: dataIn1 = 32'd5971
; 
32'd159659: dataIn1 = 32'd5973
; 
32'd159660: dataIn1 = 32'd7324
; 
32'd159661: dataIn1 = 32'd7331
; 
32'd159662: dataIn1 = 32'd4845
; 
32'd159663: dataIn1 = 32'd4849
; 
32'd159664: dataIn1 = 32'd5956
; 
32'd159665: dataIn1 = 32'd5964
; 
32'd159666: dataIn1 = 32'd5974
; 
32'd159667: dataIn1 = 32'd5975
; 
32'd159668: dataIn1 = 32'd5976
; 
32'd159669: dataIn1 = 32'd4845
; 
32'd159670: dataIn1 = 32'd4852
; 
32'd159671: dataIn1 = 32'd5958
; 
32'd159672: dataIn1 = 32'd5974
; 
32'd159673: dataIn1 = 32'd5975
; 
32'd159674: dataIn1 = 32'd5976
; 
32'd159675: dataIn1 = 32'd5977
; 
32'd159676: dataIn1 = 32'd4849
; 
32'd159677: dataIn1 = 32'd4852
; 
32'd159678: dataIn1 = 32'd5967
; 
32'd159679: dataIn1 = 32'd5974
; 
32'd159680: dataIn1 = 32'd5975
; 
32'd159681: dataIn1 = 32'd5976
; 
32'd159682: dataIn1 = 32'd5978
; 
32'd159683: dataIn1 = 32'd1105
; 
32'd159684: dataIn1 = 32'd4852
; 
32'd159685: dataIn1 = 32'd5958
; 
32'd159686: dataIn1 = 32'd5975
; 
32'd159687: dataIn1 = 32'd5977
; 
32'd159688: dataIn1 = 32'd7294
; 
32'd159689: dataIn1 = 32'd7326
; 
32'd159690: dataIn1 = 32'd2625
; 
32'd159691: dataIn1 = 32'd4852
; 
32'd159692: dataIn1 = 32'd5967
; 
32'd159693: dataIn1 = 32'd5976
; 
32'd159694: dataIn1 = 32'd5978
; 
32'd159695: dataIn1 = 32'd7325
; 
32'd159696: dataIn1 = 32'd7328
; 
32'd159697: dataIn1 = 32'd4662
; 
32'd159698: dataIn1 = 32'd4847
; 
32'd159699: dataIn1 = 32'd4850
; 
32'd159700: dataIn1 = 32'd5913
; 
32'd159701: dataIn1 = 32'd5965
; 
32'd159702: dataIn1 = 32'd5979
; 
32'd159703: dataIn1 = 32'd131
; 
32'd159704: dataIn1 = 32'd4621
; 
32'd159705: dataIn1 = 32'd4666
; 
32'd159706: dataIn1 = 32'd5922
; 
32'd159707: dataIn1 = 32'd5980
; 
32'd159708: dataIn1 = 32'd5981
; 
32'd159709: dataIn1 = 32'd5982
; 
32'd159710: dataIn1 = 32'd4666
; 
32'd159711: dataIn1 = 32'd4682
; 
32'd159712: dataIn1 = 32'd4854
; 
32'd159713: dataIn1 = 32'd5980
; 
32'd159714: dataIn1 = 32'd5981
; 
32'd159715: dataIn1 = 32'd5982
; 
32'd159716: dataIn1 = 32'd131
; 
32'd159717: dataIn1 = 32'd4635
; 
32'd159718: dataIn1 = 32'd4682
; 
32'd159719: dataIn1 = 32'd5980
; 
32'd159720: dataIn1 = 32'd5981
; 
32'd159721: dataIn1 = 32'd5982
; 
32'd159722: dataIn1 = 32'd6699
; 
32'd159723: dataIn1 = 32'd4857
; 
32'd159724: dataIn1 = 32'd4858
; 
32'd159725: dataIn1 = 32'd4859
; 
32'd159726: dataIn1 = 32'd5983
; 
32'd159727: dataIn1 = 32'd5984
; 
32'd159728: dataIn1 = 32'd5985
; 
32'd159729: dataIn1 = 32'd2626
; 
32'd159730: dataIn1 = 32'd4859
; 
32'd159731: dataIn1 = 32'd5983
; 
32'd159732: dataIn1 = 32'd5984
; 
32'd159733: dataIn1 = 32'd5985
; 
32'd159734: dataIn1 = 32'd5991
; 
32'd159735: dataIn1 = 32'd5994
; 
32'd159736: dataIn1 = 32'd2626
; 
32'd159737: dataIn1 = 32'd4858
; 
32'd159738: dataIn1 = 32'd5983
; 
32'd159739: dataIn1 = 32'd5984
; 
32'd159740: dataIn1 = 32'd5985
; 
32'd159741: dataIn1 = 32'd5986
; 
32'd159742: dataIn1 = 32'd5989
; 
32'd159743: dataIn1 = 32'd4858
; 
32'd159744: dataIn1 = 32'd4860
; 
32'd159745: dataIn1 = 32'd5985
; 
32'd159746: dataIn1 = 32'd5986
; 
32'd159747: dataIn1 = 32'd5987
; 
32'd159748: dataIn1 = 32'd5988
; 
32'd159749: dataIn1 = 32'd5989
; 
32'd159750: dataIn1 = 32'd4844
; 
32'd159751: dataIn1 = 32'd4860
; 
32'd159752: dataIn1 = 32'd5959
; 
32'd159753: dataIn1 = 32'd5986
; 
32'd159754: dataIn1 = 32'd5987
; 
32'd159755: dataIn1 = 32'd5988
; 
32'd159756: dataIn1 = 32'd5990
; 
32'd159757: dataIn1 = 32'd2624
; 
32'd159758: dataIn1 = 32'd4844
; 
32'd159759: dataIn1 = 32'd4858
; 
32'd159760: dataIn1 = 32'd5986
; 
32'd159761: dataIn1 = 32'd5987
; 
32'd159762: dataIn1 = 32'd5988
; 
32'd159763: dataIn1 = 32'd2626
; 
32'd159764: dataIn1 = 32'd4860
; 
32'd159765: dataIn1 = 32'd5985
; 
32'd159766: dataIn1 = 32'd5986
; 
32'd159767: dataIn1 = 32'd5989
; 
32'd159768: dataIn1 = 32'd7341
; 
32'd159769: dataIn1 = 32'd7345
; 
32'd159770: dataIn1 = 32'd1105
; 
32'd159771: dataIn1 = 32'd4860
; 
32'd159772: dataIn1 = 32'd5959
; 
32'd159773: dataIn1 = 32'd5987
; 
32'd159774: dataIn1 = 32'd5990
; 
32'd159775: dataIn1 = 32'd7295
; 
32'd159776: dataIn1 = 32'd7344
; 
32'd159777: dataIn1 = 32'd4859
; 
32'd159778: dataIn1 = 32'd4861
; 
32'd159779: dataIn1 = 32'd5984
; 
32'd159780: dataIn1 = 32'd5991
; 
32'd159781: dataIn1 = 32'd5992
; 
32'd159782: dataIn1 = 32'd5993
; 
32'd159783: dataIn1 = 32'd5994
; 
32'd159784: dataIn1 = 32'd2569
; 
32'd159785: dataIn1 = 32'd4678
; 
32'd159786: dataIn1 = 32'd4859
; 
32'd159787: dataIn1 = 32'd5991
; 
32'd159788: dataIn1 = 32'd5992
; 
32'd159789: dataIn1 = 32'd5993
; 
32'd159790: dataIn1 = 32'd4678
; 
32'd159791: dataIn1 = 32'd4861
; 
32'd159792: dataIn1 = 32'd5940
; 
32'd159793: dataIn1 = 32'd5991
; 
32'd159794: dataIn1 = 32'd5992
; 
32'd159795: dataIn1 = 32'd5993
; 
32'd159796: dataIn1 = 32'd5995
; 
32'd159797: dataIn1 = 32'd2626
; 
32'd159798: dataIn1 = 32'd4861
; 
32'd159799: dataIn1 = 32'd5984
; 
32'd159800: dataIn1 = 32'd5991
; 
32'd159801: dataIn1 = 32'd5994
; 
32'd159802: dataIn1 = 32'd7340
; 
32'd159803: dataIn1 = 32'd7353
; 
32'd159804: dataIn1 = 32'd6
; 
32'd159805: dataIn1 = 32'd4861
; 
32'd159806: dataIn1 = 32'd5940
; 
32'd159807: dataIn1 = 32'd5993
; 
32'd159808: dataIn1 = 32'd5995
; 
32'd159809: dataIn1 = 32'd7354
; 
32'd159810: dataIn1 = 32'd8963
; 
32'd159811: dataIn1 = 32'd4863
; 
32'd159812: dataIn1 = 32'd4864
; 
32'd159813: dataIn1 = 32'd5996
; 
32'd159814: dataIn1 = 32'd5997
; 
32'd159815: dataIn1 = 32'd5998
; 
32'd159816: dataIn1 = 32'd5999
; 
32'd159817: dataIn1 = 32'd6000
; 
32'd159818: dataIn1 = 32'd4862
; 
32'd159819: dataIn1 = 32'd4864
; 
32'd159820: dataIn1 = 32'd5996
; 
32'd159821: dataIn1 = 32'd5997
; 
32'd159822: dataIn1 = 32'd5998
; 
32'd159823: dataIn1 = 32'd6001
; 
32'd159824: dataIn1 = 32'd6002
; 
32'd159825: dataIn1 = 32'd4862
; 
32'd159826: dataIn1 = 32'd4863
; 
32'd159827: dataIn1 = 32'd5996
; 
32'd159828: dataIn1 = 32'd5997
; 
32'd159829: dataIn1 = 32'd5998
; 
32'd159830: dataIn1 = 32'd6003
; 
32'd159831: dataIn1 = 32'd6004
; 
32'd159832: dataIn1 = 32'd2627
; 
32'd159833: dataIn1 = 32'd4864
; 
32'd159834: dataIn1 = 32'd5996
; 
32'd159835: dataIn1 = 32'd5999
; 
32'd159836: dataIn1 = 32'd6000
; 
32'd159837: dataIn1 = 32'd6014
; 
32'd159838: dataIn1 = 32'd6017
; 
32'd159839: dataIn1 = 32'd2627
; 
32'd159840: dataIn1 = 32'd4863
; 
32'd159841: dataIn1 = 32'd5996
; 
32'd159842: dataIn1 = 32'd5999
; 
32'd159843: dataIn1 = 32'd6000
; 
32'd159844: dataIn1 = 32'd6009
; 
32'd159845: dataIn1 = 32'd6012
; 
32'd159846: dataIn1 = 32'd2628
; 
32'd159847: dataIn1 = 32'd4864
; 
32'd159848: dataIn1 = 32'd5997
; 
32'd159849: dataIn1 = 32'd6001
; 
32'd159850: dataIn1 = 32'd6002
; 
32'd159851: dataIn1 = 32'd6015
; 
32'd159852: dataIn1 = 32'd6018
; 
32'd159853: dataIn1 = 32'd2628
; 
32'd159854: dataIn1 = 32'd4862
; 
32'd159855: dataIn1 = 32'd5997
; 
32'd159856: dataIn1 = 32'd6001
; 
32'd159857: dataIn1 = 32'd6002
; 
32'd159858: dataIn1 = 32'd6005
; 
32'd159859: dataIn1 = 32'd6006
; 
32'd159860: dataIn1 = 32'd2629
; 
32'd159861: dataIn1 = 32'd4863
; 
32'd159862: dataIn1 = 32'd5998
; 
32'd159863: dataIn1 = 32'd6003
; 
32'd159864: dataIn1 = 32'd6004
; 
32'd159865: dataIn1 = 32'd6011
; 
32'd159866: dataIn1 = 32'd6013
; 
32'd159867: dataIn1 = 32'd2629
; 
32'd159868: dataIn1 = 32'd4862
; 
32'd159869: dataIn1 = 32'd5998
; 
32'd159870: dataIn1 = 32'd6003
; 
32'd159871: dataIn1 = 32'd6004
; 
32'd159872: dataIn1 = 32'd6007
; 
32'd159873: dataIn1 = 32'd6008
; 
32'd159874: dataIn1 = 32'd2628
; 
32'd159875: dataIn1 = 32'd4866
; 
32'd159876: dataIn1 = 32'd6002
; 
32'd159877: dataIn1 = 32'd6005
; 
32'd159878: dataIn1 = 32'd6006
; 
32'd159879: dataIn1 = 32'd6048
; 
32'd159880: dataIn1 = 32'd6701
; 
32'd159881: dataIn1 = 32'd4862
; 
32'd159882: dataIn1 = 32'd4866
; 
32'd159883: dataIn1 = 32'd6002
; 
32'd159884: dataIn1 = 32'd6005
; 
32'd159885: dataIn1 = 32'd6006
; 
32'd159886: dataIn1 = 32'd6008
; 
32'd159887: dataIn1 = 32'd6700
; 
32'd159888: dataIn1 = 32'd2629
; 
32'd159889: dataIn1 = 32'd4865
; 
32'd159890: dataIn1 = 32'd4881
; 
32'd159891: dataIn1 = 32'd6004
; 
32'd159892: dataIn1 = 32'd6007
; 
32'd159893: dataIn1 = 32'd6008
; 
32'd159894: dataIn1 = 32'd4862
; 
32'd159895: dataIn1 = 32'd4865
; 
32'd159896: dataIn1 = 32'd6004
; 
32'd159897: dataIn1 = 32'd6006
; 
32'd159898: dataIn1 = 32'd6007
; 
32'd159899: dataIn1 = 32'd6008
; 
32'd159900: dataIn1 = 32'd6700
; 
32'd159901: dataIn1 = 32'd4863
; 
32'd159902: dataIn1 = 32'd4868
; 
32'd159903: dataIn1 = 32'd6000
; 
32'd159904: dataIn1 = 32'd6009
; 
32'd159905: dataIn1 = 32'd6010
; 
32'd159906: dataIn1 = 32'd6011
; 
32'd159907: dataIn1 = 32'd6012
; 
32'd159908: dataIn1 = 32'd4867
; 
32'd159909: dataIn1 = 32'd4868
; 
32'd159910: dataIn1 = 32'd6009
; 
32'd159911: dataIn1 = 32'd6010
; 
32'd159912: dataIn1 = 32'd6011
; 
32'd159913: dataIn1 = 32'd6697
; 
32'd159914: dataIn1 = 32'd6702
; 
32'd159915: dataIn1 = 32'd4863
; 
32'd159916: dataIn1 = 32'd4867
; 
32'd159917: dataIn1 = 32'd6003
; 
32'd159918: dataIn1 = 32'd6009
; 
32'd159919: dataIn1 = 32'd6010
; 
32'd159920: dataIn1 = 32'd6011
; 
32'd159921: dataIn1 = 32'd6013
; 
32'd159922: dataIn1 = 32'd2627
; 
32'd159923: dataIn1 = 32'd4868
; 
32'd159924: dataIn1 = 32'd6000
; 
32'd159925: dataIn1 = 32'd6009
; 
32'd159926: dataIn1 = 32'd6012
; 
32'd159927: dataIn1 = 32'd6025
; 
32'd159928: dataIn1 = 32'd6035
; 
32'd159929: dataIn1 = 32'd2629
; 
32'd159930: dataIn1 = 32'd4867
; 
32'd159931: dataIn1 = 32'd4882
; 
32'd159932: dataIn1 = 32'd6003
; 
32'd159933: dataIn1 = 32'd6011
; 
32'd159934: dataIn1 = 32'd6013
; 
32'd159935: dataIn1 = 32'd4864
; 
32'd159936: dataIn1 = 32'd4870
; 
32'd159937: dataIn1 = 32'd5999
; 
32'd159938: dataIn1 = 32'd6014
; 
32'd159939: dataIn1 = 32'd6015
; 
32'd159940: dataIn1 = 32'd6016
; 
32'd159941: dataIn1 = 32'd6017
; 
32'd159942: dataIn1 = 32'd4864
; 
32'd159943: dataIn1 = 32'd4869
; 
32'd159944: dataIn1 = 32'd6001
; 
32'd159945: dataIn1 = 32'd6014
; 
32'd159946: dataIn1 = 32'd6015
; 
32'd159947: dataIn1 = 32'd6016
; 
32'd159948: dataIn1 = 32'd6018
; 
32'd159949: dataIn1 = 32'd4869
; 
32'd159950: dataIn1 = 32'd4870
; 
32'd159951: dataIn1 = 32'd6014
; 
32'd159952: dataIn1 = 32'd6015
; 
32'd159953: dataIn1 = 32'd6016
; 
32'd159954: dataIn1 = 32'd6019
; 
32'd159955: dataIn1 = 32'd6020
; 
32'd159956: dataIn1 = 32'd2627
; 
32'd159957: dataIn1 = 32'd4870
; 
32'd159958: dataIn1 = 32'd5999
; 
32'd159959: dataIn1 = 32'd6014
; 
32'd159960: dataIn1 = 32'd6017
; 
32'd159961: dataIn1 = 32'd6024
; 
32'd159962: dataIn1 = 32'd6038
; 
32'd159963: dataIn1 = 32'd2628
; 
32'd159964: dataIn1 = 32'd4869
; 
32'd159965: dataIn1 = 32'd6001
; 
32'd159966: dataIn1 = 32'd6015
; 
32'd159967: dataIn1 = 32'd6018
; 
32'd159968: dataIn1 = 32'd6046
; 
32'd159969: dataIn1 = 32'd6057
; 
32'd159970: dataIn1 = 32'd1106
; 
32'd159971: dataIn1 = 32'd4870
; 
32'd159972: dataIn1 = 32'd6016
; 
32'd159973: dataIn1 = 32'd6019
; 
32'd159974: dataIn1 = 32'd6020
; 
32'd159975: dataIn1 = 32'd6040
; 
32'd159976: dataIn1 = 32'd6042
; 
32'd159977: dataIn1 = 32'd1106
; 
32'd159978: dataIn1 = 32'd4869
; 
32'd159979: dataIn1 = 32'd6016
; 
32'd159980: dataIn1 = 32'd6019
; 
32'd159981: dataIn1 = 32'd6020
; 
32'd159982: dataIn1 = 32'd6058
; 
32'd159983: dataIn1 = 32'd6060
; 
32'd159984: dataIn1 = 32'd4872
; 
32'd159985: dataIn1 = 32'd4873
; 
32'd159986: dataIn1 = 32'd6021
; 
32'd159987: dataIn1 = 32'd6022
; 
32'd159988: dataIn1 = 32'd6023
; 
32'd159989: dataIn1 = 32'd6024
; 
32'd159990: dataIn1 = 32'd6025
; 
32'd159991: dataIn1 = 32'd4871
; 
32'd159992: dataIn1 = 32'd4873
; 
32'd159993: dataIn1 = 32'd6021
; 
32'd159994: dataIn1 = 32'd6022
; 
32'd159995: dataIn1 = 32'd6023
; 
32'd159996: dataIn1 = 32'd6026
; 
32'd159997: dataIn1 = 32'd6027
; 
32'd159998: dataIn1 = 32'd4871
; 
32'd159999: dataIn1 = 32'd4872
; 
32'd160000: dataIn1 = 32'd6021
; 
32'd160001: dataIn1 = 32'd6022
; 
32'd160002: dataIn1 = 32'd6023
; 
32'd160003: dataIn1 = 32'd6028
; 
32'd160004: dataIn1 = 32'd6029
; 
32'd160005: dataIn1 = 32'd2627
; 
32'd160006: dataIn1 = 32'd4873
; 
32'd160007: dataIn1 = 32'd6017
; 
32'd160008: dataIn1 = 32'd6021
; 
32'd160009: dataIn1 = 32'd6024
; 
32'd160010: dataIn1 = 32'd6025
; 
32'd160011: dataIn1 = 32'd6038
; 
32'd160012: dataIn1 = 32'd2627
; 
32'd160013: dataIn1 = 32'd4872
; 
32'd160014: dataIn1 = 32'd6012
; 
32'd160015: dataIn1 = 32'd6021
; 
32'd160016: dataIn1 = 32'd6024
; 
32'd160017: dataIn1 = 32'd6025
; 
32'd160018: dataIn1 = 32'd6035
; 
32'd160019: dataIn1 = 32'd2630
; 
32'd160020: dataIn1 = 32'd4873
; 
32'd160021: dataIn1 = 32'd6022
; 
32'd160022: dataIn1 = 32'd6026
; 
32'd160023: dataIn1 = 32'd6027
; 
32'd160024: dataIn1 = 32'd6039
; 
32'd160025: dataIn1 = 32'd6041
; 
32'd160026: dataIn1 = 32'd2630
; 
32'd160027: dataIn1 = 32'd4871
; 
32'd160028: dataIn1 = 32'd6022
; 
32'd160029: dataIn1 = 32'd6026
; 
32'd160030: dataIn1 = 32'd6027
; 
32'd160031: dataIn1 = 32'd6031
; 
32'd160032: dataIn1 = 32'd6034
; 
32'd160033: dataIn1 = 32'd2562
; 
32'd160034: dataIn1 = 32'd4872
; 
32'd160035: dataIn1 = 32'd5911
; 
32'd160036: dataIn1 = 32'd6023
; 
32'd160037: dataIn1 = 32'd6028
; 
32'd160038: dataIn1 = 32'd6029
; 
32'd160039: dataIn1 = 32'd6037
; 
32'd160040: dataIn1 = 32'd2562
; 
32'd160041: dataIn1 = 32'd4871
; 
32'd160042: dataIn1 = 32'd5905
; 
32'd160043: dataIn1 = 32'd6023
; 
32'd160044: dataIn1 = 32'd6028
; 
32'd160045: dataIn1 = 32'd6029
; 
32'd160046: dataIn1 = 32'd6032
; 
32'd160047: dataIn1 = 32'd4659
; 
32'd160048: dataIn1 = 32'd4874
; 
32'd160049: dataIn1 = 32'd5903
; 
32'd160050: dataIn1 = 32'd6030
; 
32'd160051: dataIn1 = 32'd6031
; 
32'd160052: dataIn1 = 32'd6032
; 
32'd160053: dataIn1 = 32'd6033
; 
32'd160054: dataIn1 = 32'd4871
; 
32'd160055: dataIn1 = 32'd4874
; 
32'd160056: dataIn1 = 32'd6027
; 
32'd160057: dataIn1 = 32'd6030
; 
32'd160058: dataIn1 = 32'd6031
; 
32'd160059: dataIn1 = 32'd6032
; 
32'd160060: dataIn1 = 32'd6034
; 
32'd160061: dataIn1 = 32'd4659
; 
32'd160062: dataIn1 = 32'd4871
; 
32'd160063: dataIn1 = 32'd5905
; 
32'd160064: dataIn1 = 32'd6029
; 
32'd160065: dataIn1 = 32'd6030
; 
32'd160066: dataIn1 = 32'd6031
; 
32'd160067: dataIn1 = 32'd6032
; 
32'd160068: dataIn1 = 32'd130
; 
32'd160069: dataIn1 = 32'd4874
; 
32'd160070: dataIn1 = 32'd5903
; 
32'd160071: dataIn1 = 32'd6030
; 
32'd160072: dataIn1 = 32'd6033
; 
32'd160073: dataIn1 = 32'd7238
; 
32'd160074: dataIn1 = 32'd7277
; 
32'd160075: dataIn1 = 32'd2630
; 
32'd160076: dataIn1 = 32'd4874
; 
32'd160077: dataIn1 = 32'd6027
; 
32'd160078: dataIn1 = 32'd6031
; 
32'd160079: dataIn1 = 32'd6034
; 
32'd160080: dataIn1 = 32'd7267
; 
32'd160081: dataIn1 = 32'd7276
; 
32'd160082: dataIn1 = 32'd4868
; 
32'd160083: dataIn1 = 32'd4872
; 
32'd160084: dataIn1 = 32'd6012
; 
32'd160085: dataIn1 = 32'd6025
; 
32'd160086: dataIn1 = 32'd6035
; 
32'd160087: dataIn1 = 32'd6036
; 
32'd160088: dataIn1 = 32'd6037
; 
32'd160089: dataIn1 = 32'd4661
; 
32'd160090: dataIn1 = 32'd4868
; 
32'd160091: dataIn1 = 32'd5910
; 
32'd160092: dataIn1 = 32'd6035
; 
32'd160093: dataIn1 = 32'd6036
; 
32'd160094: dataIn1 = 32'd6037
; 
32'd160095: dataIn1 = 32'd6697
; 
32'd160096: dataIn1 = 32'd4661
; 
32'd160097: dataIn1 = 32'd4872
; 
32'd160098: dataIn1 = 32'd5911
; 
32'd160099: dataIn1 = 32'd6028
; 
32'd160100: dataIn1 = 32'd6035
; 
32'd160101: dataIn1 = 32'd6036
; 
32'd160102: dataIn1 = 32'd6037
; 
32'd160103: dataIn1 = 32'd4870
; 
32'd160104: dataIn1 = 32'd4873
; 
32'd160105: dataIn1 = 32'd6017
; 
32'd160106: dataIn1 = 32'd6024
; 
32'd160107: dataIn1 = 32'd6038
; 
32'd160108: dataIn1 = 32'd6039
; 
32'd160109: dataIn1 = 32'd6040
; 
32'd160110: dataIn1 = 32'd4873
; 
32'd160111: dataIn1 = 32'd4875
; 
32'd160112: dataIn1 = 32'd6026
; 
32'd160113: dataIn1 = 32'd6038
; 
32'd160114: dataIn1 = 32'd6039
; 
32'd160115: dataIn1 = 32'd6040
; 
32'd160116: dataIn1 = 32'd6041
; 
32'd160117: dataIn1 = 32'd4870
; 
32'd160118: dataIn1 = 32'd4875
; 
32'd160119: dataIn1 = 32'd6019
; 
32'd160120: dataIn1 = 32'd6038
; 
32'd160121: dataIn1 = 32'd6039
; 
32'd160122: dataIn1 = 32'd6040
; 
32'd160123: dataIn1 = 32'd6042
; 
32'd160124: dataIn1 = 32'd2630
; 
32'd160125: dataIn1 = 32'd4875
; 
32'd160126: dataIn1 = 32'd6026
; 
32'd160127: dataIn1 = 32'd6039
; 
32'd160128: dataIn1 = 32'd6041
; 
32'd160129: dataIn1 = 32'd7266
; 
32'd160130: dataIn1 = 32'd7279
; 
32'd160131: dataIn1 = 32'd1106
; 
32'd160132: dataIn1 = 32'd4875
; 
32'd160133: dataIn1 = 32'd6019
; 
32'd160134: dataIn1 = 32'd6040
; 
32'd160135: dataIn1 = 32'd6042
; 
32'd160136: dataIn1 = 32'd7255
; 
32'd160137: dataIn1 = 32'd7281
; 
32'd160138: dataIn1 = 32'd4877
; 
32'd160139: dataIn1 = 32'd4878
; 
32'd160140: dataIn1 = 32'd6043
; 
32'd160141: dataIn1 = 32'd6044
; 
32'd160142: dataIn1 = 32'd6045
; 
32'd160143: dataIn1 = 32'd6047
; 
32'd160144: dataIn1 = 32'd6051
; 
32'd160145: dataIn1 = 32'd2631
; 
32'd160146: dataIn1 = 32'd4878
; 
32'd160147: dataIn1 = 32'd6043
; 
32'd160148: dataIn1 = 32'd6044
; 
32'd160149: dataIn1 = 32'd6045
; 
32'd160150: dataIn1 = 32'd6056
; 
32'd160151: dataIn1 = 32'd6059
; 
32'd160152: dataIn1 = 32'd2631
; 
32'd160153: dataIn1 = 32'd4877
; 
32'd160154: dataIn1 = 32'd6043
; 
32'd160155: dataIn1 = 32'd6044
; 
32'd160156: dataIn1 = 32'd6045
; 
32'd160157: dataIn1 = 32'd6052
; 
32'd160158: dataIn1 = 32'd6703
; 
32'd160159: dataIn1 = 32'd2628
; 
32'd160160: dataIn1 = 32'd4878
; 
32'd160161: dataIn1 = 32'd6018
; 
32'd160162: dataIn1 = 32'd6046
; 
32'd160163: dataIn1 = 32'd6047
; 
32'd160164: dataIn1 = 32'd6048
; 
32'd160165: dataIn1 = 32'd6057
; 
32'd160166: dataIn1 = 32'd4876
; 
32'd160167: dataIn1 = 32'd4878
; 
32'd160168: dataIn1 = 32'd6043
; 
32'd160169: dataIn1 = 32'd6046
; 
32'd160170: dataIn1 = 32'd6047
; 
32'd160171: dataIn1 = 32'd6048
; 
32'd160172: dataIn1 = 32'd6051
; 
32'd160173: dataIn1 = 32'd2628
; 
32'd160174: dataIn1 = 32'd4876
; 
32'd160175: dataIn1 = 32'd6005
; 
32'd160176: dataIn1 = 32'd6046
; 
32'd160177: dataIn1 = 32'd6047
; 
32'd160178: dataIn1 = 32'd6048
; 
32'd160179: dataIn1 = 32'd6701
; 
32'd160180: dataIn1 = 32'd2307
; 
32'd160181: dataIn1 = 32'd4877
; 
32'd160182: dataIn1 = 32'd5739
; 
32'd160183: dataIn1 = 32'd6049
; 
32'd160184: dataIn1 = 32'd6050
; 
32'd160185: dataIn1 = 32'd6051
; 
32'd160186: dataIn1 = 32'd6054
; 
32'd160187: dataIn1 = 32'd2307
; 
32'd160188: dataIn1 = 32'd4876
; 
32'd160189: dataIn1 = 32'd5744
; 
32'd160190: dataIn1 = 32'd6049
; 
32'd160191: dataIn1 = 32'd6050
; 
32'd160192: dataIn1 = 32'd6051
; 
32'd160193: dataIn1 = 32'd6696
; 
32'd160194: dataIn1 = 32'd4876
; 
32'd160195: dataIn1 = 32'd4877
; 
32'd160196: dataIn1 = 32'd6043
; 
32'd160197: dataIn1 = 32'd6047
; 
32'd160198: dataIn1 = 32'd6049
; 
32'd160199: dataIn1 = 32'd6050
; 
32'd160200: dataIn1 = 32'd6051
; 
32'd160201: dataIn1 = 32'd4877
; 
32'd160202: dataIn1 = 32'd4879
; 
32'd160203: dataIn1 = 32'd6045
; 
32'd160204: dataIn1 = 32'd6052
; 
32'd160205: dataIn1 = 32'd6053
; 
32'd160206: dataIn1 = 32'd6054
; 
32'd160207: dataIn1 = 32'd6703
; 
32'd160208: dataIn1 = 32'd3919
; 
32'd160209: dataIn1 = 32'd4879
; 
32'd160210: dataIn1 = 32'd5740
; 
32'd160211: dataIn1 = 32'd6052
; 
32'd160212: dataIn1 = 32'd6053
; 
32'd160213: dataIn1 = 32'd6054
; 
32'd160214: dataIn1 = 32'd6055
; 
32'd160215: dataIn1 = 32'd3919
; 
32'd160216: dataIn1 = 32'd4877
; 
32'd160217: dataIn1 = 32'd5739
; 
32'd160218: dataIn1 = 32'd6049
; 
32'd160219: dataIn1 = 32'd6052
; 
32'd160220: dataIn1 = 32'd6053
; 
32'd160221: dataIn1 = 32'd6054
; 
32'd160222: dataIn1 = 32'd5
; 
32'd160223: dataIn1 = 32'd4879
; 
32'd160224: dataIn1 = 32'd5740
; 
32'd160225: dataIn1 = 32'd6053
; 
32'd160226: dataIn1 = 32'd6055
; 
32'd160227: dataIn1 = 32'd7256
; 
32'd160228: dataIn1 = 32'd8924
; 
32'd160229: dataIn1 = 32'd4878
; 
32'd160230: dataIn1 = 32'd4880
; 
32'd160231: dataIn1 = 32'd6044
; 
32'd160232: dataIn1 = 32'd6056
; 
32'd160233: dataIn1 = 32'd6057
; 
32'd160234: dataIn1 = 32'd6058
; 
32'd160235: dataIn1 = 32'd6059
; 
32'd160236: dataIn1 = 32'd4869
; 
32'd160237: dataIn1 = 32'd4878
; 
32'd160238: dataIn1 = 32'd6018
; 
32'd160239: dataIn1 = 32'd6046
; 
32'd160240: dataIn1 = 32'd6056
; 
32'd160241: dataIn1 = 32'd6057
; 
32'd160242: dataIn1 = 32'd6058
; 
32'd160243: dataIn1 = 32'd4869
; 
32'd160244: dataIn1 = 32'd4880
; 
32'd160245: dataIn1 = 32'd6020
; 
32'd160246: dataIn1 = 32'd6056
; 
32'd160247: dataIn1 = 32'd6057
; 
32'd160248: dataIn1 = 32'd6058
; 
32'd160249: dataIn1 = 32'd6060
; 
32'd160250: dataIn1 = 32'd2631
; 
32'd160251: dataIn1 = 32'd4880
; 
32'd160252: dataIn1 = 32'd6044
; 
32'd160253: dataIn1 = 32'd6056
; 
32'd160254: dataIn1 = 32'd6059
; 
32'd160255: dataIn1 = 32'd7260
; 
32'd160256: dataIn1 = 32'd9274
; 
32'd160257: dataIn1 = 32'd1106
; 
32'd160258: dataIn1 = 32'd4880
; 
32'd160259: dataIn1 = 32'd6020
; 
32'd160260: dataIn1 = 32'd6058
; 
32'd160261: dataIn1 = 32'd6060
; 
32'd160262: dataIn1 = 32'd7254
; 
32'd160263: dataIn1 = 32'd7261
; 
32'd160264: dataIn1 = 32'd2564
; 
32'd160265: dataIn1 = 32'd4672
; 
32'd160266: dataIn1 = 32'd4883
; 
32'd160267: dataIn1 = 32'd6061
; 
32'd160268: dataIn1 = 32'd6062
; 
32'd160269: dataIn1 = 32'd6063
; 
32'd160270: dataIn1 = 32'd3912
; 
32'd160271: dataIn1 = 32'd4883
; 
32'd160272: dataIn1 = 32'd5723
; 
32'd160273: dataIn1 = 32'd6061
; 
32'd160274: dataIn1 = 32'd6062
; 
32'd160275: dataIn1 = 32'd6063
; 
32'd160276: dataIn1 = 32'd6064
; 
32'd160277: dataIn1 = 32'd3912
; 
32'd160278: dataIn1 = 32'd4672
; 
32'd160279: dataIn1 = 32'd5721
; 
32'd160280: dataIn1 = 32'd5936
; 
32'd160281: dataIn1 = 32'd6061
; 
32'd160282: dataIn1 = 32'd6062
; 
32'd160283: dataIn1 = 32'd6063
; 
32'd160284: dataIn1 = 32'd2306
; 
32'd160285: dataIn1 = 32'd4881
; 
32'd160286: dataIn1 = 32'd4883
; 
32'd160287: dataIn1 = 32'd5723
; 
32'd160288: dataIn1 = 32'd6062
; 
32'd160289: dataIn1 = 32'd6064
; 
32'd160290: dataIn1 = 32'd6
; 
32'd160291: dataIn1 = 32'd4901
; 
32'd160292: dataIn1 = 32'd5938
; 
32'd160293: dataIn1 = 32'd6065
; 
32'd160294: dataIn1 = 32'd6066
; 
32'd160295: dataIn1 = 32'd7458
; 
32'd160296: dataIn1 = 32'd8962
; 
32'd160297: dataIn1 = 32'd4679
; 
32'd160298: dataIn1 = 32'd4899
; 
32'd160299: dataIn1 = 32'd4901
; 
32'd160300: dataIn1 = 32'd5938
; 
32'd160301: dataIn1 = 32'd6065
; 
32'd160302: dataIn1 = 32'd6066
; 
32'd160303: dataIn1 = 32'd6067
; 
32'd160304: dataIn1 = 32'd7056
; 
32'd160305: dataIn1 = 32'd7057
; 
32'd160306: dataIn1 = 32'd7061
; 
32'd160307: dataIn1 = 32'd7063
; 
32'd160308: dataIn1 = 32'd7065
; 
32'd160309: dataIn1 = 32'd7066
; 
32'd160310: dataIn1 = 32'd6068
; 
32'd160311: dataIn1 = 32'd6072
; 
32'd160312: dataIn1 = 32'd6073
; 
32'd160313: dataIn1 = 32'd7055
; 
32'd160314: dataIn1 = 32'd7057
; 
32'd160315: dataIn1 = 32'd7059
; 
32'd160316: dataIn1 = 32'd7062
; 
32'd160317: dataIn1 = 32'd6069
; 
32'd160318: dataIn1 = 32'd7055
; 
32'd160319: dataIn1 = 32'd7056
; 
32'd160320: dataIn1 = 32'd7058
; 
32'd160321: dataIn1 = 32'd7060
; 
32'd160322: dataIn1 = 32'd7071
; 
32'd160323: dataIn1 = 32'd7072
; 
32'd160324: dataIn1 = 32'd6070
; 
32'd160325: dataIn1 = 32'd7064
; 
32'd160326: dataIn1 = 32'd7066
; 
32'd160327: dataIn1 = 32'd7068
; 
32'd160328: dataIn1 = 32'd7070
; 
32'd160329: dataIn1 = 32'd7104
; 
32'd160330: dataIn1 = 32'd7106
; 
32'd160331: dataIn1 = 32'd6071
; 
32'd160332: dataIn1 = 32'd7064
; 
32'd160333: dataIn1 = 32'd7065
; 
32'd160334: dataIn1 = 32'd7067
; 
32'd160335: dataIn1 = 32'd7069
; 
32'd160336: dataIn1 = 32'd7094
; 
32'd160337: dataIn1 = 32'd7095
; 
32'd160338: dataIn1 = 32'd2693
; 
32'd160339: dataIn1 = 32'd5114
; 
32'd160340: dataIn1 = 32'd6068
; 
32'd160341: dataIn1 = 32'd6072
; 
32'd160342: dataIn1 = 32'd6073
; 
32'd160343: dataIn1 = 32'd6091
; 
32'd160344: dataIn1 = 32'd6094
; 
32'd160345: dataIn1 = 32'd7062
; 
32'd160346: dataIn1 = 32'd2693
; 
32'd160347: dataIn1 = 32'd5112
; 
32'd160348: dataIn1 = 32'd6068
; 
32'd160349: dataIn1 = 32'd6072
; 
32'd160350: dataIn1 = 32'd6073
; 
32'd160351: dataIn1 = 32'd6077
; 
32'd160352: dataIn1 = 32'd6081
; 
32'd160353: dataIn1 = 32'd7059
; 
32'd160354: dataIn1 = 32'd6074
; 
32'd160355: dataIn1 = 32'd7072
; 
32'd160356: dataIn1 = 32'd7073
; 
32'd160357: dataIn1 = 32'd7075
; 
32'd160358: dataIn1 = 32'd7077
; 
32'd160359: dataIn1 = 32'd7100
; 
32'd160360: dataIn1 = 32'd7101
; 
32'd160361: dataIn1 = 32'd6075
; 
32'd160362: dataIn1 = 32'd7071
; 
32'd160363: dataIn1 = 32'd7073
; 
32'd160364: dataIn1 = 32'd7074
; 
32'd160365: dataIn1 = 32'd7076
; 
32'd160366: dataIn1 = 32'd7078
; 
32'd160367: dataIn1 = 32'd7080
; 
32'd160368: dataIn1 = 32'd5115
; 
32'd160369: dataIn1 = 32'd5116
; 
32'd160370: dataIn1 = 32'd6076
; 
32'd160371: dataIn1 = 32'd6077
; 
32'd160372: dataIn1 = 32'd6078
; 
32'd160373: dataIn1 = 32'd6079
; 
32'd160374: dataIn1 = 32'd6080
; 
32'd160375: dataIn1 = 32'd7082
; 
32'd160376: dataIn1 = 32'd5112
; 
32'd160377: dataIn1 = 32'd5116
; 
32'd160378: dataIn1 = 32'd6073
; 
32'd160379: dataIn1 = 32'd6076
; 
32'd160380: dataIn1 = 32'd6077
; 
32'd160381: dataIn1 = 32'd6078
; 
32'd160382: dataIn1 = 32'd6081
; 
32'd160383: dataIn1 = 32'd7081
; 
32'd160384: dataIn1 = 32'd6076
; 
32'd160385: dataIn1 = 32'd6077
; 
32'd160386: dataIn1 = 32'd6078
; 
32'd160387: dataIn1 = 32'd7078
; 
32'd160388: dataIn1 = 32'd7079
; 
32'd160389: dataIn1 = 32'd7081
; 
32'd160390: dataIn1 = 32'd7082
; 
32'd160391: dataIn1 = 32'd1119
; 
32'd160392: dataIn1 = 32'd5116
; 
32'd160393: dataIn1 = 32'd6076
; 
32'd160394: dataIn1 = 32'd6079
; 
32'd160395: dataIn1 = 32'd6080
; 
32'd160396: dataIn1 = 32'd6705
; 
32'd160397: dataIn1 = 32'd1119
; 
32'd160398: dataIn1 = 32'd5115
; 
32'd160399: dataIn1 = 32'd6076
; 
32'd160400: dataIn1 = 32'd6079
; 
32'd160401: dataIn1 = 32'd6080
; 
32'd160402: dataIn1 = 32'd6128
; 
32'd160403: dataIn1 = 32'd6131
; 
32'd160404: dataIn1 = 32'd7192
; 
32'd160405: dataIn1 = 32'd2693
; 
32'd160406: dataIn1 = 32'd5116
; 
32'd160407: dataIn1 = 32'd6073
; 
32'd160408: dataIn1 = 32'd6077
; 
32'd160409: dataIn1 = 32'd6081
; 
32'd160410: dataIn1 = 32'd6704
; 
32'd160411: dataIn1 = 32'd6082
; 
32'd160412: dataIn1 = 32'd7079
; 
32'd160413: dataIn1 = 32'd7080
; 
32'd160414: dataIn1 = 32'd7083
; 
32'd160415: dataIn1 = 32'd7084
; 
32'd160416: dataIn1 = 32'd7201
; 
32'd160417: dataIn1 = 32'd7202
; 
32'd160418: dataIn1 = 32'd6083
; 
32'd160419: dataIn1 = 32'd7086
; 
32'd160420: dataIn1 = 32'd7087
; 
32'd160421: dataIn1 = 32'd7091
; 
32'd160422: dataIn1 = 32'd7093
; 
32'd160423: dataIn1 = 32'd7095
; 
32'd160424: dataIn1 = 32'd7096
; 
32'd160425: dataIn1 = 32'd6084
; 
32'd160426: dataIn1 = 32'd7085
; 
32'd160427: dataIn1 = 32'd7087
; 
32'd160428: dataIn1 = 32'd7089
; 
32'd160429: dataIn1 = 32'd7092
; 
32'd160430: dataIn1 = 32'd9792
; 
32'd160431: dataIn1 = 32'd9793
; 
32'd160432: dataIn1 = 32'd6085
; 
32'd160433: dataIn1 = 32'd7085
; 
32'd160434: dataIn1 = 32'd7086
; 
32'd160435: dataIn1 = 32'd7088
; 
32'd160436: dataIn1 = 32'd7090
; 
32'd160437: dataIn1 = 32'd7099
; 
32'd160438: dataIn1 = 32'd7100
; 
32'd160439: dataIn1 = 32'd6086
; 
32'd160440: dataIn1 = 32'd7094
; 
32'd160441: dataIn1 = 32'd7096
; 
32'd160442: dataIn1 = 32'd7097
; 
32'd160443: dataIn1 = 32'd7098
; 
32'd160444: dataIn1 = 32'd7141
; 
32'd160445: dataIn1 = 32'd7143
; 
32'd160446: dataIn1 = 32'd6087
; 
32'd160447: dataIn1 = 32'd9678
; 
32'd160448: dataIn1 = 32'd9679
; 
32'd160449: dataIn1 = 32'd9701
; 
32'd160450: dataIn1 = 32'd9702
; 
32'd160451: dataIn1 = 32'd9793
; 
32'd160452: dataIn1 = 32'd9794
; 
32'd160453: dataIn1 = 32'd6088
; 
32'd160454: dataIn1 = 32'd9677
; 
32'd160455: dataIn1 = 32'd9678
; 
32'd160456: dataIn1 = 32'd9721
; 
32'd160457: dataIn1 = 32'd9722
; 
32'd160458: dataIn1 = 32'd9791
; 
32'd160459: dataIn1 = 32'd9792
; 
32'd160460: dataIn1 = 32'd6089
; 
32'd160461: dataIn1 = 32'd7099
; 
32'd160462: dataIn1 = 32'd7101
; 
32'd160463: dataIn1 = 32'd7102
; 
32'd160464: dataIn1 = 32'd7103
; 
32'd160465: dataIn1 = 32'd7203
; 
32'd160466: dataIn1 = 32'd7205
; 
32'd160467: dataIn1 = 32'd6090
; 
32'd160468: dataIn1 = 32'd6091
; 
32'd160469: dataIn1 = 32'd6092
; 
32'd160470: dataIn1 = 32'd7105
; 
32'd160471: dataIn1 = 32'd7106
; 
32'd160472: dataIn1 = 32'd7109
; 
32'd160473: dataIn1 = 32'd7110
; 
32'd160474: dataIn1 = 32'd5114
; 
32'd160475: dataIn1 = 32'd5119
; 
32'd160476: dataIn1 = 32'd6072
; 
32'd160477: dataIn1 = 32'd6090
; 
32'd160478: dataIn1 = 32'd6091
; 
32'd160479: dataIn1 = 32'd6092
; 
32'd160480: dataIn1 = 32'd6094
; 
32'd160481: dataIn1 = 32'd7110
; 
32'd160482: dataIn1 = 32'd5119
; 
32'd160483: dataIn1 = 32'd5120
; 
32'd160484: dataIn1 = 32'd6090
; 
32'd160485: dataIn1 = 32'd6091
; 
32'd160486: dataIn1 = 32'd6092
; 
32'd160487: dataIn1 = 32'd6095
; 
32'd160488: dataIn1 = 32'd6096
; 
32'd160489: dataIn1 = 32'd7109
; 
32'd160490: dataIn1 = 32'd6093
; 
32'd160491: dataIn1 = 32'd7104
; 
32'd160492: dataIn1 = 32'd7105
; 
32'd160493: dataIn1 = 32'd7107
; 
32'd160494: dataIn1 = 32'd7108
; 
32'd160495: dataIn1 = 32'd7155
; 
32'd160496: dataIn1 = 32'd7156
; 
32'd160497: dataIn1 = 32'd2693
; 
32'd160498: dataIn1 = 32'd5119
; 
32'd160499: dataIn1 = 32'd6072
; 
32'd160500: dataIn1 = 32'd6091
; 
32'd160501: dataIn1 = 32'd6094
; 
32'd160502: dataIn1 = 32'd6707
; 
32'd160503: dataIn1 = 32'd1120
; 
32'd160504: dataIn1 = 32'd5120
; 
32'd160505: dataIn1 = 32'd6092
; 
32'd160506: dataIn1 = 32'd6095
; 
32'd160507: dataIn1 = 32'd6096
; 
32'd160508: dataIn1 = 32'd6116
; 
32'd160509: dataIn1 = 32'd6118
; 
32'd160510: dataIn1 = 32'd7151
; 
32'd160511: dataIn1 = 32'd1120
; 
32'd160512: dataIn1 = 32'd5119
; 
32'd160513: dataIn1 = 32'd6092
; 
32'd160514: dataIn1 = 32'd6095
; 
32'd160515: dataIn1 = 32'd6096
; 
32'd160516: dataIn1 = 32'd6706
; 
32'd160517: dataIn1 = 32'd6097
; 
32'd160518: dataIn1 = 32'd7112
; 
32'd160519: dataIn1 = 32'd7113
; 
32'd160520: dataIn1 = 32'd7117
; 
32'd160521: dataIn1 = 32'd7119
; 
32'd160522: dataIn1 = 32'd7121
; 
32'd160523: dataIn1 = 32'd7122
; 
32'd160524: dataIn1 = 32'd6098
; 
32'd160525: dataIn1 = 32'd7111
; 
32'd160526: dataIn1 = 32'd7113
; 
32'd160527: dataIn1 = 32'd7115
; 
32'd160528: dataIn1 = 32'd7118
; 
32'd160529: dataIn1 = 32'd7127
; 
32'd160530: dataIn1 = 32'd7129
; 
32'd160531: dataIn1 = 32'd6099
; 
32'd160532: dataIn1 = 32'd7111
; 
32'd160533: dataIn1 = 32'd7112
; 
32'd160534: dataIn1 = 32'd7114
; 
32'd160535: dataIn1 = 32'd7116
; 
32'd160536: dataIn1 = 32'd9800
; 
32'd160537: dataIn1 = 32'd9801
; 
32'd160538: dataIn1 = 32'd6100
; 
32'd160539: dataIn1 = 32'd7120
; 
32'd160540: dataIn1 = 32'd7122
; 
32'd160541: dataIn1 = 32'd7124
; 
32'd160542: dataIn1 = 32'd7126
; 
32'd160543: dataIn1 = 32'd7155
; 
32'd160544: dataIn1 = 32'd7157
; 
32'd160545: dataIn1 = 32'd6101
; 
32'd160546: dataIn1 = 32'd7120
; 
32'd160547: dataIn1 = 32'd7121
; 
32'd160548: dataIn1 = 32'd7123
; 
32'd160549: dataIn1 = 32'd7125
; 
32'd160550: dataIn1 = 32'd7141
; 
32'd160551: dataIn1 = 32'd7142
; 
32'd160552: dataIn1 = 32'd6102
; 
32'd160553: dataIn1 = 32'd7128
; 
32'd160554: dataIn1 = 32'd7129
; 
32'd160555: dataIn1 = 32'd7132
; 
32'd160556: dataIn1 = 32'd7133
; 
32'd160557: dataIn1 = 32'd7159
; 
32'd160558: dataIn1 = 32'd7160
; 
32'd160559: dataIn1 = 32'd6103
; 
32'd160560: dataIn1 = 32'd7127
; 
32'd160561: dataIn1 = 32'd7128
; 
32'd160562: dataIn1 = 32'd7130
; 
32'd160563: dataIn1 = 32'd7131
; 
32'd160564: dataIn1 = 32'd7134
; 
32'd160565: dataIn1 = 32'd7135
; 
32'd160566: dataIn1 = 32'd6104
; 
32'd160567: dataIn1 = 32'd9681
; 
32'd160568: dataIn1 = 32'd9682
; 
32'd160569: dataIn1 = 32'd9706
; 
32'd160570: dataIn1 = 32'd9707
; 
32'd160571: dataIn1 = 32'd9799
; 
32'd160572: dataIn1 = 32'd9800
; 
32'd160573: dataIn1 = 32'd6105
; 
32'd160574: dataIn1 = 32'd9680
; 
32'd160575: dataIn1 = 32'd9682
; 
32'd160576: dataIn1 = 32'd9692
; 
32'd160577: dataIn1 = 32'd9694
; 
32'd160578: dataIn1 = 32'd9801
; 
32'd160579: dataIn1 = 32'd9802
; 
32'd160580: dataIn1 = 32'd6106
; 
32'd160581: dataIn1 = 32'd9684
; 
32'd160582: dataIn1 = 32'd9685
; 
32'd160583: dataIn1 = 32'd9687
; 
32'd160584: dataIn1 = 32'd9688
; 
32'd160585: dataIn1 = 32'd9805
; 
32'd160586: dataIn1 = 32'd9806
; 
32'd160587: dataIn1 = 32'd6107
; 
32'd160588: dataIn1 = 32'd7134
; 
32'd160589: dataIn1 = 32'd7136
; 
32'd160590: dataIn1 = 32'd7137
; 
32'd160591: dataIn1 = 32'd7139
; 
32'd160592: dataIn1 = 32'd9804
; 
32'd160593: dataIn1 = 32'd9805
; 
32'd160594: dataIn1 = 32'd6108
; 
32'd160595: dataIn1 = 32'd9683
; 
32'd160596: dataIn1 = 32'd9684
; 
32'd160597: dataIn1 = 32'd9692
; 
32'd160598: dataIn1 = 32'd9693
; 
32'd160599: dataIn1 = 32'd9803
; 
32'd160600: dataIn1 = 32'd9804
; 
32'd160601: dataIn1 = 32'd6109
; 
32'd160602: dataIn1 = 32'd9686
; 
32'd160603: dataIn1 = 32'd9688
; 
32'd160604: dataIn1 = 32'd9690
; 
32'd160605: dataIn1 = 32'd9756
; 
32'd160606: dataIn1 = 32'd9807
; 
32'd160607: dataIn1 = 32'd9808
; 
32'd160608: dataIn1 = 32'd6110
; 
32'd160609: dataIn1 = 32'd7135
; 
32'd160610: dataIn1 = 32'd7136
; 
32'd160611: dataIn1 = 32'd7138
; 
32'd160612: dataIn1 = 32'd7140
; 
32'd160613: dataIn1 = 32'd9378
; 
32'd160614: dataIn1 = 32'd9379
; 
32'd160615: dataIn1 = 32'd6111
; 
32'd160616: dataIn1 = 32'd7142
; 
32'd160617: dataIn1 = 32'd7143
; 
32'd160618: dataIn1 = 32'd7144
; 
32'd160619: dataIn1 = 32'd7145
; 
32'd160620: dataIn1 = 32'd9796
; 
32'd160621: dataIn1 = 32'd9797
; 
32'd160622: dataIn1 = 32'd6112
; 
32'd160623: dataIn1 = 32'd9697
; 
32'd160624: dataIn1 = 32'd9699
; 
32'd160625: dataIn1 = 32'd9700
; 
32'd160626: dataIn1 = 32'd9702
; 
32'd160627: dataIn1 = 32'd9795
; 
32'd160628: dataIn1 = 32'd9796
; 
32'd160629: dataIn1 = 32'd6113
; 
32'd160630: dataIn1 = 32'd9697
; 
32'd160631: dataIn1 = 32'd9698
; 
32'd160632: dataIn1 = 32'd9705
; 
32'd160633: dataIn1 = 32'd9706
; 
32'd160634: dataIn1 = 32'd9797
; 
32'd160635: dataIn1 = 32'd9798
; 
32'd160636: dataIn1 = 32'd6114
; 
32'd160637: dataIn1 = 32'd7147
; 
32'd160638: dataIn1 = 32'd7148
; 
32'd160639: dataIn1 = 32'd7152
; 
32'd160640: dataIn1 = 32'd7154
; 
32'd160641: dataIn1 = 32'd7156
; 
32'd160642: dataIn1 = 32'd7157
; 
32'd160643: dataIn1 = 32'd6115
; 
32'd160644: dataIn1 = 32'd7146
; 
32'd160645: dataIn1 = 32'd7148
; 
32'd160646: dataIn1 = 32'd7150
; 
32'd160647: dataIn1 = 32'd7153
; 
32'd160648: dataIn1 = 32'd7158
; 
32'd160649: dataIn1 = 32'd7160
; 
32'd160650: dataIn1 = 32'd6095
; 
32'd160651: dataIn1 = 32'd6116
; 
32'd160652: dataIn1 = 32'd6118
; 
32'd160653: dataIn1 = 32'd7146
; 
32'd160654: dataIn1 = 32'd7147
; 
32'd160655: dataIn1 = 32'd7149
; 
32'd160656: dataIn1 = 32'd7151
; 
32'd160657: dataIn1 = 32'd6117
; 
32'd160658: dataIn1 = 32'd7158
; 
32'd160659: dataIn1 = 32'd7159
; 
32'd160660: dataIn1 = 32'd7161
; 
32'd160661: dataIn1 = 32'd7162
; 
32'd160662: dataIn1 = 32'd9380
; 
32'd160663: dataIn1 = 32'd9382
; 
32'd160664: dataIn1 = 32'd1120
; 
32'd160665: dataIn1 = 32'd5125
; 
32'd160666: dataIn1 = 32'd6095
; 
32'd160667: dataIn1 = 32'd6116
; 
32'd160668: dataIn1 = 32'd6118
; 
32'd160669: dataIn1 = 32'd6817
; 
32'd160670: dataIn1 = 32'd6820
; 
32'd160671: dataIn1 = 32'd7149
; 
32'd160672: dataIn1 = 32'd6119
; 
32'd160673: dataIn1 = 32'd7164
; 
32'd160674: dataIn1 = 32'd7165
; 
32'd160675: dataIn1 = 32'd7169
; 
32'd160676: dataIn1 = 32'd7171
; 
32'd160677: dataIn1 = 32'd9777
; 
32'd160678: dataIn1 = 32'd9785
; 
32'd160679: dataIn1 = 32'd6120
; 
32'd160680: dataIn1 = 32'd7163
; 
32'd160681: dataIn1 = 32'd7165
; 
32'd160682: dataIn1 = 32'd7167
; 
32'd160683: dataIn1 = 32'd7170
; 
32'd160684: dataIn1 = 32'd7172
; 
32'd160685: dataIn1 = 32'd7174
; 
32'd160686: dataIn1 = 32'd6121
; 
32'd160687: dataIn1 = 32'd7163
; 
32'd160688: dataIn1 = 32'd7164
; 
32'd160689: dataIn1 = 32'd7166
; 
32'd160690: dataIn1 = 32'd7168
; 
32'd160691: dataIn1 = 32'd7179
; 
32'd160692: dataIn1 = 32'd7180
; 
32'd160693: dataIn1 = 32'd6122
; 
32'd160694: dataIn1 = 32'd9710
; 
32'd160695: dataIn1 = 32'd9712
; 
32'd160696: dataIn1 = 32'd9726
; 
32'd160697: dataIn1 = 32'd9728
; 
32'd160698: dataIn1 = 32'd9759
; 
32'd160699: dataIn1 = 32'd9777
; 
32'd160700: dataIn1 = 32'd6123
; 
32'd160701: dataIn1 = 32'd9710
; 
32'd160702: dataIn1 = 32'd9711
; 
32'd160703: dataIn1 = 32'd9716
; 
32'd160704: dataIn1 = 32'd9717
; 
32'd160705: dataIn1 = 32'd9785
; 
32'd160706: dataIn1 = 32'd9786
; 
32'd160707: dataIn1 = 32'd6124
; 
32'd160708: dataIn1 = 32'd7173
; 
32'd160709: dataIn1 = 32'd7174
; 
32'd160710: dataIn1 = 32'd7177
; 
32'd160711: dataIn1 = 32'd7178
; 
32'd160712: dataIn1 = 32'd7216
; 
32'd160713: dataIn1 = 32'd7217
; 
32'd160714: dataIn1 = 32'd6125
; 
32'd160715: dataIn1 = 32'd7172
; 
32'd160716: dataIn1 = 32'd7173
; 
32'd160717: dataIn1 = 32'd7175
; 
32'd160718: dataIn1 = 32'd7176
; 
32'd160719: dataIn1 = 32'd7195
; 
32'd160720: dataIn1 = 32'd7196
; 
32'd160721: dataIn1 = 32'd6126
; 
32'd160722: dataIn1 = 32'd7180
; 
32'd160723: dataIn1 = 32'd7181
; 
32'd160724: dataIn1 = 32'd7183
; 
32'd160725: dataIn1 = 32'd7185
; 
32'd160726: dataIn1 = 32'd7204
; 
32'd160727: dataIn1 = 32'd7205
; 
32'd160728: dataIn1 = 32'd6127
; 
32'd160729: dataIn1 = 32'd7179
; 
32'd160730: dataIn1 = 32'd7181
; 
32'd160731: dataIn1 = 32'd7182
; 
32'd160732: dataIn1 = 32'd7184
; 
32'd160733: dataIn1 = 32'd7200
; 
32'd160734: dataIn1 = 32'd7202
; 
32'd160735: dataIn1 = 32'd6080
; 
32'd160736: dataIn1 = 32'd6128
; 
32'd160737: dataIn1 = 32'd6131
; 
32'd160738: dataIn1 = 32'd7187
; 
32'd160739: dataIn1 = 32'd7188
; 
32'd160740: dataIn1 = 32'd7192
; 
32'd160741: dataIn1 = 32'd7194
; 
32'd160742: dataIn1 = 32'd6129
; 
32'd160743: dataIn1 = 32'd7186
; 
32'd160744: dataIn1 = 32'd7188
; 
32'd160745: dataIn1 = 32'd7190
; 
32'd160746: dataIn1 = 32'd7193
; 
32'd160747: dataIn1 = 32'd7195
; 
32'd160748: dataIn1 = 32'd7197
; 
32'd160749: dataIn1 = 32'd6130
; 
32'd160750: dataIn1 = 32'd7186
; 
32'd160751: dataIn1 = 32'd7187
; 
32'd160752: dataIn1 = 32'd7189
; 
32'd160753: dataIn1 = 32'd7191
; 
32'd160754: dataIn1 = 32'd7200
; 
32'd160755: dataIn1 = 32'd7201
; 
32'd160756: dataIn1 = 32'd1119
; 
32'd160757: dataIn1 = 32'd5129
; 
32'd160758: dataIn1 = 32'd6080
; 
32'd160759: dataIn1 = 32'd6128
; 
32'd160760: dataIn1 = 32'd6131
; 
32'd160761: dataIn1 = 32'd6592
; 
32'd160762: dataIn1 = 32'd6594
; 
32'd160763: dataIn1 = 32'd7194
; 
32'd160764: dataIn1 = 32'd6132
; 
32'd160765: dataIn1 = 32'd7196
; 
32'd160766: dataIn1 = 32'd7197
; 
32'd160767: dataIn1 = 32'd7198
; 
32'd160768: dataIn1 = 32'd7199
; 
32'd160769: dataIn1 = 32'd8916
; 
32'd160770: dataIn1 = 32'd8917
; 
32'd160771: dataIn1 = 32'd6133
; 
32'd160772: dataIn1 = 32'd9714
; 
32'd160773: dataIn1 = 32'd9715
; 
32'd160774: dataIn1 = 32'd9717
; 
32'd160775: dataIn1 = 32'd9718
; 
32'd160776: dataIn1 = 32'd9787
; 
32'd160777: dataIn1 = 32'd9788
; 
32'd160778: dataIn1 = 32'd6134
; 
32'd160779: dataIn1 = 32'd9713
; 
32'd160780: dataIn1 = 32'd9715
; 
32'd160781: dataIn1 = 32'd9721
; 
32'd160782: dataIn1 = 32'd9723
; 
32'd160783: dataIn1 = 32'd9789
; 
32'd160784: dataIn1 = 32'd9790
; 
32'd160785: dataIn1 = 32'd6135
; 
32'd160786: dataIn1 = 32'd7203
; 
32'd160787: dataIn1 = 32'd7204
; 
32'd160788: dataIn1 = 32'd7206
; 
32'd160789: dataIn1 = 32'd7207
; 
32'd160790: dataIn1 = 32'd9788
; 
32'd160791: dataIn1 = 32'd9789
; 
32'd160792: dataIn1 = 32'd6136
; 
32'd160793: dataIn1 = 32'd7209
; 
32'd160794: dataIn1 = 32'd7210
; 
32'd160795: dataIn1 = 32'd7214
; 
32'd160796: dataIn1 = 32'd9727
; 
32'd160797: dataIn1 = 32'd9728
; 
32'd160798: dataIn1 = 32'd9731
; 
32'd160799: dataIn1 = 32'd6137
; 
32'd160800: dataIn1 = 32'd7208
; 
32'd160801: dataIn1 = 32'd7210
; 
32'd160802: dataIn1 = 32'd7212
; 
32'd160803: dataIn1 = 32'd7213
; 
32'd160804: dataIn1 = 32'd7215
; 
32'd160805: dataIn1 = 32'd7217
; 
32'd160806: dataIn1 = 32'd4817
; 
32'd160807: dataIn1 = 32'd6138
; 
32'd160808: dataIn1 = 32'd7208
; 
32'd160809: dataIn1 = 32'd7209
; 
32'd160810: dataIn1 = 32'd7211
; 
32'd160811: dataIn1 = 32'd7220
; 
32'd160812: dataIn1 = 32'd9758
; 
32'd160813: dataIn1 = 32'd6139
; 
32'd160814: dataIn1 = 32'd7215
; 
32'd160815: dataIn1 = 32'd7216
; 
32'd160816: dataIn1 = 32'd7218
; 
32'd160817: dataIn1 = 32'd7219
; 
32'd160818: dataIn1 = 32'd8906
; 
32'd160819: dataIn1 = 32'd8907
; 
32'd160820: dataIn1 = 32'd4
; 
32'd160821: dataIn1 = 32'd4817
; 
32'd160822: dataIn1 = 32'd6140
; 
32'd160823: dataIn1 = 32'd7220
; 
32'd160824: dataIn1 = 32'd7221
; 
32'd160825: dataIn1 = 32'd8902
; 
32'd160826: dataIn1 = 32'd8904
; 
32'd160827: dataIn1 = 32'd6141
; 
32'd160828: dataIn1 = 32'd6142
; 
32'd160829: dataIn1 = 32'd6143
; 
32'd160830: dataIn1 = 32'd7241
; 
32'd160831: dataIn1 = 32'd7242
; 
32'd160832: dataIn1 = 32'd7244
; 
32'd160833: dataIn1 = 32'd7246
; 
32'd160834: dataIn1 = 32'd2699
; 
32'd160835: dataIn1 = 32'd5131
; 
32'd160836: dataIn1 = 32'd6141
; 
32'd160837: dataIn1 = 32'd6142
; 
32'd160838: dataIn1 = 32'd6143
; 
32'd160839: dataIn1 = 32'd6144
; 
32'd160840: dataIn1 = 32'd6145
; 
32'd160841: dataIn1 = 32'd7246
; 
32'd160842: dataIn1 = 32'd5131
; 
32'd160843: dataIn1 = 32'd5132
; 
32'd160844: dataIn1 = 32'd5133
; 
32'd160845: dataIn1 = 32'd6141
; 
32'd160846: dataIn1 = 32'd6142
; 
32'd160847: dataIn1 = 32'd6143
; 
32'd160848: dataIn1 = 32'd7244
; 
32'd160849: dataIn1 = 32'd2699
; 
32'd160850: dataIn1 = 32'd5134
; 
32'd160851: dataIn1 = 32'd6142
; 
32'd160852: dataIn1 = 32'd6144
; 
32'd160853: dataIn1 = 32'd6145
; 
32'd160854: dataIn1 = 32'd6176
; 
32'd160855: dataIn1 = 32'd6179
; 
32'd160856: dataIn1 = 32'd7310
; 
32'd160857: dataIn1 = 32'd5131
; 
32'd160858: dataIn1 = 32'd5134
; 
32'd160859: dataIn1 = 32'd5135
; 
32'd160860: dataIn1 = 32'd6142
; 
32'd160861: dataIn1 = 32'd6144
; 
32'd160862: dataIn1 = 32'd6145
; 
32'd160863: dataIn1 = 32'd6146
; 
32'd160864: dataIn1 = 32'd6150
; 
32'd160865: dataIn1 = 32'd7223
; 
32'd160866: dataIn1 = 32'd7224
; 
32'd160867: dataIn1 = 32'd7228
; 
32'd160868: dataIn1 = 32'd7230
; 
32'd160869: dataIn1 = 32'd7232
; 
32'd160870: dataIn1 = 32'd6147
; 
32'd160871: dataIn1 = 32'd7222
; 
32'd160872: dataIn1 = 32'd7224
; 
32'd160873: dataIn1 = 32'd7226
; 
32'd160874: dataIn1 = 32'd7229
; 
32'd160875: dataIn1 = 32'd7233
; 
32'd160876: dataIn1 = 32'd7235
; 
32'd160877: dataIn1 = 32'd6148
; 
32'd160878: dataIn1 = 32'd7222
; 
32'd160879: dataIn1 = 32'd7223
; 
32'd160880: dataIn1 = 32'd7225
; 
32'd160881: dataIn1 = 32'd7227
; 
32'd160882: dataIn1 = 32'd7240
; 
32'd160883: dataIn1 = 32'd7241
; 
32'd160884: dataIn1 = 32'd2697
; 
32'd160885: dataIn1 = 32'd6149
; 
32'd160886: dataIn1 = 32'd6150
; 
32'd160887: dataIn1 = 32'd7231
; 
32'd160888: dataIn1 = 32'd7232
; 
32'd160889: dataIn1 = 32'd7272
; 
32'd160890: dataIn1 = 32'd7274
; 
32'd160891: dataIn1 = 32'd2697
; 
32'd160892: dataIn1 = 32'd5132
; 
32'd160893: dataIn1 = 32'd5133
; 
32'd160894: dataIn1 = 32'd6146
; 
32'd160895: dataIn1 = 32'd6149
; 
32'd160896: dataIn1 = 32'd6150
; 
32'd160897: dataIn1 = 32'd7228
; 
32'd160898: dataIn1 = 32'd7232
; 
32'd160899: dataIn1 = 32'd6151
; 
32'd160900: dataIn1 = 32'd7234
; 
32'd160901: dataIn1 = 32'd7235
; 
32'd160902: dataIn1 = 32'd7238
; 
32'd160903: dataIn1 = 32'd7239
; 
32'd160904: dataIn1 = 32'd7277
; 
32'd160905: dataIn1 = 32'd7278
; 
32'd160906: dataIn1 = 32'd6152
; 
32'd160907: dataIn1 = 32'd7233
; 
32'd160908: dataIn1 = 32'd7234
; 
32'd160909: dataIn1 = 32'd7236
; 
32'd160910: dataIn1 = 32'd7237
; 
32'd160911: dataIn1 = 32'd7329
; 
32'd160912: dataIn1 = 32'd7330
; 
32'd160913: dataIn1 = 32'd6153
; 
32'd160914: dataIn1 = 32'd7240
; 
32'd160915: dataIn1 = 32'd7242
; 
32'd160916: dataIn1 = 32'd7243
; 
32'd160917: dataIn1 = 32'd7245
; 
32'd160918: dataIn1 = 32'd7332
; 
32'd160919: dataIn1 = 32'd7334
; 
32'd160920: dataIn1 = 32'd5142
; 
32'd160921: dataIn1 = 32'd6154
; 
32'd160922: dataIn1 = 32'd6157
; 
32'd160923: dataIn1 = 32'd9733
; 
32'd160924: dataIn1 = 32'd9734
; 
32'd160925: dataIn1 = 32'd9761
; 
32'd160926: dataIn1 = 32'd9762
; 
32'd160927: dataIn1 = 32'd5142
; 
32'd160928: dataIn1 = 32'd6155
; 
32'd160929: dataIn1 = 32'd9668
; 
32'd160930: dataIn1 = 32'd9732
; 
32'd160931: dataIn1 = 32'd9734
; 
32'd160932: dataIn1 = 32'd9760
; 
32'd160933: dataIn1 = 32'd10150
; 
32'd160934: dataIn1 = 32'd6156
; 
32'd160935: dataIn1 = 32'd7247
; 
32'd160936: dataIn1 = 32'd7248
; 
32'd160937: dataIn1 = 32'd7250
; 
32'd160938: dataIn1 = 32'd7252
; 
32'd160939: dataIn1 = 32'd9732
; 
32'd160940: dataIn1 = 32'd9733
; 
32'd160941: dataIn1 = 32'd2697
; 
32'd160942: dataIn1 = 32'd5139
; 
32'd160943: dataIn1 = 32'd5142
; 
32'd160944: dataIn1 = 32'd6154
; 
32'd160945: dataIn1 = 32'd6157
; 
32'd160946: dataIn1 = 32'd6158
; 
32'd160947: dataIn1 = 32'd9762
; 
32'd160948: dataIn1 = 32'd2697
; 
32'd160949: dataIn1 = 32'd6157
; 
32'd160950: dataIn1 = 32'd6158
; 
32'd160951: dataIn1 = 32'd7272
; 
32'd160952: dataIn1 = 32'd7273
; 
32'd160953: dataIn1 = 32'd7275
; 
32'd160954: dataIn1 = 32'd9762
; 
32'd160955: dataIn1 = 32'd6159
; 
32'd160956: dataIn1 = 32'd7248
; 
32'd160957: dataIn1 = 32'd7249
; 
32'd160958: dataIn1 = 32'd7253
; 
32'd160959: dataIn1 = 32'd7255
; 
32'd160960: dataIn1 = 32'd7280
; 
32'd160961: dataIn1 = 32'd7281
; 
32'd160962: dataIn1 = 32'd6160
; 
32'd160963: dataIn1 = 32'd7247
; 
32'd160964: dataIn1 = 32'd7249
; 
32'd160965: dataIn1 = 32'd7251
; 
32'd160966: dataIn1 = 32'd7254
; 
32'd160967: dataIn1 = 32'd7259
; 
32'd160968: dataIn1 = 32'd7261
; 
32'd160969: dataIn1 = 32'd6161
; 
32'd160970: dataIn1 = 32'd7257
; 
32'd160971: dataIn1 = 32'd7258
; 
32'd160972: dataIn1 = 32'd9232
; 
32'd160973: dataIn1 = 32'd9286
; 
32'd160974: dataIn1 = 32'd9778
; 
32'd160975: dataIn1 = 32'd10151
; 
32'd160976: dataIn1 = 32'd6162
; 
32'd160977: dataIn1 = 32'd10119
; 
32'd160978: dataIn1 = 32'd10121
; 
32'd160979: dataIn1 = 32'd10123
; 
32'd160980: dataIn1 = 32'd10124
; 
32'd160981: dataIn1 = 32'd10151
; 
32'd160982: dataIn1 = 32'd10220
; 
32'd160983: dataIn1 = 32'd6163
; 
32'd160984: dataIn1 = 32'd7259
; 
32'd160985: dataIn1 = 32'd7260
; 
32'd160986: dataIn1 = 32'd7262
; 
32'd160987: dataIn1 = 32'd9274
; 
32'd160988: dataIn1 = 32'd9286
; 
32'd160989: dataIn1 = 32'd10220
; 
32'd160990: dataIn1 = 32'd6164
; 
32'd160991: dataIn1 = 32'd7256
; 
32'd160992: dataIn1 = 32'd7258
; 
32'd160993: dataIn1 = 32'd8921
; 
32'd160994: dataIn1 = 32'd8922
; 
32'd160995: dataIn1 = 32'd8924
; 
32'd160996: dataIn1 = 32'd9767
; 
32'd160997: dataIn1 = 32'd6165
; 
32'd160998: dataIn1 = 32'd7264
; 
32'd160999: dataIn1 = 32'd7265
; 
32'd161000: dataIn1 = 32'd7269
; 
32'd161001: dataIn1 = 32'd7271
; 
32'd161002: dataIn1 = 32'd7273
; 
32'd161003: dataIn1 = 32'd7274
; 
32'd161004: dataIn1 = 32'd6166
; 
32'd161005: dataIn1 = 32'd7263
; 
32'd161006: dataIn1 = 32'd7265
; 
32'd161007: dataIn1 = 32'd7267
; 
32'd161008: dataIn1 = 32'd7270
; 
32'd161009: dataIn1 = 32'd7276
; 
32'd161010: dataIn1 = 32'd7278
; 
32'd161011: dataIn1 = 32'd6167
; 
32'd161012: dataIn1 = 32'd7263
; 
32'd161013: dataIn1 = 32'd7264
; 
32'd161014: dataIn1 = 32'd7266
; 
32'd161015: dataIn1 = 32'd7268
; 
32'd161016: dataIn1 = 32'd7279
; 
32'd161017: dataIn1 = 32'd7280
; 
32'd161018: dataIn1 = 32'd6168
; 
32'd161019: dataIn1 = 32'd7283
; 
32'd161020: dataIn1 = 32'd7284
; 
32'd161021: dataIn1 = 32'd7288
; 
32'd161022: dataIn1 = 32'd7290
; 
32'd161023: dataIn1 = 32'd7292
; 
32'd161024: dataIn1 = 32'd7293
; 
32'd161025: dataIn1 = 32'd6169
; 
32'd161026: dataIn1 = 32'd7282
; 
32'd161027: dataIn1 = 32'd7284
; 
32'd161028: dataIn1 = 32'd7286
; 
32'd161029: dataIn1 = 32'd7289
; 
32'd161030: dataIn1 = 32'd7298
; 
32'd161031: dataIn1 = 32'd7300
; 
32'd161032: dataIn1 = 32'd6170
; 
32'd161033: dataIn1 = 32'd7282
; 
32'd161034: dataIn1 = 32'd7283
; 
32'd161035: dataIn1 = 32'd7285
; 
32'd161036: dataIn1 = 32'd7287
; 
32'd161037: dataIn1 = 32'd7305
; 
32'd161038: dataIn1 = 32'd7306
; 
32'd161039: dataIn1 = 32'd6171
; 
32'd161040: dataIn1 = 32'd7291
; 
32'd161041: dataIn1 = 32'd7293
; 
32'd161042: dataIn1 = 32'd7295
; 
32'd161043: dataIn1 = 32'd7297
; 
32'd161044: dataIn1 = 32'd7344
; 
32'd161045: dataIn1 = 32'd7346
; 
32'd161046: dataIn1 = 32'd6172
; 
32'd161047: dataIn1 = 32'd7291
; 
32'd161048: dataIn1 = 32'd7292
; 
32'd161049: dataIn1 = 32'd7294
; 
32'd161050: dataIn1 = 32'd7296
; 
32'd161051: dataIn1 = 32'd7326
; 
32'd161052: dataIn1 = 32'd7327
; 
32'd161053: dataIn1 = 32'd6173
; 
32'd161054: dataIn1 = 32'd7299
; 
32'd161055: dataIn1 = 32'd7300
; 
32'd161056: dataIn1 = 32'd7303
; 
32'd161057: dataIn1 = 32'd7304
; 
32'd161058: dataIn1 = 32'd7348
; 
32'd161059: dataIn1 = 32'd7349
; 
32'd161060: dataIn1 = 32'd6174
; 
32'd161061: dataIn1 = 32'd7298
; 
32'd161062: dataIn1 = 32'd7299
; 
32'd161063: dataIn1 = 32'd7301
; 
32'd161064: dataIn1 = 32'd7302
; 
32'd161065: dataIn1 = 32'd7312
; 
32'd161066: dataIn1 = 32'd7313
; 
32'd161067: dataIn1 = 32'd6175
; 
32'd161068: dataIn1 = 32'd7306
; 
32'd161069: dataIn1 = 32'd7307
; 
32'd161070: dataIn1 = 32'd7309
; 
32'd161071: dataIn1 = 32'd7311
; 
32'd161072: dataIn1 = 32'd7333
; 
32'd161073: dataIn1 = 32'd7334
; 
32'd161074: dataIn1 = 32'd6144
; 
32'd161075: dataIn1 = 32'd6176
; 
32'd161076: dataIn1 = 32'd6179
; 
32'd161077: dataIn1 = 32'd7305
; 
32'd161078: dataIn1 = 32'd7307
; 
32'd161079: dataIn1 = 32'd7308
; 
32'd161080: dataIn1 = 32'd7310
; 
32'd161081: dataIn1 = 32'd1121
; 
32'd161082: dataIn1 = 32'd5134
; 
32'd161083: dataIn1 = 32'd5148
; 
32'd161084: dataIn1 = 32'd6177
; 
32'd161085: dataIn1 = 32'd6178
; 
32'd161086: dataIn1 = 32'd6179
; 
32'd161087: dataIn1 = 32'd5148
; 
32'd161088: dataIn1 = 32'd6177
; 
32'd161089: dataIn1 = 32'd6178
; 
32'd161090: dataIn1 = 32'd6179
; 
32'd161091: dataIn1 = 32'd7312
; 
32'd161092: dataIn1 = 32'd7314
; 
32'd161093: dataIn1 = 32'd7315
; 
32'd161094: dataIn1 = 32'd5134
; 
32'd161095: dataIn1 = 32'd5145
; 
32'd161096: dataIn1 = 32'd6144
; 
32'd161097: dataIn1 = 32'd6176
; 
32'd161098: dataIn1 = 32'd6177
; 
32'd161099: dataIn1 = 32'd6178
; 
32'd161100: dataIn1 = 32'd6179
; 
32'd161101: dataIn1 = 32'd7308
; 
32'd161102: dataIn1 = 32'd7315
; 
32'd161103: dataIn1 = 32'd5148
; 
32'd161104: dataIn1 = 32'd6180
; 
32'd161105: dataIn1 = 32'd6610
; 
32'd161106: dataIn1 = 32'd7313
; 
32'd161107: dataIn1 = 32'd7314
; 
32'd161108: dataIn1 = 32'd7316
; 
32'd161109: dataIn1 = 32'd8975
; 
32'd161110: dataIn1 = 32'd6181
; 
32'd161111: dataIn1 = 32'd7318
; 
32'd161112: dataIn1 = 32'd7319
; 
32'd161113: dataIn1 = 32'd7323
; 
32'd161114: dataIn1 = 32'd7325
; 
32'd161115: dataIn1 = 32'd7327
; 
32'd161116: dataIn1 = 32'd7328
; 
32'd161117: dataIn1 = 32'd6182
; 
32'd161118: dataIn1 = 32'd7317
; 
32'd161119: dataIn1 = 32'd7319
; 
32'd161120: dataIn1 = 32'd7321
; 
32'd161121: dataIn1 = 32'd7324
; 
32'd161122: dataIn1 = 32'd7329
; 
32'd161123: dataIn1 = 32'd7331
; 
32'd161124: dataIn1 = 32'd6183
; 
32'd161125: dataIn1 = 32'd7317
; 
32'd161126: dataIn1 = 32'd7318
; 
32'd161127: dataIn1 = 32'd7320
; 
32'd161128: dataIn1 = 32'd7322
; 
32'd161129: dataIn1 = 32'd7332
; 
32'd161130: dataIn1 = 32'd7333
; 
32'd161131: dataIn1 = 32'd6184
; 
32'd161132: dataIn1 = 32'd7336
; 
32'd161133: dataIn1 = 32'd7337
; 
32'd161134: dataIn1 = 32'd7341
; 
32'd161135: dataIn1 = 32'd7343
; 
32'd161136: dataIn1 = 32'd7345
; 
32'd161137: dataIn1 = 32'd7346
; 
32'd161138: dataIn1 = 32'd6185
; 
32'd161139: dataIn1 = 32'd7335
; 
32'd161140: dataIn1 = 32'd7337
; 
32'd161141: dataIn1 = 32'd7339
; 
32'd161142: dataIn1 = 32'd7342
; 
32'd161143: dataIn1 = 32'd7347
; 
32'd161144: dataIn1 = 32'd7349
; 
32'd161145: dataIn1 = 32'd6186
; 
32'd161146: dataIn1 = 32'd7335
; 
32'd161147: dataIn1 = 32'd7336
; 
32'd161148: dataIn1 = 32'd7338
; 
32'd161149: dataIn1 = 32'd7340
; 
32'd161150: dataIn1 = 32'd7352
; 
32'd161151: dataIn1 = 32'd7353
; 
32'd161152: dataIn1 = 32'd6187
; 
32'd161153: dataIn1 = 32'd7347
; 
32'd161154: dataIn1 = 32'd7348
; 
32'd161155: dataIn1 = 32'd7350
; 
32'd161156: dataIn1 = 32'd7351
; 
32'd161157: dataIn1 = 32'd8965
; 
32'd161158: dataIn1 = 32'd8966
; 
32'd161159: dataIn1 = 32'd6188
; 
32'd161160: dataIn1 = 32'd7352
; 
32'd161161: dataIn1 = 32'd7354
; 
32'd161162: dataIn1 = 32'd7355
; 
32'd161163: dataIn1 = 32'd8959
; 
32'd161164: dataIn1 = 32'd8961
; 
32'd161165: dataIn1 = 32'd8963
; 
32'd161166: dataIn1 = 32'd6189
; 
32'd161167: dataIn1 = 32'd7357
; 
32'd161168: dataIn1 = 32'd7358
; 
32'd161169: dataIn1 = 32'd7362
; 
32'd161170: dataIn1 = 32'd7364
; 
32'd161171: dataIn1 = 32'd7366
; 
32'd161172: dataIn1 = 32'd7367
; 
32'd161173: dataIn1 = 32'd6190
; 
32'd161174: dataIn1 = 32'd6744
; 
32'd161175: dataIn1 = 32'd6745
; 
32'd161176: dataIn1 = 32'd7356
; 
32'd161177: dataIn1 = 32'd7358
; 
32'd161178: dataIn1 = 32'd7360
; 
32'd161179: dataIn1 = 32'd7363
; 
32'd161180: dataIn1 = 32'd6191
; 
32'd161181: dataIn1 = 32'd7356
; 
32'd161182: dataIn1 = 32'd7357
; 
32'd161183: dataIn1 = 32'd7359
; 
32'd161184: dataIn1 = 32'd7361
; 
32'd161185: dataIn1 = 32'd7372
; 
32'd161186: dataIn1 = 32'd7373
; 
32'd161187: dataIn1 = 32'd6192
; 
32'd161188: dataIn1 = 32'd7365
; 
32'd161189: dataIn1 = 32'd7367
; 
32'd161190: dataIn1 = 32'd7369
; 
32'd161191: dataIn1 = 32'd7371
; 
32'd161192: dataIn1 = 32'd7412
; 
32'd161193: dataIn1 = 32'd7414
; 
32'd161194: dataIn1 = 32'd6193
; 
32'd161195: dataIn1 = 32'd7365
; 
32'd161196: dataIn1 = 32'd7366
; 
32'd161197: dataIn1 = 32'd7368
; 
32'd161198: dataIn1 = 32'd7370
; 
32'd161199: dataIn1 = 32'd7395
; 
32'd161200: dataIn1 = 32'd7396
; 
32'd161201: dataIn1 = 32'd6194
; 
32'd161202: dataIn1 = 32'd7373
; 
32'd161203: dataIn1 = 32'd7374
; 
32'd161204: dataIn1 = 32'd7376
; 
32'd161205: dataIn1 = 32'd7378
; 
32'd161206: dataIn1 = 32'd7408
; 
32'd161207: dataIn1 = 32'd7409
; 
32'd161208: dataIn1 = 32'd6195
; 
32'd161209: dataIn1 = 32'd7372
; 
32'd161210: dataIn1 = 32'd7374
; 
32'd161211: dataIn1 = 32'd7375
; 
32'd161212: dataIn1 = 32'd7377
; 
32'd161213: dataIn1 = 32'd7379
; 
32'd161214: dataIn1 = 32'd7381
; 
32'd161215: dataIn1 = 32'd6196
; 
32'd161216: dataIn1 = 32'd7380
; 
32'd161217: dataIn1 = 32'd7381
; 
32'd161218: dataIn1 = 32'd7384
; 
32'd161219: dataIn1 = 32'd7385
; 
32'd161220: dataIn1 = 32'd7557
; 
32'd161221: dataIn1 = 32'd7558
; 
32'd161222: dataIn1 = 32'd6197
; 
32'd161223: dataIn1 = 32'd6746
; 
32'd161224: dataIn1 = 32'd6747
; 
32'd161225: dataIn1 = 32'd7379
; 
32'd161226: dataIn1 = 32'd7380
; 
32'd161227: dataIn1 = 32'd7382
; 
32'd161228: dataIn1 = 32'd7383
; 
32'd161229: dataIn1 = 32'd6198
; 
32'd161230: dataIn1 = 32'd7387
; 
32'd161231: dataIn1 = 32'd7388
; 
32'd161232: dataIn1 = 32'd7392
; 
32'd161233: dataIn1 = 32'd7394
; 
32'd161234: dataIn1 = 32'd7396
; 
32'd161235: dataIn1 = 32'd7397
; 
32'd161236: dataIn1 = 32'd6199
; 
32'd161237: dataIn1 = 32'd7386
; 
32'd161238: dataIn1 = 32'd7388
; 
32'd161239: dataIn1 = 32'd7390
; 
32'd161240: dataIn1 = 32'd7393
; 
32'd161241: dataIn1 = 32'd7400
; 
32'd161242: dataIn1 = 32'd7402
; 
32'd161243: dataIn1 = 32'd6200
; 
32'd161244: dataIn1 = 32'd7386
; 
32'd161245: dataIn1 = 32'd7387
; 
32'd161246: dataIn1 = 32'd7389
; 
32'd161247: dataIn1 = 32'd7391
; 
32'd161248: dataIn1 = 32'd7407
; 
32'd161249: dataIn1 = 32'd7408
; 
32'd161250: dataIn1 = 32'd6201
; 
32'd161251: dataIn1 = 32'd7395
; 
32'd161252: dataIn1 = 32'd7397
; 
32'd161253: dataIn1 = 32'd7398
; 
32'd161254: dataIn1 = 32'd7399
; 
32'd161255: dataIn1 = 32'd7482
; 
32'd161256: dataIn1 = 32'd7484
; 
32'd161257: dataIn1 = 32'd6202
; 
32'd161258: dataIn1 = 32'd7401
; 
32'd161259: dataIn1 = 32'd7402
; 
32'd161260: dataIn1 = 32'd7405
; 
32'd161261: dataIn1 = 32'd7406
; 
32'd161262: dataIn1 = 32'd7486
; 
32'd161263: dataIn1 = 32'd7487
; 
32'd161264: dataIn1 = 32'd6203
; 
32'd161265: dataIn1 = 32'd7400
; 
32'd161266: dataIn1 = 32'd7401
; 
32'd161267: dataIn1 = 32'd7403
; 
32'd161268: dataIn1 = 32'd7404
; 
32'd161269: dataIn1 = 32'd7573
; 
32'd161270: dataIn1 = 32'd7574
; 
32'd161271: dataIn1 = 32'd6204
; 
32'd161272: dataIn1 = 32'd7407
; 
32'd161273: dataIn1 = 32'd7409
; 
32'd161274: dataIn1 = 32'd7410
; 
32'd161275: dataIn1 = 32'd7411
; 
32'd161276: dataIn1 = 32'd7578
; 
32'd161277: dataIn1 = 32'd7580
; 
32'd161278: dataIn1 = 32'd6205
; 
32'd161279: dataIn1 = 32'd6748
; 
32'd161280: dataIn1 = 32'd6749
; 
32'd161281: dataIn1 = 32'd7413
; 
32'd161282: dataIn1 = 32'd7414
; 
32'd161283: dataIn1 = 32'd7417
; 
32'd161284: dataIn1 = 32'd7418
; 
32'd161285: dataIn1 = 32'd6206
; 
32'd161286: dataIn1 = 32'd7412
; 
32'd161287: dataIn1 = 32'd7413
; 
32'd161288: dataIn1 = 32'd7415
; 
32'd161289: dataIn1 = 32'd7416
; 
32'd161290: dataIn1 = 32'd7504
; 
32'd161291: dataIn1 = 32'd7505
; 
32'd161292: dataIn1 = 32'd6207
; 
32'd161293: dataIn1 = 32'd7420
; 
32'd161294: dataIn1 = 32'd7421
; 
32'd161295: dataIn1 = 32'd7425
; 
32'd161296: dataIn1 = 32'd7427
; 
32'd161297: dataIn1 = 32'd7429
; 
32'd161298: dataIn1 = 32'd7430
; 
32'd161299: dataIn1 = 32'd6208
; 
32'd161300: dataIn1 = 32'd7419
; 
32'd161301: dataIn1 = 32'd7421
; 
32'd161302: dataIn1 = 32'd7423
; 
32'd161303: dataIn1 = 32'd7426
; 
32'd161304: dataIn1 = 32'd7435
; 
32'd161305: dataIn1 = 32'd7437
; 
32'd161306: dataIn1 = 32'd6209
; 
32'd161307: dataIn1 = 32'd7419
; 
32'd161308: dataIn1 = 32'd7420
; 
32'd161309: dataIn1 = 32'd7422
; 
32'd161310: dataIn1 = 32'd7424
; 
32'd161311: dataIn1 = 32'd7442
; 
32'd161312: dataIn1 = 32'd7443
; 
32'd161313: dataIn1 = 32'd6210
; 
32'd161314: dataIn1 = 32'd7428
; 
32'd161315: dataIn1 = 32'd7430
; 
32'd161316: dataIn1 = 32'd7432
; 
32'd161317: dataIn1 = 32'd7434
; 
32'd161318: dataIn1 = 32'd7504
; 
32'd161319: dataIn1 = 32'd7506
; 
32'd161320: dataIn1 = 32'd6211
; 
32'd161321: dataIn1 = 32'd7428
; 
32'd161322: dataIn1 = 32'd7429
; 
32'd161323: dataIn1 = 32'd7431
; 
32'd161324: dataIn1 = 32'd7433
; 
32'd161325: dataIn1 = 32'd7482
; 
32'd161326: dataIn1 = 32'd7483
; 
32'd161327: dataIn1 = 32'd6212
; 
32'd161328: dataIn1 = 32'd7436
; 
32'd161329: dataIn1 = 32'd7437
; 
32'd161330: dataIn1 = 32'd7440
; 
32'd161331: dataIn1 = 32'd7441
; 
32'd161332: dataIn1 = 32'd7508
; 
32'd161333: dataIn1 = 32'd7509
; 
32'd161334: dataIn1 = 32'd6213
; 
32'd161335: dataIn1 = 32'd7435
; 
32'd161336: dataIn1 = 32'd7436
; 
32'd161337: dataIn1 = 32'd7438
; 
32'd161338: dataIn1 = 32'd7439
; 
32'd161339: dataIn1 = 32'd7463
; 
32'd161340: dataIn1 = 32'd7464
; 
32'd161341: dataIn1 = 32'd6214
; 
32'd161342: dataIn1 = 32'd7443
; 
32'd161343: dataIn1 = 32'd7444
; 
32'd161344: dataIn1 = 32'd7446
; 
32'd161345: dataIn1 = 32'd7448
; 
32'd161346: dataIn1 = 32'd7491
; 
32'd161347: dataIn1 = 32'd7492
; 
32'd161348: dataIn1 = 32'd6215
; 
32'd161349: dataIn1 = 32'd7442
; 
32'd161350: dataIn1 = 32'd7444
; 
32'd161351: dataIn1 = 32'd7445
; 
32'd161352: dataIn1 = 32'd7447
; 
32'd161353: dataIn1 = 32'd7468
; 
32'd161354: dataIn1 = 32'd7470
; 
32'd161355: dataIn1 = 32'd6216
; 
32'd161356: dataIn1 = 32'd7450
; 
32'd161357: dataIn1 = 32'd7451
; 
32'd161358: dataIn1 = 32'd7455
; 
32'd161359: dataIn1 = 32'd7457
; 
32'd161360: dataIn1 = 32'd7459
; 
32'd161361: dataIn1 = 32'd7460
; 
32'd161362: dataIn1 = 32'd6217
; 
32'd161363: dataIn1 = 32'd7449
; 
32'd161364: dataIn1 = 32'd7451
; 
32'd161365: dataIn1 = 32'd7453
; 
32'd161366: dataIn1 = 32'd7456
; 
32'd161367: dataIn1 = 32'd7463
; 
32'd161368: dataIn1 = 32'd7465
; 
32'd161369: dataIn1 = 32'd6218
; 
32'd161370: dataIn1 = 32'd7449
; 
32'd161371: dataIn1 = 32'd7450
; 
32'd161372: dataIn1 = 32'd7452
; 
32'd161373: dataIn1 = 32'd7454
; 
32'd161374: dataIn1 = 32'd7468
; 
32'd161375: dataIn1 = 32'd7469
; 
32'd161376: dataIn1 = 32'd6219
; 
32'd161377: dataIn1 = 32'd7458
; 
32'd161378: dataIn1 = 32'd7460
; 
32'd161379: dataIn1 = 32'd7462
; 
32'd161380: dataIn1 = 32'd8959
; 
32'd161381: dataIn1 = 32'd8960
; 
32'd161382: dataIn1 = 32'd8962
; 
32'd161383: dataIn1 = 32'd6220
; 
32'd161384: dataIn1 = 32'd7464
; 
32'd161385: dataIn1 = 32'd7465
; 
32'd161386: dataIn1 = 32'd7466
; 
32'd161387: dataIn1 = 32'd7467
; 
32'd161388: dataIn1 = 32'd8968
; 
32'd161389: dataIn1 = 32'd8969
; 
32'd161390: dataIn1 = 32'd6221
; 
32'd161391: dataIn1 = 32'd7474
; 
32'd161392: dataIn1 = 32'd7475
; 
32'd161393: dataIn1 = 32'd7479
; 
32'd161394: dataIn1 = 32'd7481
; 
32'd161395: dataIn1 = 32'd7483
; 
32'd161396: dataIn1 = 32'd7484
; 
32'd161397: dataIn1 = 32'd6222
; 
32'd161398: dataIn1 = 32'd7473
; 
32'd161399: dataIn1 = 32'd7475
; 
32'd161400: dataIn1 = 32'd7477
; 
32'd161401: dataIn1 = 32'd7480
; 
32'd161402: dataIn1 = 32'd7485
; 
32'd161403: dataIn1 = 32'd7487
; 
32'd161404: dataIn1 = 32'd6223
; 
32'd161405: dataIn1 = 32'd7473
; 
32'd161406: dataIn1 = 32'd7474
; 
32'd161407: dataIn1 = 32'd7476
; 
32'd161408: dataIn1 = 32'd7478
; 
32'd161409: dataIn1 = 32'd7490
; 
32'd161410: dataIn1 = 32'd7491
; 
32'd161411: dataIn1 = 32'd6224
; 
32'd161412: dataIn1 = 32'd7496
; 
32'd161413: dataIn1 = 32'd7497
; 
32'd161414: dataIn1 = 32'd7501
; 
32'd161415: dataIn1 = 32'd7503
; 
32'd161416: dataIn1 = 32'd7505
; 
32'd161417: dataIn1 = 32'd7506
; 
32'd161418: dataIn1 = 32'd6225
; 
32'd161419: dataIn1 = 32'd7495
; 
32'd161420: dataIn1 = 32'd7497
; 
32'd161421: dataIn1 = 32'd7499
; 
32'd161422: dataIn1 = 32'd7502
; 
32'd161423: dataIn1 = 32'd7507
; 
32'd161424: dataIn1 = 32'd7509
; 
32'd161425: dataIn1 = 32'd6226
; 
32'd161426: dataIn1 = 32'd6750
; 
32'd161427: dataIn1 = 32'd6751
; 
32'd161428: dataIn1 = 32'd7495
; 
32'd161429: dataIn1 = 32'd7496
; 
32'd161430: dataIn1 = 32'd7498
; 
32'd161431: dataIn1 = 32'd7500
; 
32'd161432: dataIn1 = 32'd6227
; 
32'd161433: dataIn1 = 32'd7507
; 
32'd161434: dataIn1 = 32'd7508
; 
32'd161435: dataIn1 = 32'd7510
; 
32'd161436: dataIn1 = 32'd7511
; 
32'd161437: dataIn1 = 32'd8970
; 
32'd161438: dataIn1 = 32'd8972
; 
32'd161439: dataIn1 = 32'd6228
; 
32'd161440: dataIn1 = 32'd7513
; 
32'd161441: dataIn1 = 32'd7514
; 
32'd161442: dataIn1 = 32'd7518
; 
32'd161443: dataIn1 = 32'd7520
; 
32'd161444: dataIn1 = 32'd7522
; 
32'd161445: dataIn1 = 32'd7523
; 
32'd161446: dataIn1 = 32'd6229
; 
32'd161447: dataIn1 = 32'd7512
; 
32'd161448: dataIn1 = 32'd7514
; 
32'd161449: dataIn1 = 32'd7516
; 
32'd161450: dataIn1 = 32'd7519
; 
32'd161451: dataIn1 = 32'd7528
; 
32'd161452: dataIn1 = 32'd7530
; 
32'd161453: dataIn1 = 32'd6230
; 
32'd161454: dataIn1 = 32'd7512
; 
32'd161455: dataIn1 = 32'd7513
; 
32'd161456: dataIn1 = 32'd7515
; 
32'd161457: dataIn1 = 32'd7517
; 
32'd161458: dataIn1 = 32'd7535
; 
32'd161459: dataIn1 = 32'd7536
; 
32'd161460: dataIn1 = 32'd6231
; 
32'd161461: dataIn1 = 32'd7521
; 
32'd161462: dataIn1 = 32'd7523
; 
32'd161463: dataIn1 = 32'd7525
; 
32'd161464: dataIn1 = 32'd7527
; 
32'd161465: dataIn1 = 32'd7590
; 
32'd161466: dataIn1 = 32'd7592
; 
32'd161467: dataIn1 = 32'd6232
; 
32'd161468: dataIn1 = 32'd7521
; 
32'd161469: dataIn1 = 32'd7522
; 
32'd161470: dataIn1 = 32'd7524
; 
32'd161471: dataIn1 = 32'd7526
; 
32'd161472: dataIn1 = 32'd7568
; 
32'd161473: dataIn1 = 32'd7569
; 
32'd161474: dataIn1 = 32'd6233
; 
32'd161475: dataIn1 = 32'd7529
; 
32'd161476: dataIn1 = 32'd7530
; 
32'd161477: dataIn1 = 32'd7533
; 
32'd161478: dataIn1 = 32'd7534
; 
32'd161479: dataIn1 = 32'd7596
; 
32'd161480: dataIn1 = 32'd7597
; 
32'd161481: dataIn1 = 32'd6234
; 
32'd161482: dataIn1 = 32'd7528
; 
32'd161483: dataIn1 = 32'd7529
; 
32'd161484: dataIn1 = 32'd7531
; 
32'd161485: dataIn1 = 32'd7532
; 
32'd161486: dataIn1 = 32'd7551
; 
32'd161487: dataIn1 = 32'd7552
; 
32'd161488: dataIn1 = 32'd6235
; 
32'd161489: dataIn1 = 32'd7536
; 
32'd161490: dataIn1 = 32'd7537
; 
32'd161491: dataIn1 = 32'd7539
; 
32'd161492: dataIn1 = 32'd7541
; 
32'd161493: dataIn1 = 32'd7579
; 
32'd161494: dataIn1 = 32'd7580
; 
32'd161495: dataIn1 = 32'd6236
; 
32'd161496: dataIn1 = 32'd7535
; 
32'd161497: dataIn1 = 32'd7537
; 
32'd161498: dataIn1 = 32'd7538
; 
32'd161499: dataIn1 = 32'd7540
; 
32'd161500: dataIn1 = 32'd7556
; 
32'd161501: dataIn1 = 32'd7558
; 
32'd161502: dataIn1 = 32'd6237
; 
32'd161503: dataIn1 = 32'd6752
; 
32'd161504: dataIn1 = 32'd6753
; 
32'd161505: dataIn1 = 32'd7543
; 
32'd161506: dataIn1 = 32'd7544
; 
32'd161507: dataIn1 = 32'd7548
; 
32'd161508: dataIn1 = 32'd7550
; 
32'd161509: dataIn1 = 32'd6238
; 
32'd161510: dataIn1 = 32'd7542
; 
32'd161511: dataIn1 = 32'd7544
; 
32'd161512: dataIn1 = 32'd7546
; 
32'd161513: dataIn1 = 32'd7549
; 
32'd161514: dataIn1 = 32'd7551
; 
32'd161515: dataIn1 = 32'd7553
; 
32'd161516: dataIn1 = 32'd6239
; 
32'd161517: dataIn1 = 32'd7542
; 
32'd161518: dataIn1 = 32'd7543
; 
32'd161519: dataIn1 = 32'd7545
; 
32'd161520: dataIn1 = 32'd7547
; 
32'd161521: dataIn1 = 32'd7556
; 
32'd161522: dataIn1 = 32'd7557
; 
32'd161523: dataIn1 = 32'd6240
; 
32'd161524: dataIn1 = 32'd7552
; 
32'd161525: dataIn1 = 32'd7553
; 
32'd161526: dataIn1 = 32'd7554
; 
32'd161527: dataIn1 = 32'd7555
; 
32'd161528: dataIn1 = 32'd9022
; 
32'd161529: dataIn1 = 32'd9023
; 
32'd161530: dataIn1 = 32'd6241
; 
32'd161531: dataIn1 = 32'd7560
; 
32'd161532: dataIn1 = 32'd7561
; 
32'd161533: dataIn1 = 32'd7565
; 
32'd161534: dataIn1 = 32'd7567
; 
32'd161535: dataIn1 = 32'd7569
; 
32'd161536: dataIn1 = 32'd7570
; 
32'd161537: dataIn1 = 32'd6242
; 
32'd161538: dataIn1 = 32'd7559
; 
32'd161539: dataIn1 = 32'd7561
; 
32'd161540: dataIn1 = 32'd7563
; 
32'd161541: dataIn1 = 32'd7566
; 
32'd161542: dataIn1 = 32'd7573
; 
32'd161543: dataIn1 = 32'd7575
; 
32'd161544: dataIn1 = 32'd6243
; 
32'd161545: dataIn1 = 32'd7559
; 
32'd161546: dataIn1 = 32'd7560
; 
32'd161547: dataIn1 = 32'd7562
; 
32'd161548: dataIn1 = 32'd7564
; 
32'd161549: dataIn1 = 32'd7578
; 
32'd161550: dataIn1 = 32'd7579
; 
32'd161551: dataIn1 = 32'd6244
; 
32'd161552: dataIn1 = 32'd7582
; 
32'd161553: dataIn1 = 32'd7583
; 
32'd161554: dataIn1 = 32'd7587
; 
32'd161555: dataIn1 = 32'd7589
; 
32'd161556: dataIn1 = 32'd7591
; 
32'd161557: dataIn1 = 32'd7592
; 
32'd161558: dataIn1 = 32'd6245
; 
32'd161559: dataIn1 = 32'd7581
; 
32'd161560: dataIn1 = 32'd7583
; 
32'd161561: dataIn1 = 32'd7585
; 
32'd161562: dataIn1 = 32'd7588
; 
32'd161563: dataIn1 = 32'd7595
; 
32'd161564: dataIn1 = 32'd7597
; 
32'd161565: dataIn1 = 32'd6246
; 
32'd161566: dataIn1 = 32'd7581
; 
32'd161567: dataIn1 = 32'd7582
; 
32'd161568: dataIn1 = 32'd7584
; 
32'd161569: dataIn1 = 32'd7586
; 
32'd161570: dataIn1 = 32'd7600
; 
32'd161571: dataIn1 = 32'd7601
; 
32'd161572: dataIn1 = 32'd6247
; 
32'd161573: dataIn1 = 32'd7595
; 
32'd161574: dataIn1 = 32'd7596
; 
32'd161575: dataIn1 = 32'd7598
; 
32'd161576: dataIn1 = 32'd7599
; 
32'd161577: dataIn1 = 32'd9012
; 
32'd161578: dataIn1 = 32'd9013
; 
32'd161579: dataIn1 = 32'd6248
; 
32'd161580: dataIn1 = 32'd7600
; 
32'd161581: dataIn1 = 32'd7602
; 
32'd161582: dataIn1 = 32'd7603
; 
32'd161583: dataIn1 = 32'd7605
; 
32'd161584: dataIn1 = 32'd9008
; 
32'd161585: dataIn1 = 32'd9010
; 
32'd161586: dataIn1 = 32'd6249
; 
32'd161587: dataIn1 = 32'd7608
; 
32'd161588: dataIn1 = 32'd7609
; 
32'd161589: dataIn1 = 32'd7613
; 
32'd161590: dataIn1 = 32'd7615
; 
32'd161591: dataIn1 = 32'd7617
; 
32'd161592: dataIn1 = 32'd7618
; 
32'd161593: dataIn1 = 32'd6250
; 
32'd161594: dataIn1 = 32'd6754
; 
32'd161595: dataIn1 = 32'd6755
; 
32'd161596: dataIn1 = 32'd7607
; 
32'd161597: dataIn1 = 32'd7609
; 
32'd161598: dataIn1 = 32'd7611
; 
32'd161599: dataIn1 = 32'd7614
; 
32'd161600: dataIn1 = 32'd6251
; 
32'd161601: dataIn1 = 32'd7607
; 
32'd161602: dataIn1 = 32'd7608
; 
32'd161603: dataIn1 = 32'd7610
; 
32'd161604: dataIn1 = 32'd7612
; 
32'd161605: dataIn1 = 32'd7623
; 
32'd161606: dataIn1 = 32'd7624
; 
32'd161607: dataIn1 = 32'd6252
; 
32'd161608: dataIn1 = 32'd7616
; 
32'd161609: dataIn1 = 32'd7618
; 
32'd161610: dataIn1 = 32'd7620
; 
32'd161611: dataIn1 = 32'd7622
; 
32'd161612: dataIn1 = 32'd7663
; 
32'd161613: dataIn1 = 32'd7665
; 
32'd161614: dataIn1 = 32'd6253
; 
32'd161615: dataIn1 = 32'd7616
; 
32'd161616: dataIn1 = 32'd7617
; 
32'd161617: dataIn1 = 32'd7619
; 
32'd161618: dataIn1 = 32'd7621
; 
32'd161619: dataIn1 = 32'd7646
; 
32'd161620: dataIn1 = 32'd7647
; 
32'd161621: dataIn1 = 32'd6254
; 
32'd161622: dataIn1 = 32'd7624
; 
32'd161623: dataIn1 = 32'd7625
; 
32'd161624: dataIn1 = 32'd7627
; 
32'd161625: dataIn1 = 32'd7629
; 
32'd161626: dataIn1 = 32'd7659
; 
32'd161627: dataIn1 = 32'd7660
; 
32'd161628: dataIn1 = 32'd6255
; 
32'd161629: dataIn1 = 32'd7623
; 
32'd161630: dataIn1 = 32'd7625
; 
32'd161631: dataIn1 = 32'd7626
; 
32'd161632: dataIn1 = 32'd7628
; 
32'd161633: dataIn1 = 32'd7630
; 
32'd161634: dataIn1 = 32'd7632
; 
32'd161635: dataIn1 = 32'd6256
; 
32'd161636: dataIn1 = 32'd7631
; 
32'd161637: dataIn1 = 32'd7632
; 
32'd161638: dataIn1 = 32'd7635
; 
32'd161639: dataIn1 = 32'd7636
; 
32'd161640: dataIn1 = 32'd7810
; 
32'd161641: dataIn1 = 32'd7811
; 
32'd161642: dataIn1 = 32'd6257
; 
32'd161643: dataIn1 = 32'd6756
; 
32'd161644: dataIn1 = 32'd6757
; 
32'd161645: dataIn1 = 32'd7630
; 
32'd161646: dataIn1 = 32'd7631
; 
32'd161647: dataIn1 = 32'd7633
; 
32'd161648: dataIn1 = 32'd7634
; 
32'd161649: dataIn1 = 32'd6258
; 
32'd161650: dataIn1 = 32'd7638
; 
32'd161651: dataIn1 = 32'd7639
; 
32'd161652: dataIn1 = 32'd7643
; 
32'd161653: dataIn1 = 32'd7645
; 
32'd161654: dataIn1 = 32'd7647
; 
32'd161655: dataIn1 = 32'd7648
; 
32'd161656: dataIn1 = 32'd6259
; 
32'd161657: dataIn1 = 32'd7637
; 
32'd161658: dataIn1 = 32'd7639
; 
32'd161659: dataIn1 = 32'd7641
; 
32'd161660: dataIn1 = 32'd7644
; 
32'd161661: dataIn1 = 32'd7651
; 
32'd161662: dataIn1 = 32'd7653
; 
32'd161663: dataIn1 = 32'd6260
; 
32'd161664: dataIn1 = 32'd7637
; 
32'd161665: dataIn1 = 32'd7638
; 
32'd161666: dataIn1 = 32'd7640
; 
32'd161667: dataIn1 = 32'd7642
; 
32'd161668: dataIn1 = 32'd7658
; 
32'd161669: dataIn1 = 32'd7659
; 
32'd161670: dataIn1 = 32'd6261
; 
32'd161671: dataIn1 = 32'd7646
; 
32'd161672: dataIn1 = 32'd7648
; 
32'd161673: dataIn1 = 32'd7649
; 
32'd161674: dataIn1 = 32'd7650
; 
32'd161675: dataIn1 = 32'd7735
; 
32'd161676: dataIn1 = 32'd7737
; 
32'd161677: dataIn1 = 32'd6262
; 
32'd161678: dataIn1 = 32'd7652
; 
32'd161679: dataIn1 = 32'd7653
; 
32'd161680: dataIn1 = 32'd7656
; 
32'd161681: dataIn1 = 32'd7657
; 
32'd161682: dataIn1 = 32'd7739
; 
32'd161683: dataIn1 = 32'd7740
; 
32'd161684: dataIn1 = 32'd6263
; 
32'd161685: dataIn1 = 32'd7651
; 
32'd161686: dataIn1 = 32'd7652
; 
32'd161687: dataIn1 = 32'd7654
; 
32'd161688: dataIn1 = 32'd7655
; 
32'd161689: dataIn1 = 32'd7826
; 
32'd161690: dataIn1 = 32'd7827
; 
32'd161691: dataIn1 = 32'd6264
; 
32'd161692: dataIn1 = 32'd7658
; 
32'd161693: dataIn1 = 32'd7660
; 
32'd161694: dataIn1 = 32'd7661
; 
32'd161695: dataIn1 = 32'd7662
; 
32'd161696: dataIn1 = 32'd7831
; 
32'd161697: dataIn1 = 32'd7833
; 
32'd161698: dataIn1 = 32'd6265
; 
32'd161699: dataIn1 = 32'd6758
; 
32'd161700: dataIn1 = 32'd6759
; 
32'd161701: dataIn1 = 32'd7664
; 
32'd161702: dataIn1 = 32'd7665
; 
32'd161703: dataIn1 = 32'd7668
; 
32'd161704: dataIn1 = 32'd7669
; 
32'd161705: dataIn1 = 32'd6266
; 
32'd161706: dataIn1 = 32'd7663
; 
32'd161707: dataIn1 = 32'd7664
; 
32'd161708: dataIn1 = 32'd7666
; 
32'd161709: dataIn1 = 32'd7667
; 
32'd161710: dataIn1 = 32'd7757
; 
32'd161711: dataIn1 = 32'd7758
; 
32'd161712: dataIn1 = 32'd6267
; 
32'd161713: dataIn1 = 32'd7671
; 
32'd161714: dataIn1 = 32'd7672
; 
32'd161715: dataIn1 = 32'd7676
; 
32'd161716: dataIn1 = 32'd7678
; 
32'd161717: dataIn1 = 32'd7680
; 
32'd161718: dataIn1 = 32'd7681
; 
32'd161719: dataIn1 = 32'd6268
; 
32'd161720: dataIn1 = 32'd7670
; 
32'd161721: dataIn1 = 32'd7672
; 
32'd161722: dataIn1 = 32'd7674
; 
32'd161723: dataIn1 = 32'd7677
; 
32'd161724: dataIn1 = 32'd7686
; 
32'd161725: dataIn1 = 32'd7688
; 
32'd161726: dataIn1 = 32'd6269
; 
32'd161727: dataIn1 = 32'd7670
; 
32'd161728: dataIn1 = 32'd7671
; 
32'd161729: dataIn1 = 32'd7673
; 
32'd161730: dataIn1 = 32'd7675
; 
32'd161731: dataIn1 = 32'd7693
; 
32'd161732: dataIn1 = 32'd7694
; 
32'd161733: dataIn1 = 32'd6270
; 
32'd161734: dataIn1 = 32'd7679
; 
32'd161735: dataIn1 = 32'd7681
; 
32'd161736: dataIn1 = 32'd7683
; 
32'd161737: dataIn1 = 32'd7685
; 
32'd161738: dataIn1 = 32'd7757
; 
32'd161739: dataIn1 = 32'd7759
; 
32'd161740: dataIn1 = 32'd6271
; 
32'd161741: dataIn1 = 32'd7679
; 
32'd161742: dataIn1 = 32'd7680
; 
32'd161743: dataIn1 = 32'd7682
; 
32'd161744: dataIn1 = 32'd7684
; 
32'd161745: dataIn1 = 32'd7735
; 
32'd161746: dataIn1 = 32'd7736
; 
32'd161747: dataIn1 = 32'd6272
; 
32'd161748: dataIn1 = 32'd7687
; 
32'd161749: dataIn1 = 32'd7688
; 
32'd161750: dataIn1 = 32'd7691
; 
32'd161751: dataIn1 = 32'd7692
; 
32'd161752: dataIn1 = 32'd7761
; 
32'd161753: dataIn1 = 32'd7762
; 
32'd161754: dataIn1 = 32'd6273
; 
32'd161755: dataIn1 = 32'd7686
; 
32'd161756: dataIn1 = 32'd7687
; 
32'd161757: dataIn1 = 32'd7689
; 
32'd161758: dataIn1 = 32'd7690
; 
32'd161759: dataIn1 = 32'd7716
; 
32'd161760: dataIn1 = 32'd7717
; 
32'd161761: dataIn1 = 32'd6274
; 
32'd161762: dataIn1 = 32'd7694
; 
32'd161763: dataIn1 = 32'd7695
; 
32'd161764: dataIn1 = 32'd7697
; 
32'd161765: dataIn1 = 32'd7699
; 
32'd161766: dataIn1 = 32'd7744
; 
32'd161767: dataIn1 = 32'd7745
; 
32'd161768: dataIn1 = 32'd6275
; 
32'd161769: dataIn1 = 32'd7693
; 
32'd161770: dataIn1 = 32'd7695
; 
32'd161771: dataIn1 = 32'd7696
; 
32'd161772: dataIn1 = 32'd7698
; 
32'd161773: dataIn1 = 32'd7721
; 
32'd161774: dataIn1 = 32'd7723
; 
32'd161775: dataIn1 = 32'd6276
; 
32'd161776: dataIn1 = 32'd7701
; 
32'd161777: dataIn1 = 32'd7702
; 
32'd161778: dataIn1 = 32'd7706
; 
32'd161779: dataIn1 = 32'd7708
; 
32'd161780: dataIn1 = 32'd7710
; 
32'd161781: dataIn1 = 32'd7711
; 
32'd161782: dataIn1 = 32'd6277
; 
32'd161783: dataIn1 = 32'd7700
; 
32'd161784: dataIn1 = 32'd7702
; 
32'd161785: dataIn1 = 32'd7704
; 
32'd161786: dataIn1 = 32'd7707
; 
32'd161787: dataIn1 = 32'd7716
; 
32'd161788: dataIn1 = 32'd7718
; 
32'd161789: dataIn1 = 32'd6278
; 
32'd161790: dataIn1 = 32'd7700
; 
32'd161791: dataIn1 = 32'd7701
; 
32'd161792: dataIn1 = 32'd7703
; 
32'd161793: dataIn1 = 32'd7705
; 
32'd161794: dataIn1 = 32'd7721
; 
32'd161795: dataIn1 = 32'd7722
; 
32'd161796: dataIn1 = 32'd6279
; 
32'd161797: dataIn1 = 32'd7709
; 
32'd161798: dataIn1 = 32'd7711
; 
32'd161799: dataIn1 = 32'd7713
; 
32'd161800: dataIn1 = 32'd7715
; 
32'd161801: dataIn1 = 32'd9008
; 
32'd161802: dataIn1 = 32'd9009
; 
32'd161803: dataIn1 = 32'd6280
; 
32'd161804: dataIn1 = 32'd7717
; 
32'd161805: dataIn1 = 32'd7718
; 
32'd161806: dataIn1 = 32'd7719
; 
32'd161807: dataIn1 = 32'd7720
; 
32'd161808: dataIn1 = 32'd9015
; 
32'd161809: dataIn1 = 32'd9016
; 
32'd161810: dataIn1 = 32'd6281
; 
32'd161811: dataIn1 = 32'd7727
; 
32'd161812: dataIn1 = 32'd7728
; 
32'd161813: dataIn1 = 32'd7732
; 
32'd161814: dataIn1 = 32'd7734
; 
32'd161815: dataIn1 = 32'd7736
; 
32'd161816: dataIn1 = 32'd7737
; 
32'd161817: dataIn1 = 32'd6282
; 
32'd161818: dataIn1 = 32'd7726
; 
32'd161819: dataIn1 = 32'd7728
; 
32'd161820: dataIn1 = 32'd7730
; 
32'd161821: dataIn1 = 32'd7733
; 
32'd161822: dataIn1 = 32'd7738
; 
32'd161823: dataIn1 = 32'd7740
; 
32'd161824: dataIn1 = 32'd6283
; 
32'd161825: dataIn1 = 32'd7726
; 
32'd161826: dataIn1 = 32'd7727
; 
32'd161827: dataIn1 = 32'd7729
; 
32'd161828: dataIn1 = 32'd7731
; 
32'd161829: dataIn1 = 32'd7743
; 
32'd161830: dataIn1 = 32'd7744
; 
32'd161831: dataIn1 = 32'd6284
; 
32'd161832: dataIn1 = 32'd7749
; 
32'd161833: dataIn1 = 32'd7750
; 
32'd161834: dataIn1 = 32'd7754
; 
32'd161835: dataIn1 = 32'd7756
; 
32'd161836: dataIn1 = 32'd7758
; 
32'd161837: dataIn1 = 32'd7759
; 
32'd161838: dataIn1 = 32'd6285
; 
32'd161839: dataIn1 = 32'd7748
; 
32'd161840: dataIn1 = 32'd7750
; 
32'd161841: dataIn1 = 32'd7752
; 
32'd161842: dataIn1 = 32'd7755
; 
32'd161843: dataIn1 = 32'd7760
; 
32'd161844: dataIn1 = 32'd7762
; 
32'd161845: dataIn1 = 32'd6286
; 
32'd161846: dataIn1 = 32'd6760
; 
32'd161847: dataIn1 = 32'd6761
; 
32'd161848: dataIn1 = 32'd7748
; 
32'd161849: dataIn1 = 32'd7749
; 
32'd161850: dataIn1 = 32'd7751
; 
32'd161851: dataIn1 = 32'd7753
; 
32'd161852: dataIn1 = 32'd6287
; 
32'd161853: dataIn1 = 32'd7760
; 
32'd161854: dataIn1 = 32'd7761
; 
32'd161855: dataIn1 = 32'd7763
; 
32'd161856: dataIn1 = 32'd7764
; 
32'd161857: dataIn1 = 32'd9017
; 
32'd161858: dataIn1 = 32'd9019
; 
32'd161859: dataIn1 = 32'd6288
; 
32'd161860: dataIn1 = 32'd7766
; 
32'd161861: dataIn1 = 32'd7767
; 
32'd161862: dataIn1 = 32'd7771
; 
32'd161863: dataIn1 = 32'd7773
; 
32'd161864: dataIn1 = 32'd7775
; 
32'd161865: dataIn1 = 32'd7776
; 
32'd161866: dataIn1 = 32'd6289
; 
32'd161867: dataIn1 = 32'd7765
; 
32'd161868: dataIn1 = 32'd7767
; 
32'd161869: dataIn1 = 32'd7769
; 
32'd161870: dataIn1 = 32'd7772
; 
32'd161871: dataIn1 = 32'd7781
; 
32'd161872: dataIn1 = 32'd7783
; 
32'd161873: dataIn1 = 32'd6290
; 
32'd161874: dataIn1 = 32'd7765
; 
32'd161875: dataIn1 = 32'd7766
; 
32'd161876: dataIn1 = 32'd7768
; 
32'd161877: dataIn1 = 32'd7770
; 
32'd161878: dataIn1 = 32'd7788
; 
32'd161879: dataIn1 = 32'd7789
; 
32'd161880: dataIn1 = 32'd6291
; 
32'd161881: dataIn1 = 32'd7774
; 
32'd161882: dataIn1 = 32'd7776
; 
32'd161883: dataIn1 = 32'd7778
; 
32'd161884: dataIn1 = 32'd7780
; 
32'd161885: dataIn1 = 32'd7843
; 
32'd161886: dataIn1 = 32'd7845
; 
32'd161887: dataIn1 = 32'd6292
; 
32'd161888: dataIn1 = 32'd7774
; 
32'd161889: dataIn1 = 32'd7775
; 
32'd161890: dataIn1 = 32'd7777
; 
32'd161891: dataIn1 = 32'd7779
; 
32'd161892: dataIn1 = 32'd7821
; 
32'd161893: dataIn1 = 32'd7822
; 
32'd161894: dataIn1 = 32'd6293
; 
32'd161895: dataIn1 = 32'd7782
; 
32'd161896: dataIn1 = 32'd7783
; 
32'd161897: dataIn1 = 32'd7786
; 
32'd161898: dataIn1 = 32'd7787
; 
32'd161899: dataIn1 = 32'd7849
; 
32'd161900: dataIn1 = 32'd7850
; 
32'd161901: dataIn1 = 32'd6294
; 
32'd161902: dataIn1 = 32'd7781
; 
32'd161903: dataIn1 = 32'd7782
; 
32'd161904: dataIn1 = 32'd7784
; 
32'd161905: dataIn1 = 32'd7785
; 
32'd161906: dataIn1 = 32'd7804
; 
32'd161907: dataIn1 = 32'd7805
; 
32'd161908: dataIn1 = 32'd6295
; 
32'd161909: dataIn1 = 32'd7789
; 
32'd161910: dataIn1 = 32'd7790
; 
32'd161911: dataIn1 = 32'd7792
; 
32'd161912: dataIn1 = 32'd7794
; 
32'd161913: dataIn1 = 32'd7832
; 
32'd161914: dataIn1 = 32'd7833
; 
32'd161915: dataIn1 = 32'd6296
; 
32'd161916: dataIn1 = 32'd7788
; 
32'd161917: dataIn1 = 32'd7790
; 
32'd161918: dataIn1 = 32'd7791
; 
32'd161919: dataIn1 = 32'd7793
; 
32'd161920: dataIn1 = 32'd7809
; 
32'd161921: dataIn1 = 32'd7811
; 
32'd161922: dataIn1 = 32'd6297
; 
32'd161923: dataIn1 = 32'd6762
; 
32'd161924: dataIn1 = 32'd6763
; 
32'd161925: dataIn1 = 32'd7796
; 
32'd161926: dataIn1 = 32'd7797
; 
32'd161927: dataIn1 = 32'd7801
; 
32'd161928: dataIn1 = 32'd7803
; 
32'd161929: dataIn1 = 32'd6298
; 
32'd161930: dataIn1 = 32'd7795
; 
32'd161931: dataIn1 = 32'd7797
; 
32'd161932: dataIn1 = 32'd7799
; 
32'd161933: dataIn1 = 32'd7802
; 
32'd161934: dataIn1 = 32'd7804
; 
32'd161935: dataIn1 = 32'd7806
; 
32'd161936: dataIn1 = 32'd6299
; 
32'd161937: dataIn1 = 32'd7795
; 
32'd161938: dataIn1 = 32'd7796
; 
32'd161939: dataIn1 = 32'd7798
; 
32'd161940: dataIn1 = 32'd7800
; 
32'd161941: dataIn1 = 32'd7809
; 
32'd161942: dataIn1 = 32'd7810
; 
32'd161943: dataIn1 = 32'd6300
; 
32'd161944: dataIn1 = 32'd7805
; 
32'd161945: dataIn1 = 32'd7806
; 
32'd161946: dataIn1 = 32'd7807
; 
32'd161947: dataIn1 = 32'd7808
; 
32'd161948: dataIn1 = 32'd9074
; 
32'd161949: dataIn1 = 32'd9075
; 
32'd161950: dataIn1 = 32'd6301
; 
32'd161951: dataIn1 = 32'd7813
; 
32'd161952: dataIn1 = 32'd7814
; 
32'd161953: dataIn1 = 32'd7818
; 
32'd161954: dataIn1 = 32'd7820
; 
32'd161955: dataIn1 = 32'd7822
; 
32'd161956: dataIn1 = 32'd7823
; 
32'd161957: dataIn1 = 32'd6302
; 
32'd161958: dataIn1 = 32'd7812
; 
32'd161959: dataIn1 = 32'd7814
; 
32'd161960: dataIn1 = 32'd7816
; 
32'd161961: dataIn1 = 32'd7819
; 
32'd161962: dataIn1 = 32'd7826
; 
32'd161963: dataIn1 = 32'd7828
; 
32'd161964: dataIn1 = 32'd6303
; 
32'd161965: dataIn1 = 32'd7812
; 
32'd161966: dataIn1 = 32'd7813
; 
32'd161967: dataIn1 = 32'd7815
; 
32'd161968: dataIn1 = 32'd7817
; 
32'd161969: dataIn1 = 32'd7831
; 
32'd161970: dataIn1 = 32'd7832
; 
32'd161971: dataIn1 = 32'd6304
; 
32'd161972: dataIn1 = 32'd7835
; 
32'd161973: dataIn1 = 32'd7836
; 
32'd161974: dataIn1 = 32'd7840
; 
32'd161975: dataIn1 = 32'd7842
; 
32'd161976: dataIn1 = 32'd7844
; 
32'd161977: dataIn1 = 32'd7845
; 
32'd161978: dataIn1 = 32'd6305
; 
32'd161979: dataIn1 = 32'd7834
; 
32'd161980: dataIn1 = 32'd7836
; 
32'd161981: dataIn1 = 32'd7838
; 
32'd161982: dataIn1 = 32'd7841
; 
32'd161983: dataIn1 = 32'd7848
; 
32'd161984: dataIn1 = 32'd7850
; 
32'd161985: dataIn1 = 32'd6306
; 
32'd161986: dataIn1 = 32'd7834
; 
32'd161987: dataIn1 = 32'd7835
; 
32'd161988: dataIn1 = 32'd7837
; 
32'd161989: dataIn1 = 32'd7839
; 
32'd161990: dataIn1 = 32'd7853
; 
32'd161991: dataIn1 = 32'd7854
; 
32'd161992: dataIn1 = 32'd6307
; 
32'd161993: dataIn1 = 32'd7848
; 
32'd161994: dataIn1 = 32'd7849
; 
32'd161995: dataIn1 = 32'd7851
; 
32'd161996: dataIn1 = 32'd7852
; 
32'd161997: dataIn1 = 32'd9064
; 
32'd161998: dataIn1 = 32'd9065
; 
32'd161999: dataIn1 = 32'd6308
; 
32'd162000: dataIn1 = 32'd7853
; 
32'd162001: dataIn1 = 32'd7855
; 
32'd162002: dataIn1 = 32'd7856
; 
32'd162003: dataIn1 = 32'd7858
; 
32'd162004: dataIn1 = 32'd9060
; 
32'd162005: dataIn1 = 32'd9062
; 
32'd162006: dataIn1 = 32'd6309
; 
32'd162007: dataIn1 = 32'd7861
; 
32'd162008: dataIn1 = 32'd7862
; 
32'd162009: dataIn1 = 32'd7866
; 
32'd162010: dataIn1 = 32'd7868
; 
32'd162011: dataIn1 = 32'd7870
; 
32'd162012: dataIn1 = 32'd7871
; 
32'd162013: dataIn1 = 32'd6310
; 
32'd162014: dataIn1 = 32'd6314
; 
32'd162015: dataIn1 = 32'd6315
; 
32'd162016: dataIn1 = 32'd7860
; 
32'd162017: dataIn1 = 32'd7862
; 
32'd162018: dataIn1 = 32'd7864
; 
32'd162019: dataIn1 = 32'd7867
; 
32'd162020: dataIn1 = 32'd6311
; 
32'd162021: dataIn1 = 32'd7860
; 
32'd162022: dataIn1 = 32'd7861
; 
32'd162023: dataIn1 = 32'd7863
; 
32'd162024: dataIn1 = 32'd7865
; 
32'd162025: dataIn1 = 32'd7876
; 
32'd162026: dataIn1 = 32'd7877
; 
32'd162027: dataIn1 = 32'd6312
; 
32'd162028: dataIn1 = 32'd7869
; 
32'd162029: dataIn1 = 32'd7871
; 
32'd162030: dataIn1 = 32'd7873
; 
32'd162031: dataIn1 = 32'd7875
; 
32'd162032: dataIn1 = 32'd7916
; 
32'd162033: dataIn1 = 32'd7918
; 
32'd162034: dataIn1 = 32'd6313
; 
32'd162035: dataIn1 = 32'd7869
; 
32'd162036: dataIn1 = 32'd7870
; 
32'd162037: dataIn1 = 32'd7872
; 
32'd162038: dataIn1 = 32'd7874
; 
32'd162039: dataIn1 = 32'd7899
; 
32'd162040: dataIn1 = 32'd7900
; 
32'd162041: dataIn1 = 32'd2715
; 
32'd162042: dataIn1 = 32'd5190
; 
32'd162043: dataIn1 = 32'd6310
; 
32'd162044: dataIn1 = 32'd6314
; 
32'd162045: dataIn1 = 32'd6315
; 
32'd162046: dataIn1 = 32'd6334
; 
32'd162047: dataIn1 = 32'd6335
; 
32'd162048: dataIn1 = 32'd7867
; 
32'd162049: dataIn1 = 32'd2715
; 
32'd162050: dataIn1 = 32'd5188
; 
32'd162051: dataIn1 = 32'd6310
; 
32'd162052: dataIn1 = 32'd6314
; 
32'd162053: dataIn1 = 32'd6315
; 
32'd162054: dataIn1 = 32'd6321
; 
32'd162055: dataIn1 = 32'd6322
; 
32'd162056: dataIn1 = 32'd7864
; 
32'd162057: dataIn1 = 32'd6316
; 
32'd162058: dataIn1 = 32'd7877
; 
32'd162059: dataIn1 = 32'd7878
; 
32'd162060: dataIn1 = 32'd7880
; 
32'd162061: dataIn1 = 32'd7882
; 
32'd162062: dataIn1 = 32'd7912
; 
32'd162063: dataIn1 = 32'd7913
; 
32'd162064: dataIn1 = 32'd6317
; 
32'd162065: dataIn1 = 32'd7876
; 
32'd162066: dataIn1 = 32'd7878
; 
32'd162067: dataIn1 = 32'd7879
; 
32'd162068: dataIn1 = 32'd7881
; 
32'd162069: dataIn1 = 32'd7883
; 
32'd162070: dataIn1 = 32'd7885
; 
32'd162071: dataIn1 = 32'd5191
; 
32'd162072: dataIn1 = 32'd5192
; 
32'd162073: dataIn1 = 32'd6318
; 
32'd162074: dataIn1 = 32'd6319
; 
32'd162075: dataIn1 = 32'd6320
; 
32'd162076: dataIn1 = 32'd6322
; 
32'd162077: dataIn1 = 32'd6324
; 
32'd162078: dataIn1 = 32'd7887
; 
32'd162079: dataIn1 = 32'd1127
; 
32'd162080: dataIn1 = 32'd5192
; 
32'd162081: dataIn1 = 32'd6318
; 
32'd162082: dataIn1 = 32'd6319
; 
32'd162083: dataIn1 = 32'd6320
; 
32'd162084: dataIn1 = 32'd6709
; 
32'd162085: dataIn1 = 32'd1127
; 
32'd162086: dataIn1 = 32'd5191
; 
32'd162087: dataIn1 = 32'd6318
; 
32'd162088: dataIn1 = 32'd6319
; 
32'd162089: dataIn1 = 32'd6320
; 
32'd162090: dataIn1 = 32'd6370
; 
32'd162091: dataIn1 = 32'd6373
; 
32'd162092: dataIn1 = 32'd8054
; 
32'd162093: dataIn1 = 32'd2715
; 
32'd162094: dataIn1 = 32'd5192
; 
32'd162095: dataIn1 = 32'd6315
; 
32'd162096: dataIn1 = 32'd6321
; 
32'd162097: dataIn1 = 32'd6322
; 
32'd162098: dataIn1 = 32'd6708
; 
32'd162099: dataIn1 = 32'd5188
; 
32'd162100: dataIn1 = 32'd5192
; 
32'd162101: dataIn1 = 32'd6315
; 
32'd162102: dataIn1 = 32'd6318
; 
32'd162103: dataIn1 = 32'd6321
; 
32'd162104: dataIn1 = 32'd6322
; 
32'd162105: dataIn1 = 32'd6324
; 
32'd162106: dataIn1 = 32'd7886
; 
32'd162107: dataIn1 = 32'd6323
; 
32'd162108: dataIn1 = 32'd7884
; 
32'd162109: dataIn1 = 32'd7885
; 
32'd162110: dataIn1 = 32'd7888
; 
32'd162111: dataIn1 = 32'd7889
; 
32'd162112: dataIn1 = 32'd8063
; 
32'd162113: dataIn1 = 32'd8064
; 
32'd162114: dataIn1 = 32'd6318
; 
32'd162115: dataIn1 = 32'd6322
; 
32'd162116: dataIn1 = 32'd6324
; 
32'd162117: dataIn1 = 32'd7883
; 
32'd162118: dataIn1 = 32'd7884
; 
32'd162119: dataIn1 = 32'd7886
; 
32'd162120: dataIn1 = 32'd7887
; 
32'd162121: dataIn1 = 32'd6325
; 
32'd162122: dataIn1 = 32'd7891
; 
32'd162123: dataIn1 = 32'd7892
; 
32'd162124: dataIn1 = 32'd7896
; 
32'd162125: dataIn1 = 32'd7898
; 
32'd162126: dataIn1 = 32'd7900
; 
32'd162127: dataIn1 = 32'd7901
; 
32'd162128: dataIn1 = 32'd6326
; 
32'd162129: dataIn1 = 32'd7890
; 
32'd162130: dataIn1 = 32'd7892
; 
32'd162131: dataIn1 = 32'd7894
; 
32'd162132: dataIn1 = 32'd7897
; 
32'd162133: dataIn1 = 32'd7904
; 
32'd162134: dataIn1 = 32'd7906
; 
32'd162135: dataIn1 = 32'd6327
; 
32'd162136: dataIn1 = 32'd7890
; 
32'd162137: dataIn1 = 32'd7891
; 
32'd162138: dataIn1 = 32'd7893
; 
32'd162139: dataIn1 = 32'd7895
; 
32'd162140: dataIn1 = 32'd7911
; 
32'd162141: dataIn1 = 32'd7912
; 
32'd162142: dataIn1 = 32'd6328
; 
32'd162143: dataIn1 = 32'd7899
; 
32'd162144: dataIn1 = 32'd7901
; 
32'd162145: dataIn1 = 32'd7902
; 
32'd162146: dataIn1 = 32'd7903
; 
32'd162147: dataIn1 = 32'd7988
; 
32'd162148: dataIn1 = 32'd7990
; 
32'd162149: dataIn1 = 32'd6329
; 
32'd162150: dataIn1 = 32'd7905
; 
32'd162151: dataIn1 = 32'd7906
; 
32'd162152: dataIn1 = 32'd7909
; 
32'd162153: dataIn1 = 32'd7910
; 
32'd162154: dataIn1 = 32'd7992
; 
32'd162155: dataIn1 = 32'd7993
; 
32'd162156: dataIn1 = 32'd6330
; 
32'd162157: dataIn1 = 32'd7904
; 
32'd162158: dataIn1 = 32'd7905
; 
32'd162159: dataIn1 = 32'd7907
; 
32'd162160: dataIn1 = 32'd7908
; 
32'd162161: dataIn1 = 32'd8079
; 
32'd162162: dataIn1 = 32'd8080
; 
32'd162163: dataIn1 = 32'd6331
; 
32'd162164: dataIn1 = 32'd7911
; 
32'd162165: dataIn1 = 32'd7913
; 
32'd162166: dataIn1 = 32'd7914
; 
32'd162167: dataIn1 = 32'd7915
; 
32'd162168: dataIn1 = 32'd8084
; 
32'd162169: dataIn1 = 32'd8086
; 
32'd162170: dataIn1 = 32'd6332
; 
32'd162171: dataIn1 = 32'd6334
; 
32'd162172: dataIn1 = 32'd6338
; 
32'd162173: dataIn1 = 32'd7917
; 
32'd162174: dataIn1 = 32'd7918
; 
32'd162175: dataIn1 = 32'd7921
; 
32'd162176: dataIn1 = 32'd7922
; 
32'd162177: dataIn1 = 32'd6333
; 
32'd162178: dataIn1 = 32'd7916
; 
32'd162179: dataIn1 = 32'd7917
; 
32'd162180: dataIn1 = 32'd7919
; 
32'd162181: dataIn1 = 32'd7920
; 
32'd162182: dataIn1 = 32'd8010
; 
32'd162183: dataIn1 = 32'd8011
; 
32'd162184: dataIn1 = 32'd5190
; 
32'd162185: dataIn1 = 32'd5195
; 
32'd162186: dataIn1 = 32'd6314
; 
32'd162187: dataIn1 = 32'd6332
; 
32'd162188: dataIn1 = 32'd6334
; 
32'd162189: dataIn1 = 32'd6335
; 
32'd162190: dataIn1 = 32'd6338
; 
32'd162191: dataIn1 = 32'd7922
; 
32'd162192: dataIn1 = 32'd2715
; 
32'd162193: dataIn1 = 32'd5195
; 
32'd162194: dataIn1 = 32'd6314
; 
32'd162195: dataIn1 = 32'd6334
; 
32'd162196: dataIn1 = 32'd6335
; 
32'd162197: dataIn1 = 32'd6711
; 
32'd162198: dataIn1 = 32'd1128
; 
32'd162199: dataIn1 = 32'd5196
; 
32'd162200: dataIn1 = 32'd6336
; 
32'd162201: dataIn1 = 32'd6337
; 
32'd162202: dataIn1 = 32'd6338
; 
32'd162203: dataIn1 = 32'd6358
; 
32'd162204: dataIn1 = 32'd6360
; 
32'd162205: dataIn1 = 32'd8006
; 
32'd162206: dataIn1 = 32'd1128
; 
32'd162207: dataIn1 = 32'd5195
; 
32'd162208: dataIn1 = 32'd6336
; 
32'd162209: dataIn1 = 32'd6337
; 
32'd162210: dataIn1 = 32'd6338
; 
32'd162211: dataIn1 = 32'd6710
; 
32'd162212: dataIn1 = 32'd5195
; 
32'd162213: dataIn1 = 32'd5196
; 
32'd162214: dataIn1 = 32'd6332
; 
32'd162215: dataIn1 = 32'd6334
; 
32'd162216: dataIn1 = 32'd6336
; 
32'd162217: dataIn1 = 32'd6337
; 
32'd162218: dataIn1 = 32'd6338
; 
32'd162219: dataIn1 = 32'd7921
; 
32'd162220: dataIn1 = 32'd6339
; 
32'd162221: dataIn1 = 32'd7924
; 
32'd162222: dataIn1 = 32'd7925
; 
32'd162223: dataIn1 = 32'd7929
; 
32'd162224: dataIn1 = 32'd7931
; 
32'd162225: dataIn1 = 32'd7933
; 
32'd162226: dataIn1 = 32'd7934
; 
32'd162227: dataIn1 = 32'd6340
; 
32'd162228: dataIn1 = 32'd7923
; 
32'd162229: dataIn1 = 32'd7925
; 
32'd162230: dataIn1 = 32'd7927
; 
32'd162231: dataIn1 = 32'd7930
; 
32'd162232: dataIn1 = 32'd7939
; 
32'd162233: dataIn1 = 32'd7941
; 
32'd162234: dataIn1 = 32'd6341
; 
32'd162235: dataIn1 = 32'd7923
; 
32'd162236: dataIn1 = 32'd7924
; 
32'd162237: dataIn1 = 32'd7926
; 
32'd162238: dataIn1 = 32'd7928
; 
32'd162239: dataIn1 = 32'd7946
; 
32'd162240: dataIn1 = 32'd7947
; 
32'd162241: dataIn1 = 32'd6342
; 
32'd162242: dataIn1 = 32'd7932
; 
32'd162243: dataIn1 = 32'd7934
; 
32'd162244: dataIn1 = 32'd7936
; 
32'd162245: dataIn1 = 32'd7938
; 
32'd162246: dataIn1 = 32'd8010
; 
32'd162247: dataIn1 = 32'd8012
; 
32'd162248: dataIn1 = 32'd6343
; 
32'd162249: dataIn1 = 32'd7932
; 
32'd162250: dataIn1 = 32'd7933
; 
32'd162251: dataIn1 = 32'd7935
; 
32'd162252: dataIn1 = 32'd7937
; 
32'd162253: dataIn1 = 32'd7988
; 
32'd162254: dataIn1 = 32'd7989
; 
32'd162255: dataIn1 = 32'd6344
; 
32'd162256: dataIn1 = 32'd7940
; 
32'd162257: dataIn1 = 32'd7941
; 
32'd162258: dataIn1 = 32'd7944
; 
32'd162259: dataIn1 = 32'd7945
; 
32'd162260: dataIn1 = 32'd8014
; 
32'd162261: dataIn1 = 32'd8015
; 
32'd162262: dataIn1 = 32'd6345
; 
32'd162263: dataIn1 = 32'd7939
; 
32'd162264: dataIn1 = 32'd7940
; 
32'd162265: dataIn1 = 32'd7942
; 
32'd162266: dataIn1 = 32'd7943
; 
32'd162267: dataIn1 = 32'd7969
; 
32'd162268: dataIn1 = 32'd7970
; 
32'd162269: dataIn1 = 32'd6346
; 
32'd162270: dataIn1 = 32'd7947
; 
32'd162271: dataIn1 = 32'd7948
; 
32'd162272: dataIn1 = 32'd7950
; 
32'd162273: dataIn1 = 32'd7952
; 
32'd162274: dataIn1 = 32'd7997
; 
32'd162275: dataIn1 = 32'd7998
; 
32'd162276: dataIn1 = 32'd6347
; 
32'd162277: dataIn1 = 32'd7946
; 
32'd162278: dataIn1 = 32'd7948
; 
32'd162279: dataIn1 = 32'd7949
; 
32'd162280: dataIn1 = 32'd7951
; 
32'd162281: dataIn1 = 32'd7974
; 
32'd162282: dataIn1 = 32'd7976
; 
32'd162283: dataIn1 = 32'd6348
; 
32'd162284: dataIn1 = 32'd7954
; 
32'd162285: dataIn1 = 32'd7955
; 
32'd162286: dataIn1 = 32'd7959
; 
32'd162287: dataIn1 = 32'd7961
; 
32'd162288: dataIn1 = 32'd7963
; 
32'd162289: dataIn1 = 32'd7964
; 
32'd162290: dataIn1 = 32'd6349
; 
32'd162291: dataIn1 = 32'd7953
; 
32'd162292: dataIn1 = 32'd7955
; 
32'd162293: dataIn1 = 32'd7957
; 
32'd162294: dataIn1 = 32'd7960
; 
32'd162295: dataIn1 = 32'd7969
; 
32'd162296: dataIn1 = 32'd7971
; 
32'd162297: dataIn1 = 32'd6350
; 
32'd162298: dataIn1 = 32'd7953
; 
32'd162299: dataIn1 = 32'd7954
; 
32'd162300: dataIn1 = 32'd7956
; 
32'd162301: dataIn1 = 32'd7958
; 
32'd162302: dataIn1 = 32'd7974
; 
32'd162303: dataIn1 = 32'd7975
; 
32'd162304: dataIn1 = 32'd6351
; 
32'd162305: dataIn1 = 32'd7962
; 
32'd162306: dataIn1 = 32'd7964
; 
32'd162307: dataIn1 = 32'd7966
; 
32'd162308: dataIn1 = 32'd7968
; 
32'd162309: dataIn1 = 32'd9060
; 
32'd162310: dataIn1 = 32'd9061
; 
32'd162311: dataIn1 = 32'd6352
; 
32'd162312: dataIn1 = 32'd7970
; 
32'd162313: dataIn1 = 32'd7971
; 
32'd162314: dataIn1 = 32'd7972
; 
32'd162315: dataIn1 = 32'd7973
; 
32'd162316: dataIn1 = 32'd9067
; 
32'd162317: dataIn1 = 32'd9068
; 
32'd162318: dataIn1 = 32'd6353
; 
32'd162319: dataIn1 = 32'd7980
; 
32'd162320: dataIn1 = 32'd7981
; 
32'd162321: dataIn1 = 32'd7985
; 
32'd162322: dataIn1 = 32'd7987
; 
32'd162323: dataIn1 = 32'd7989
; 
32'd162324: dataIn1 = 32'd7990
; 
32'd162325: dataIn1 = 32'd6354
; 
32'd162326: dataIn1 = 32'd7979
; 
32'd162327: dataIn1 = 32'd7981
; 
32'd162328: dataIn1 = 32'd7983
; 
32'd162329: dataIn1 = 32'd7986
; 
32'd162330: dataIn1 = 32'd7991
; 
32'd162331: dataIn1 = 32'd7993
; 
32'd162332: dataIn1 = 32'd6355
; 
32'd162333: dataIn1 = 32'd7979
; 
32'd162334: dataIn1 = 32'd7980
; 
32'd162335: dataIn1 = 32'd7982
; 
32'd162336: dataIn1 = 32'd7984
; 
32'd162337: dataIn1 = 32'd7996
; 
32'd162338: dataIn1 = 32'd7997
; 
32'd162339: dataIn1 = 32'd6356
; 
32'd162340: dataIn1 = 32'd8002
; 
32'd162341: dataIn1 = 32'd8003
; 
32'd162342: dataIn1 = 32'd8007
; 
32'd162343: dataIn1 = 32'd8009
; 
32'd162344: dataIn1 = 32'd8011
; 
32'd162345: dataIn1 = 32'd8012
; 
32'd162346: dataIn1 = 32'd6357
; 
32'd162347: dataIn1 = 32'd8001
; 
32'd162348: dataIn1 = 32'd8003
; 
32'd162349: dataIn1 = 32'd8005
; 
32'd162350: dataIn1 = 32'd8008
; 
32'd162351: dataIn1 = 32'd8013
; 
32'd162352: dataIn1 = 32'd8015
; 
32'd162353: dataIn1 = 32'd6336
; 
32'd162354: dataIn1 = 32'd6358
; 
32'd162355: dataIn1 = 32'd6360
; 
32'd162356: dataIn1 = 32'd8001
; 
32'd162357: dataIn1 = 32'd8002
; 
32'd162358: dataIn1 = 32'd8004
; 
32'd162359: dataIn1 = 32'd8006
; 
32'd162360: dataIn1 = 32'd6359
; 
32'd162361: dataIn1 = 32'd8013
; 
32'd162362: dataIn1 = 32'd8014
; 
32'd162363: dataIn1 = 32'd8016
; 
32'd162364: dataIn1 = 32'd8017
; 
32'd162365: dataIn1 = 32'd9069
; 
32'd162366: dataIn1 = 32'd9071
; 
32'd162367: dataIn1 = 32'd1128
; 
32'd162368: dataIn1 = 32'd5201
; 
32'd162369: dataIn1 = 32'd6336
; 
32'd162370: dataIn1 = 32'd6358
; 
32'd162371: dataIn1 = 32'd6360
; 
32'd162372: dataIn1 = 32'd6637
; 
32'd162373: dataIn1 = 32'd6638
; 
32'd162374: dataIn1 = 32'd8004
; 
32'd162375: dataIn1 = 32'd6361
; 
32'd162376: dataIn1 = 32'd8019
; 
32'd162377: dataIn1 = 32'd8020
; 
32'd162378: dataIn1 = 32'd8024
; 
32'd162379: dataIn1 = 32'd8026
; 
32'd162380: dataIn1 = 32'd8028
; 
32'd162381: dataIn1 = 32'd8029
; 
32'd162382: dataIn1 = 32'd6362
; 
32'd162383: dataIn1 = 32'd8018
; 
32'd162384: dataIn1 = 32'd8020
; 
32'd162385: dataIn1 = 32'd8022
; 
32'd162386: dataIn1 = 32'd8025
; 
32'd162387: dataIn1 = 32'd8034
; 
32'd162388: dataIn1 = 32'd8036
; 
32'd162389: dataIn1 = 32'd6363
; 
32'd162390: dataIn1 = 32'd8018
; 
32'd162391: dataIn1 = 32'd8019
; 
32'd162392: dataIn1 = 32'd8021
; 
32'd162393: dataIn1 = 32'd8023
; 
32'd162394: dataIn1 = 32'd8041
; 
32'd162395: dataIn1 = 32'd8042
; 
32'd162396: dataIn1 = 32'd6364
; 
32'd162397: dataIn1 = 32'd8027
; 
32'd162398: dataIn1 = 32'd8029
; 
32'd162399: dataIn1 = 32'd8031
; 
32'd162400: dataIn1 = 32'd8033
; 
32'd162401: dataIn1 = 32'd8096
; 
32'd162402: dataIn1 = 32'd8098
; 
32'd162403: dataIn1 = 32'd6365
; 
32'd162404: dataIn1 = 32'd8027
; 
32'd162405: dataIn1 = 32'd8028
; 
32'd162406: dataIn1 = 32'd8030
; 
32'd162407: dataIn1 = 32'd8032
; 
32'd162408: dataIn1 = 32'd8074
; 
32'd162409: dataIn1 = 32'd8075
; 
32'd162410: dataIn1 = 32'd6366
; 
32'd162411: dataIn1 = 32'd8035
; 
32'd162412: dataIn1 = 32'd8036
; 
32'd162413: dataIn1 = 32'd8039
; 
32'd162414: dataIn1 = 32'd8040
; 
32'd162415: dataIn1 = 32'd8102
; 
32'd162416: dataIn1 = 32'd8103
; 
32'd162417: dataIn1 = 32'd6367
; 
32'd162418: dataIn1 = 32'd8034
; 
32'd162419: dataIn1 = 32'd8035
; 
32'd162420: dataIn1 = 32'd8037
; 
32'd162421: dataIn1 = 32'd8038
; 
32'd162422: dataIn1 = 32'd8057
; 
32'd162423: dataIn1 = 32'd8058
; 
32'd162424: dataIn1 = 32'd6368
; 
32'd162425: dataIn1 = 32'd8042
; 
32'd162426: dataIn1 = 32'd8043
; 
32'd162427: dataIn1 = 32'd8045
; 
32'd162428: dataIn1 = 32'd8047
; 
32'd162429: dataIn1 = 32'd8085
; 
32'd162430: dataIn1 = 32'd8086
; 
32'd162431: dataIn1 = 32'd6369
; 
32'd162432: dataIn1 = 32'd8041
; 
32'd162433: dataIn1 = 32'd8043
; 
32'd162434: dataIn1 = 32'd8044
; 
32'd162435: dataIn1 = 32'd8046
; 
32'd162436: dataIn1 = 32'd8062
; 
32'd162437: dataIn1 = 32'd8064
; 
32'd162438: dataIn1 = 32'd6320
; 
32'd162439: dataIn1 = 32'd6370
; 
32'd162440: dataIn1 = 32'd6373
; 
32'd162441: dataIn1 = 32'd8049
; 
32'd162442: dataIn1 = 32'd8050
; 
32'd162443: dataIn1 = 32'd8054
; 
32'd162444: dataIn1 = 32'd8056
; 
32'd162445: dataIn1 = 32'd6371
; 
32'd162446: dataIn1 = 32'd8048
; 
32'd162447: dataIn1 = 32'd8050
; 
32'd162448: dataIn1 = 32'd8052
; 
32'd162449: dataIn1 = 32'd8055
; 
32'd162450: dataIn1 = 32'd8057
; 
32'd162451: dataIn1 = 32'd8059
; 
32'd162452: dataIn1 = 32'd6372
; 
32'd162453: dataIn1 = 32'd8048
; 
32'd162454: dataIn1 = 32'd8049
; 
32'd162455: dataIn1 = 32'd8051
; 
32'd162456: dataIn1 = 32'd8053
; 
32'd162457: dataIn1 = 32'd8062
; 
32'd162458: dataIn1 = 32'd8063
; 
32'd162459: dataIn1 = 32'd1127
; 
32'd162460: dataIn1 = 32'd5205
; 
32'd162461: dataIn1 = 32'd6320
; 
32'd162462: dataIn1 = 32'd6370
; 
32'd162463: dataIn1 = 32'd6373
; 
32'd162464: dataIn1 = 32'd6659
; 
32'd162465: dataIn1 = 32'd6660
; 
32'd162466: dataIn1 = 32'd8056
; 
32'd162467: dataIn1 = 32'd6374
; 
32'd162468: dataIn1 = 32'd8058
; 
32'd162469: dataIn1 = 32'd8059
; 
32'd162470: dataIn1 = 32'd8060
; 
32'd162471: dataIn1 = 32'd8061
; 
32'd162472: dataIn1 = 32'd9125
; 
32'd162473: dataIn1 = 32'd9126
; 
32'd162474: dataIn1 = 32'd6375
; 
32'd162475: dataIn1 = 32'd8066
; 
32'd162476: dataIn1 = 32'd8067
; 
32'd162477: dataIn1 = 32'd8071
; 
32'd162478: dataIn1 = 32'd8073
; 
32'd162479: dataIn1 = 32'd8075
; 
32'd162480: dataIn1 = 32'd8076
; 
32'd162481: dataIn1 = 32'd6376
; 
32'd162482: dataIn1 = 32'd8065
; 
32'd162483: dataIn1 = 32'd8067
; 
32'd162484: dataIn1 = 32'd8069
; 
32'd162485: dataIn1 = 32'd8072
; 
32'd162486: dataIn1 = 32'd8079
; 
32'd162487: dataIn1 = 32'd8081
; 
32'd162488: dataIn1 = 32'd6377
; 
32'd162489: dataIn1 = 32'd8065
; 
32'd162490: dataIn1 = 32'd8066
; 
32'd162491: dataIn1 = 32'd8068
; 
32'd162492: dataIn1 = 32'd8070
; 
32'd162493: dataIn1 = 32'd8084
; 
32'd162494: dataIn1 = 32'd8085
; 
32'd162495: dataIn1 = 32'd6378
; 
32'd162496: dataIn1 = 32'd8088
; 
32'd162497: dataIn1 = 32'd8089
; 
32'd162498: dataIn1 = 32'd8093
; 
32'd162499: dataIn1 = 32'd8095
; 
32'd162500: dataIn1 = 32'd8097
; 
32'd162501: dataIn1 = 32'd8098
; 
32'd162502: dataIn1 = 32'd6379
; 
32'd162503: dataIn1 = 32'd8087
; 
32'd162504: dataIn1 = 32'd8089
; 
32'd162505: dataIn1 = 32'd8091
; 
32'd162506: dataIn1 = 32'd8094
; 
32'd162507: dataIn1 = 32'd8101
; 
32'd162508: dataIn1 = 32'd8103
; 
32'd162509: dataIn1 = 32'd6380
; 
32'd162510: dataIn1 = 32'd8087
; 
32'd162511: dataIn1 = 32'd8088
; 
32'd162512: dataIn1 = 32'd8090
; 
32'd162513: dataIn1 = 32'd8092
; 
32'd162514: dataIn1 = 32'd8106
; 
32'd162515: dataIn1 = 32'd8107
; 
32'd162516: dataIn1 = 32'd6381
; 
32'd162517: dataIn1 = 32'd8101
; 
32'd162518: dataIn1 = 32'd8102
; 
32'd162519: dataIn1 = 32'd8104
; 
32'd162520: dataIn1 = 32'd8105
; 
32'd162521: dataIn1 = 32'd9115
; 
32'd162522: dataIn1 = 32'd9116
; 
32'd162523: dataIn1 = 32'd6382
; 
32'd162524: dataIn1 = 32'd8106
; 
32'd162525: dataIn1 = 32'd8108
; 
32'd162526: dataIn1 = 32'd8109
; 
32'd162527: dataIn1 = 32'd8111
; 
32'd162528: dataIn1 = 32'd9111
; 
32'd162529: dataIn1 = 32'd9113
; 
32'd162530: dataIn1 = 32'd6383
; 
32'd162531: dataIn1 = 32'd8114
; 
32'd162532: dataIn1 = 32'd8115
; 
32'd162533: dataIn1 = 32'd8119
; 
32'd162534: dataIn1 = 32'd8121
; 
32'd162535: dataIn1 = 32'd8123
; 
32'd162536: dataIn1 = 32'd8124
; 
32'd162537: dataIn1 = 32'd6384
; 
32'd162538: dataIn1 = 32'd6388
; 
32'd162539: dataIn1 = 32'd6389
; 
32'd162540: dataIn1 = 32'd8113
; 
32'd162541: dataIn1 = 32'd8115
; 
32'd162542: dataIn1 = 32'd8117
; 
32'd162543: dataIn1 = 32'd8120
; 
32'd162544: dataIn1 = 32'd6385
; 
32'd162545: dataIn1 = 32'd8113
; 
32'd162546: dataIn1 = 32'd8114
; 
32'd162547: dataIn1 = 32'd8116
; 
32'd162548: dataIn1 = 32'd8118
; 
32'd162549: dataIn1 = 32'd8129
; 
32'd162550: dataIn1 = 32'd8130
; 
32'd162551: dataIn1 = 32'd6386
; 
32'd162552: dataIn1 = 32'd8122
; 
32'd162553: dataIn1 = 32'd8124
; 
32'd162554: dataIn1 = 32'd8126
; 
32'd162555: dataIn1 = 32'd8128
; 
32'd162556: dataIn1 = 32'd8169
; 
32'd162557: dataIn1 = 32'd8171
; 
32'd162558: dataIn1 = 32'd6387
; 
32'd162559: dataIn1 = 32'd8122
; 
32'd162560: dataIn1 = 32'd8123
; 
32'd162561: dataIn1 = 32'd8125
; 
32'd162562: dataIn1 = 32'd8127
; 
32'd162563: dataIn1 = 32'd8152
; 
32'd162564: dataIn1 = 32'd8153
; 
32'd162565: dataIn1 = 32'd2720
; 
32'd162566: dataIn1 = 32'd5209
; 
32'd162567: dataIn1 = 32'd6384
; 
32'd162568: dataIn1 = 32'd6388
; 
32'd162569: dataIn1 = 32'd6389
; 
32'd162570: dataIn1 = 32'd6408
; 
32'd162571: dataIn1 = 32'd6409
; 
32'd162572: dataIn1 = 32'd8120
; 
32'd162573: dataIn1 = 32'd2720
; 
32'd162574: dataIn1 = 32'd5207
; 
32'd162575: dataIn1 = 32'd6384
; 
32'd162576: dataIn1 = 32'd6388
; 
32'd162577: dataIn1 = 32'd6389
; 
32'd162578: dataIn1 = 32'd6393
; 
32'd162579: dataIn1 = 32'd6397
; 
32'd162580: dataIn1 = 32'd8117
; 
32'd162581: dataIn1 = 32'd9765
; 
32'd162582: dataIn1 = 32'd6390
; 
32'd162583: dataIn1 = 32'd8130
; 
32'd162584: dataIn1 = 32'd8131
; 
32'd162585: dataIn1 = 32'd8133
; 
32'd162586: dataIn1 = 32'd8135
; 
32'd162587: dataIn1 = 32'd8165
; 
32'd162588: dataIn1 = 32'd8166
; 
32'd162589: dataIn1 = 32'd6391
; 
32'd162590: dataIn1 = 32'd8129
; 
32'd162591: dataIn1 = 32'd8131
; 
32'd162592: dataIn1 = 32'd8132
; 
32'd162593: dataIn1 = 32'd8134
; 
32'd162594: dataIn1 = 32'd8136
; 
32'd162595: dataIn1 = 32'd8138
; 
32'd162596: dataIn1 = 32'd6392
; 
32'd162597: dataIn1 = 32'd9736
; 
32'd162598: dataIn1 = 32'd9737
; 
32'd162599: dataIn1 = 32'd9739
; 
32'd162600: dataIn1 = 32'd9741
; 
32'd162601: dataIn1 = 32'd9766
; 
32'd162602: dataIn1 = 32'd10279
; 
32'd162603: dataIn1 = 32'd6389
; 
32'd162604: dataIn1 = 32'd6393
; 
32'd162605: dataIn1 = 32'd6397
; 
32'd162606: dataIn1 = 32'd9735
; 
32'd162607: dataIn1 = 32'd9737
; 
32'd162608: dataIn1 = 32'd9738
; 
32'd162609: dataIn1 = 32'd9765
; 
32'd162610: dataIn1 = 32'd6394
; 
32'd162611: dataIn1 = 32'd8136
; 
32'd162612: dataIn1 = 32'd8137
; 
32'd162613: dataIn1 = 32'd8139
; 
32'd162614: dataIn1 = 32'd8140
; 
32'd162615: dataIn1 = 32'd9735
; 
32'd162616: dataIn1 = 32'd9736
; 
32'd162617: dataIn1 = 32'd1129
; 
32'd162618: dataIn1 = 32'd6395
; 
32'd162619: dataIn1 = 32'd9740
; 
32'd162620: dataIn1 = 32'd9741
; 
32'd162621: dataIn1 = 32'd10138
; 
32'd162622: dataIn1 = 32'd10140
; 
32'd162623: dataIn1 = 32'd10282
; 
32'd162624: dataIn1 = 32'd1129
; 
32'd162625: dataIn1 = 32'd6396
; 
32'd162626: dataIn1 = 32'd6443
; 
32'd162627: dataIn1 = 32'd10278
; 
32'd162628: dataIn1 = 32'd10279
; 
32'd162629: dataIn1 = 32'd10280
; 
32'd162630: dataIn1 = 32'd10282
; 
32'd162631: dataIn1 = 32'd2720
; 
32'd162632: dataIn1 = 32'd5211
; 
32'd162633: dataIn1 = 32'd6389
; 
32'd162634: dataIn1 = 32'd6393
; 
32'd162635: dataIn1 = 32'd6397
; 
32'd162636: dataIn1 = 32'd9738
; 
32'd162637: dataIn1 = 32'd9748
; 
32'd162638: dataIn1 = 32'd9776
; 
32'd162639: dataIn1 = 32'd6398
; 
32'd162640: dataIn1 = 32'd8137
; 
32'd162641: dataIn1 = 32'd8138
; 
32'd162642: dataIn1 = 32'd8141
; 
32'd162643: dataIn1 = 32'd8142
; 
32'd162644: dataIn1 = 32'd8315
; 
32'd162645: dataIn1 = 32'd8316
; 
32'd162646: dataIn1 = 32'd6399
; 
32'd162647: dataIn1 = 32'd8144
; 
32'd162648: dataIn1 = 32'd8145
; 
32'd162649: dataIn1 = 32'd8149
; 
32'd162650: dataIn1 = 32'd8151
; 
32'd162651: dataIn1 = 32'd8153
; 
32'd162652: dataIn1 = 32'd8154
; 
32'd162653: dataIn1 = 32'd6400
; 
32'd162654: dataIn1 = 32'd8143
; 
32'd162655: dataIn1 = 32'd8145
; 
32'd162656: dataIn1 = 32'd8147
; 
32'd162657: dataIn1 = 32'd8150
; 
32'd162658: dataIn1 = 32'd8157
; 
32'd162659: dataIn1 = 32'd8159
; 
32'd162660: dataIn1 = 32'd6401
; 
32'd162661: dataIn1 = 32'd8143
; 
32'd162662: dataIn1 = 32'd8144
; 
32'd162663: dataIn1 = 32'd8146
; 
32'd162664: dataIn1 = 32'd8148
; 
32'd162665: dataIn1 = 32'd8164
; 
32'd162666: dataIn1 = 32'd8165
; 
32'd162667: dataIn1 = 32'd6402
; 
32'd162668: dataIn1 = 32'd8152
; 
32'd162669: dataIn1 = 32'd8154
; 
32'd162670: dataIn1 = 32'd8155
; 
32'd162671: dataIn1 = 32'd8156
; 
32'd162672: dataIn1 = 32'd8241
; 
32'd162673: dataIn1 = 32'd8243
; 
32'd162674: dataIn1 = 32'd6403
; 
32'd162675: dataIn1 = 32'd8158
; 
32'd162676: dataIn1 = 32'd8159
; 
32'd162677: dataIn1 = 32'd8162
; 
32'd162678: dataIn1 = 32'd8163
; 
32'd162679: dataIn1 = 32'd8245
; 
32'd162680: dataIn1 = 32'd8246
; 
32'd162681: dataIn1 = 32'd6404
; 
32'd162682: dataIn1 = 32'd8157
; 
32'd162683: dataIn1 = 32'd8158
; 
32'd162684: dataIn1 = 32'd8160
; 
32'd162685: dataIn1 = 32'd8161
; 
32'd162686: dataIn1 = 32'd8331
; 
32'd162687: dataIn1 = 32'd8332
; 
32'd162688: dataIn1 = 32'd6405
; 
32'd162689: dataIn1 = 32'd8164
; 
32'd162690: dataIn1 = 32'd8166
; 
32'd162691: dataIn1 = 32'd8167
; 
32'd162692: dataIn1 = 32'd8168
; 
32'd162693: dataIn1 = 32'd8336
; 
32'd162694: dataIn1 = 32'd8338
; 
32'd162695: dataIn1 = 32'd6406
; 
32'd162696: dataIn1 = 32'd6408
; 
32'd162697: dataIn1 = 32'd6714
; 
32'd162698: dataIn1 = 32'd8170
; 
32'd162699: dataIn1 = 32'd8171
; 
32'd162700: dataIn1 = 32'd8174
; 
32'd162701: dataIn1 = 32'd8175
; 
32'd162702: dataIn1 = 32'd6407
; 
32'd162703: dataIn1 = 32'd8169
; 
32'd162704: dataIn1 = 32'd8170
; 
32'd162705: dataIn1 = 32'd8172
; 
32'd162706: dataIn1 = 32'd8173
; 
32'd162707: dataIn1 = 32'd8263
; 
32'd162708: dataIn1 = 32'd8264
; 
32'd162709: dataIn1 = 32'd5209
; 
32'd162710: dataIn1 = 32'd5214
; 
32'd162711: dataIn1 = 32'd6388
; 
32'd162712: dataIn1 = 32'd6406
; 
32'd162713: dataIn1 = 32'd6408
; 
32'd162714: dataIn1 = 32'd6409
; 
32'd162715: dataIn1 = 32'd6714
; 
32'd162716: dataIn1 = 32'd8175
; 
32'd162717: dataIn1 = 32'd2720
; 
32'd162718: dataIn1 = 32'd5214
; 
32'd162719: dataIn1 = 32'd6388
; 
32'd162720: dataIn1 = 32'd6408
; 
32'd162721: dataIn1 = 32'd6409
; 
32'd162722: dataIn1 = 32'd6716
; 
32'd162723: dataIn1 = 32'd6410
; 
32'd162724: dataIn1 = 32'd8177
; 
32'd162725: dataIn1 = 32'd8178
; 
32'd162726: dataIn1 = 32'd8182
; 
32'd162727: dataIn1 = 32'd8184
; 
32'd162728: dataIn1 = 32'd8186
; 
32'd162729: dataIn1 = 32'd8187
; 
32'd162730: dataIn1 = 32'd6411
; 
32'd162731: dataIn1 = 32'd8176
; 
32'd162732: dataIn1 = 32'd8178
; 
32'd162733: dataIn1 = 32'd8180
; 
32'd162734: dataIn1 = 32'd8183
; 
32'd162735: dataIn1 = 32'd8192
; 
32'd162736: dataIn1 = 32'd8194
; 
32'd162737: dataIn1 = 32'd6412
; 
32'd162738: dataIn1 = 32'd8176
; 
32'd162739: dataIn1 = 32'd8177
; 
32'd162740: dataIn1 = 32'd8179
; 
32'd162741: dataIn1 = 32'd8181
; 
32'd162742: dataIn1 = 32'd8199
; 
32'd162743: dataIn1 = 32'd8200
; 
32'd162744: dataIn1 = 32'd6413
; 
32'd162745: dataIn1 = 32'd8185
; 
32'd162746: dataIn1 = 32'd8187
; 
32'd162747: dataIn1 = 32'd8189
; 
32'd162748: dataIn1 = 32'd8191
; 
32'd162749: dataIn1 = 32'd8263
; 
32'd162750: dataIn1 = 32'd8265
; 
32'd162751: dataIn1 = 32'd6414
; 
32'd162752: dataIn1 = 32'd8185
; 
32'd162753: dataIn1 = 32'd8186
; 
32'd162754: dataIn1 = 32'd8188
; 
32'd162755: dataIn1 = 32'd8190
; 
32'd162756: dataIn1 = 32'd8241
; 
32'd162757: dataIn1 = 32'd8242
; 
32'd162758: dataIn1 = 32'd6415
; 
32'd162759: dataIn1 = 32'd8193
; 
32'd162760: dataIn1 = 32'd8194
; 
32'd162761: dataIn1 = 32'd8197
; 
32'd162762: dataIn1 = 32'd8198
; 
32'd162763: dataIn1 = 32'd8267
; 
32'd162764: dataIn1 = 32'd8268
; 
32'd162765: dataIn1 = 32'd6416
; 
32'd162766: dataIn1 = 32'd8192
; 
32'd162767: dataIn1 = 32'd8193
; 
32'd162768: dataIn1 = 32'd8195
; 
32'd162769: dataIn1 = 32'd8196
; 
32'd162770: dataIn1 = 32'd8222
; 
32'd162771: dataIn1 = 32'd8223
; 
32'd162772: dataIn1 = 32'd6417
; 
32'd162773: dataIn1 = 32'd8200
; 
32'd162774: dataIn1 = 32'd8201
; 
32'd162775: dataIn1 = 32'd8203
; 
32'd162776: dataIn1 = 32'd8205
; 
32'd162777: dataIn1 = 32'd8250
; 
32'd162778: dataIn1 = 32'd8251
; 
32'd162779: dataIn1 = 32'd6418
; 
32'd162780: dataIn1 = 32'd8199
; 
32'd162781: dataIn1 = 32'd8201
; 
32'd162782: dataIn1 = 32'd8202
; 
32'd162783: dataIn1 = 32'd8204
; 
32'd162784: dataIn1 = 32'd8227
; 
32'd162785: dataIn1 = 32'd8229
; 
32'd162786: dataIn1 = 32'd6419
; 
32'd162787: dataIn1 = 32'd8207
; 
32'd162788: dataIn1 = 32'd8208
; 
32'd162789: dataIn1 = 32'd8212
; 
32'd162790: dataIn1 = 32'd8214
; 
32'd162791: dataIn1 = 32'd8216
; 
32'd162792: dataIn1 = 32'd8217
; 
32'd162793: dataIn1 = 32'd6420
; 
32'd162794: dataIn1 = 32'd8206
; 
32'd162795: dataIn1 = 32'd8208
; 
32'd162796: dataIn1 = 32'd8210
; 
32'd162797: dataIn1 = 32'd8213
; 
32'd162798: dataIn1 = 32'd8222
; 
32'd162799: dataIn1 = 32'd8224
; 
32'd162800: dataIn1 = 32'd6421
; 
32'd162801: dataIn1 = 32'd8206
; 
32'd162802: dataIn1 = 32'd8207
; 
32'd162803: dataIn1 = 32'd8209
; 
32'd162804: dataIn1 = 32'd8211
; 
32'd162805: dataIn1 = 32'd8227
; 
32'd162806: dataIn1 = 32'd8228
; 
32'd162807: dataIn1 = 32'd6422
; 
32'd162808: dataIn1 = 32'd8215
; 
32'd162809: dataIn1 = 32'd8217
; 
32'd162810: dataIn1 = 32'd8219
; 
32'd162811: dataIn1 = 32'd8221
; 
32'd162812: dataIn1 = 32'd9111
; 
32'd162813: dataIn1 = 32'd9112
; 
32'd162814: dataIn1 = 32'd6423
; 
32'd162815: dataIn1 = 32'd8223
; 
32'd162816: dataIn1 = 32'd8224
; 
32'd162817: dataIn1 = 32'd8225
; 
32'd162818: dataIn1 = 32'd8226
; 
32'd162819: dataIn1 = 32'd9118
; 
32'd162820: dataIn1 = 32'd9119
; 
32'd162821: dataIn1 = 32'd6424
; 
32'd162822: dataIn1 = 32'd8233
; 
32'd162823: dataIn1 = 32'd8234
; 
32'd162824: dataIn1 = 32'd8238
; 
32'd162825: dataIn1 = 32'd8240
; 
32'd162826: dataIn1 = 32'd8242
; 
32'd162827: dataIn1 = 32'd8243
; 
32'd162828: dataIn1 = 32'd6425
; 
32'd162829: dataIn1 = 32'd8232
; 
32'd162830: dataIn1 = 32'd8234
; 
32'd162831: dataIn1 = 32'd8236
; 
32'd162832: dataIn1 = 32'd8239
; 
32'd162833: dataIn1 = 32'd8244
; 
32'd162834: dataIn1 = 32'd8246
; 
32'd162835: dataIn1 = 32'd6426
; 
32'd162836: dataIn1 = 32'd8232
; 
32'd162837: dataIn1 = 32'd8233
; 
32'd162838: dataIn1 = 32'd8235
; 
32'd162839: dataIn1 = 32'd8237
; 
32'd162840: dataIn1 = 32'd8249
; 
32'd162841: dataIn1 = 32'd8250
; 
32'd162842: dataIn1 = 32'd6427
; 
32'd162843: dataIn1 = 32'd8255
; 
32'd162844: dataIn1 = 32'd8256
; 
32'd162845: dataIn1 = 32'd8260
; 
32'd162846: dataIn1 = 32'd8262
; 
32'd162847: dataIn1 = 32'd8264
; 
32'd162848: dataIn1 = 32'd8265
; 
32'd162849: dataIn1 = 32'd6428
; 
32'd162850: dataIn1 = 32'd8254
; 
32'd162851: dataIn1 = 32'd8256
; 
32'd162852: dataIn1 = 32'd8258
; 
32'd162853: dataIn1 = 32'd8261
; 
32'd162854: dataIn1 = 32'd8266
; 
32'd162855: dataIn1 = 32'd8268
; 
32'd162856: dataIn1 = 32'd6429
; 
32'd162857: dataIn1 = 32'd6764
; 
32'd162858: dataIn1 = 32'd6765
; 
32'd162859: dataIn1 = 32'd8254
; 
32'd162860: dataIn1 = 32'd8255
; 
32'd162861: dataIn1 = 32'd8257
; 
32'd162862: dataIn1 = 32'd8259
; 
32'd162863: dataIn1 = 32'd6430
; 
32'd162864: dataIn1 = 32'd8266
; 
32'd162865: dataIn1 = 32'd8267
; 
32'd162866: dataIn1 = 32'd8269
; 
32'd162867: dataIn1 = 32'd8270
; 
32'd162868: dataIn1 = 32'd9120
; 
32'd162869: dataIn1 = 32'd9122
; 
32'd162870: dataIn1 = 32'd6431
; 
32'd162871: dataIn1 = 32'd8272
; 
32'd162872: dataIn1 = 32'd8273
; 
32'd162873: dataIn1 = 32'd8277
; 
32'd162874: dataIn1 = 32'd8279
; 
32'd162875: dataIn1 = 32'd8281
; 
32'd162876: dataIn1 = 32'd8282
; 
32'd162877: dataIn1 = 32'd6432
; 
32'd162878: dataIn1 = 32'd8271
; 
32'd162879: dataIn1 = 32'd8273
; 
32'd162880: dataIn1 = 32'd8275
; 
32'd162881: dataIn1 = 32'd8278
; 
32'd162882: dataIn1 = 32'd8287
; 
32'd162883: dataIn1 = 32'd8289
; 
32'd162884: dataIn1 = 32'd6433
; 
32'd162885: dataIn1 = 32'd8271
; 
32'd162886: dataIn1 = 32'd8272
; 
32'd162887: dataIn1 = 32'd8274
; 
32'd162888: dataIn1 = 32'd8276
; 
32'd162889: dataIn1 = 32'd8294
; 
32'd162890: dataIn1 = 32'd8295
; 
32'd162891: dataIn1 = 32'd6434
; 
32'd162892: dataIn1 = 32'd8280
; 
32'd162893: dataIn1 = 32'd8282
; 
32'd162894: dataIn1 = 32'd8284
; 
32'd162895: dataIn1 = 32'd8286
; 
32'd162896: dataIn1 = 32'd8348
; 
32'd162897: dataIn1 = 32'd8350
; 
32'd162898: dataIn1 = 32'd6435
; 
32'd162899: dataIn1 = 32'd8280
; 
32'd162900: dataIn1 = 32'd8281
; 
32'd162901: dataIn1 = 32'd8283
; 
32'd162902: dataIn1 = 32'd8285
; 
32'd162903: dataIn1 = 32'd8326
; 
32'd162904: dataIn1 = 32'd8327
; 
32'd162905: dataIn1 = 32'd6436
; 
32'd162906: dataIn1 = 32'd8288
; 
32'd162907: dataIn1 = 32'd8289
; 
32'd162908: dataIn1 = 32'd8292
; 
32'd162909: dataIn1 = 32'd8293
; 
32'd162910: dataIn1 = 32'd8354
; 
32'd162911: dataIn1 = 32'd8355
; 
32'd162912: dataIn1 = 32'd6437
; 
32'd162913: dataIn1 = 32'd8287
; 
32'd162914: dataIn1 = 32'd8288
; 
32'd162915: dataIn1 = 32'd8290
; 
32'd162916: dataIn1 = 32'd8291
; 
32'd162917: dataIn1 = 32'd8310
; 
32'd162918: dataIn1 = 32'd8311
; 
32'd162919: dataIn1 = 32'd6438
; 
32'd162920: dataIn1 = 32'd8295
; 
32'd162921: dataIn1 = 32'd8296
; 
32'd162922: dataIn1 = 32'd8298
; 
32'd162923: dataIn1 = 32'd8300
; 
32'd162924: dataIn1 = 32'd8337
; 
32'd162925: dataIn1 = 32'd8338
; 
32'd162926: dataIn1 = 32'd6439
; 
32'd162927: dataIn1 = 32'd8294
; 
32'd162928: dataIn1 = 32'd8296
; 
32'd162929: dataIn1 = 32'd8297
; 
32'd162930: dataIn1 = 32'd8299
; 
32'd162931: dataIn1 = 32'd8314
; 
32'd162932: dataIn1 = 32'd8316
; 
32'd162933: dataIn1 = 32'd6440
; 
32'd162934: dataIn1 = 32'd6443
; 
32'd162935: dataIn1 = 32'd8302
; 
32'd162936: dataIn1 = 32'd8303
; 
32'd162937: dataIn1 = 32'd8307
; 
32'd162938: dataIn1 = 32'd8309
; 
32'd162939: dataIn1 = 32'd10280
; 
32'd162940: dataIn1 = 32'd6441
; 
32'd162941: dataIn1 = 32'd8301
; 
32'd162942: dataIn1 = 32'd8303
; 
32'd162943: dataIn1 = 32'd8305
; 
32'd162944: dataIn1 = 32'd8308
; 
32'd162945: dataIn1 = 32'd8310
; 
32'd162946: dataIn1 = 32'd8312
; 
32'd162947: dataIn1 = 32'd6442
; 
32'd162948: dataIn1 = 32'd8301
; 
32'd162949: dataIn1 = 32'd8302
; 
32'd162950: dataIn1 = 32'd8304
; 
32'd162951: dataIn1 = 32'd8306
; 
32'd162952: dataIn1 = 32'd8314
; 
32'd162953: dataIn1 = 32'd8315
; 
32'd162954: dataIn1 = 32'd1129
; 
32'd162955: dataIn1 = 32'd5224
; 
32'd162956: dataIn1 = 32'd6396
; 
32'd162957: dataIn1 = 32'd6440
; 
32'd162958: dataIn1 = 32'd6443
; 
32'd162959: dataIn1 = 32'd6676
; 
32'd162960: dataIn1 = 32'd6678
; 
32'd162961: dataIn1 = 32'd8309
; 
32'd162962: dataIn1 = 32'd10280
; 
32'd162963: dataIn1 = 32'd6444
; 
32'd162964: dataIn1 = 32'd8311
; 
32'd162965: dataIn1 = 32'd8312
; 
32'd162966: dataIn1 = 32'd8313
; 
32'd162967: dataIn1 = 32'd9177
; 
32'd162968: dataIn1 = 32'd9178
; 
32'd162969: dataIn1 = 32'd9275
; 
32'd162970: dataIn1 = 32'd6445
; 
32'd162971: dataIn1 = 32'd8318
; 
32'd162972: dataIn1 = 32'd8319
; 
32'd162973: dataIn1 = 32'd8323
; 
32'd162974: dataIn1 = 32'd8325
; 
32'd162975: dataIn1 = 32'd8327
; 
32'd162976: dataIn1 = 32'd8328
; 
32'd162977: dataIn1 = 32'd6446
; 
32'd162978: dataIn1 = 32'd8317
; 
32'd162979: dataIn1 = 32'd8319
; 
32'd162980: dataIn1 = 32'd8321
; 
32'd162981: dataIn1 = 32'd8324
; 
32'd162982: dataIn1 = 32'd8331
; 
32'd162983: dataIn1 = 32'd8333
; 
32'd162984: dataIn1 = 32'd6447
; 
32'd162985: dataIn1 = 32'd8317
; 
32'd162986: dataIn1 = 32'd8318
; 
32'd162987: dataIn1 = 32'd8320
; 
32'd162988: dataIn1 = 32'd8322
; 
32'd162989: dataIn1 = 32'd8336
; 
32'd162990: dataIn1 = 32'd8337
; 
32'd162991: dataIn1 = 32'd6448
; 
32'd162992: dataIn1 = 32'd8340
; 
32'd162993: dataIn1 = 32'd8341
; 
32'd162994: dataIn1 = 32'd8345
; 
32'd162995: dataIn1 = 32'd8347
; 
32'd162996: dataIn1 = 32'd8349
; 
32'd162997: dataIn1 = 32'd8350
; 
32'd162998: dataIn1 = 32'd6449
; 
32'd162999: dataIn1 = 32'd8339
; 
32'd163000: dataIn1 = 32'd8341
; 
32'd163001: dataIn1 = 32'd8343
; 
32'd163002: dataIn1 = 32'd8346
; 
32'd163003: dataIn1 = 32'd8353
; 
32'd163004: dataIn1 = 32'd8355
; 
32'd163005: dataIn1 = 32'd6450
; 
32'd163006: dataIn1 = 32'd8339
; 
32'd163007: dataIn1 = 32'd8340
; 
32'd163008: dataIn1 = 32'd8342
; 
32'd163009: dataIn1 = 32'd8344
; 
32'd163010: dataIn1 = 32'd8358
; 
32'd163011: dataIn1 = 32'd8359
; 
32'd163012: dataIn1 = 32'd6451
; 
32'd163013: dataIn1 = 32'd8353
; 
32'd163014: dataIn1 = 32'd8354
; 
32'd163015: dataIn1 = 32'd8356
; 
32'd163016: dataIn1 = 32'd8357
; 
32'd163017: dataIn1 = 32'd9167
; 
32'd163018: dataIn1 = 32'd9168
; 
32'd163019: dataIn1 = 32'd6452
; 
32'd163020: dataIn1 = 32'd8358
; 
32'd163021: dataIn1 = 32'd8360
; 
32'd163022: dataIn1 = 32'd8361
; 
32'd163023: dataIn1 = 32'd8363
; 
32'd163024: dataIn1 = 32'd9163
; 
32'd163025: dataIn1 = 32'd9165
; 
32'd163026: dataIn1 = 32'd6453
; 
32'd163027: dataIn1 = 32'd8366
; 
32'd163028: dataIn1 = 32'd8367
; 
32'd163029: dataIn1 = 32'd8371
; 
32'd163030: dataIn1 = 32'd8373
; 
32'd163031: dataIn1 = 32'd8375
; 
32'd163032: dataIn1 = 32'd8376
; 
32'd163033: dataIn1 = 32'd6454
; 
32'd163034: dataIn1 = 32'd6766
; 
32'd163035: dataIn1 = 32'd6767
; 
32'd163036: dataIn1 = 32'd8365
; 
32'd163037: dataIn1 = 32'd8367
; 
32'd163038: dataIn1 = 32'd8369
; 
32'd163039: dataIn1 = 32'd8372
; 
32'd163040: dataIn1 = 32'd6455
; 
32'd163041: dataIn1 = 32'd8365
; 
32'd163042: dataIn1 = 32'd8366
; 
32'd163043: dataIn1 = 32'd8368
; 
32'd163044: dataIn1 = 32'd8370
; 
32'd163045: dataIn1 = 32'd8381
; 
32'd163046: dataIn1 = 32'd8382
; 
32'd163047: dataIn1 = 32'd6456
; 
32'd163048: dataIn1 = 32'd8374
; 
32'd163049: dataIn1 = 32'd8376
; 
32'd163050: dataIn1 = 32'd8378
; 
32'd163051: dataIn1 = 32'd8380
; 
32'd163052: dataIn1 = 32'd8421
; 
32'd163053: dataIn1 = 32'd8423
; 
32'd163054: dataIn1 = 32'd6457
; 
32'd163055: dataIn1 = 32'd8374
; 
32'd163056: dataIn1 = 32'd8375
; 
32'd163057: dataIn1 = 32'd8377
; 
32'd163058: dataIn1 = 32'd8379
; 
32'd163059: dataIn1 = 32'd8404
; 
32'd163060: dataIn1 = 32'd8405
; 
32'd163061: dataIn1 = 32'd6458
; 
32'd163062: dataIn1 = 32'd8382
; 
32'd163063: dataIn1 = 32'd8383
; 
32'd163064: dataIn1 = 32'd8385
; 
32'd163065: dataIn1 = 32'd8387
; 
32'd163066: dataIn1 = 32'd8417
; 
32'd163067: dataIn1 = 32'd8418
; 
32'd163068: dataIn1 = 32'd6459
; 
32'd163069: dataIn1 = 32'd8381
; 
32'd163070: dataIn1 = 32'd8383
; 
32'd163071: dataIn1 = 32'd8384
; 
32'd163072: dataIn1 = 32'd8386
; 
32'd163073: dataIn1 = 32'd8388
; 
32'd163074: dataIn1 = 32'd8390
; 
32'd163075: dataIn1 = 32'd6460
; 
32'd163076: dataIn1 = 32'd8389
; 
32'd163077: dataIn1 = 32'd8390
; 
32'd163078: dataIn1 = 32'd8393
; 
32'd163079: dataIn1 = 32'd8394
; 
32'd163080: dataIn1 = 32'd8568
; 
32'd163081: dataIn1 = 32'd8569
; 
32'd163082: dataIn1 = 32'd6461
; 
32'd163083: dataIn1 = 32'd6768
; 
32'd163084: dataIn1 = 32'd6769
; 
32'd163085: dataIn1 = 32'd8388
; 
32'd163086: dataIn1 = 32'd8389
; 
32'd163087: dataIn1 = 32'd8391
; 
32'd163088: dataIn1 = 32'd8392
; 
32'd163089: dataIn1 = 32'd6462
; 
32'd163090: dataIn1 = 32'd8396
; 
32'd163091: dataIn1 = 32'd8397
; 
32'd163092: dataIn1 = 32'd8401
; 
32'd163093: dataIn1 = 32'd8403
; 
32'd163094: dataIn1 = 32'd8405
; 
32'd163095: dataIn1 = 32'd8406
; 
32'd163096: dataIn1 = 32'd6463
; 
32'd163097: dataIn1 = 32'd8395
; 
32'd163098: dataIn1 = 32'd8397
; 
32'd163099: dataIn1 = 32'd8399
; 
32'd163100: dataIn1 = 32'd8402
; 
32'd163101: dataIn1 = 32'd8409
; 
32'd163102: dataIn1 = 32'd8411
; 
32'd163103: dataIn1 = 32'd6464
; 
32'd163104: dataIn1 = 32'd8395
; 
32'd163105: dataIn1 = 32'd8396
; 
32'd163106: dataIn1 = 32'd8398
; 
32'd163107: dataIn1 = 32'd8400
; 
32'd163108: dataIn1 = 32'd8416
; 
32'd163109: dataIn1 = 32'd8417
; 
32'd163110: dataIn1 = 32'd6465
; 
32'd163111: dataIn1 = 32'd8404
; 
32'd163112: dataIn1 = 32'd8406
; 
32'd163113: dataIn1 = 32'd8407
; 
32'd163114: dataIn1 = 32'd8408
; 
32'd163115: dataIn1 = 32'd8493
; 
32'd163116: dataIn1 = 32'd8495
; 
32'd163117: dataIn1 = 32'd6466
; 
32'd163118: dataIn1 = 32'd8410
; 
32'd163119: dataIn1 = 32'd8411
; 
32'd163120: dataIn1 = 32'd8414
; 
32'd163121: dataIn1 = 32'd8415
; 
32'd163122: dataIn1 = 32'd8497
; 
32'd163123: dataIn1 = 32'd8498
; 
32'd163124: dataIn1 = 32'd6467
; 
32'd163125: dataIn1 = 32'd8409
; 
32'd163126: dataIn1 = 32'd8410
; 
32'd163127: dataIn1 = 32'd8412
; 
32'd163128: dataIn1 = 32'd8413
; 
32'd163129: dataIn1 = 32'd8584
; 
32'd163130: dataIn1 = 32'd8585
; 
32'd163131: dataIn1 = 32'd6468
; 
32'd163132: dataIn1 = 32'd8416
; 
32'd163133: dataIn1 = 32'd8418
; 
32'd163134: dataIn1 = 32'd8419
; 
32'd163135: dataIn1 = 32'd8420
; 
32'd163136: dataIn1 = 32'd8589
; 
32'd163137: dataIn1 = 32'd8591
; 
32'd163138: dataIn1 = 32'd6469
; 
32'd163139: dataIn1 = 32'd6770
; 
32'd163140: dataIn1 = 32'd6771
; 
32'd163141: dataIn1 = 32'd8422
; 
32'd163142: dataIn1 = 32'd8423
; 
32'd163143: dataIn1 = 32'd8426
; 
32'd163144: dataIn1 = 32'd8427
; 
32'd163145: dataIn1 = 32'd6470
; 
32'd163146: dataIn1 = 32'd8421
; 
32'd163147: dataIn1 = 32'd8422
; 
32'd163148: dataIn1 = 32'd8424
; 
32'd163149: dataIn1 = 32'd8425
; 
32'd163150: dataIn1 = 32'd8515
; 
32'd163151: dataIn1 = 32'd8516
; 
32'd163152: dataIn1 = 32'd6471
; 
32'd163153: dataIn1 = 32'd8429
; 
32'd163154: dataIn1 = 32'd8430
; 
32'd163155: dataIn1 = 32'd8434
; 
32'd163156: dataIn1 = 32'd8436
; 
32'd163157: dataIn1 = 32'd8438
; 
32'd163158: dataIn1 = 32'd8439
; 
32'd163159: dataIn1 = 32'd6472
; 
32'd163160: dataIn1 = 32'd8428
; 
32'd163161: dataIn1 = 32'd8430
; 
32'd163162: dataIn1 = 32'd8432
; 
32'd163163: dataIn1 = 32'd8435
; 
32'd163164: dataIn1 = 32'd8444
; 
32'd163165: dataIn1 = 32'd8446
; 
32'd163166: dataIn1 = 32'd6473
; 
32'd163167: dataIn1 = 32'd8428
; 
32'd163168: dataIn1 = 32'd8429
; 
32'd163169: dataIn1 = 32'd8431
; 
32'd163170: dataIn1 = 32'd8433
; 
32'd163171: dataIn1 = 32'd8451
; 
32'd163172: dataIn1 = 32'd8452
; 
32'd163173: dataIn1 = 32'd6474
; 
32'd163174: dataIn1 = 32'd8437
; 
32'd163175: dataIn1 = 32'd8439
; 
32'd163176: dataIn1 = 32'd8441
; 
32'd163177: dataIn1 = 32'd8443
; 
32'd163178: dataIn1 = 32'd8515
; 
32'd163179: dataIn1 = 32'd8517
; 
32'd163180: dataIn1 = 32'd6475
; 
32'd163181: dataIn1 = 32'd8437
; 
32'd163182: dataIn1 = 32'd8438
; 
32'd163183: dataIn1 = 32'd8440
; 
32'd163184: dataIn1 = 32'd8442
; 
32'd163185: dataIn1 = 32'd8493
; 
32'd163186: dataIn1 = 32'd8494
; 
32'd163187: dataIn1 = 32'd6476
; 
32'd163188: dataIn1 = 32'd8445
; 
32'd163189: dataIn1 = 32'd8446
; 
32'd163190: dataIn1 = 32'd8449
; 
32'd163191: dataIn1 = 32'd8450
; 
32'd163192: dataIn1 = 32'd8519
; 
32'd163193: dataIn1 = 32'd8520
; 
32'd163194: dataIn1 = 32'd6477
; 
32'd163195: dataIn1 = 32'd8444
; 
32'd163196: dataIn1 = 32'd8445
; 
32'd163197: dataIn1 = 32'd8447
; 
32'd163198: dataIn1 = 32'd8448
; 
32'd163199: dataIn1 = 32'd8474
; 
32'd163200: dataIn1 = 32'd8475
; 
32'd163201: dataIn1 = 32'd6478
; 
32'd163202: dataIn1 = 32'd8452
; 
32'd163203: dataIn1 = 32'd8453
; 
32'd163204: dataIn1 = 32'd8455
; 
32'd163205: dataIn1 = 32'd8457
; 
32'd163206: dataIn1 = 32'd8502
; 
32'd163207: dataIn1 = 32'd8503
; 
32'd163208: dataIn1 = 32'd6479
; 
32'd163209: dataIn1 = 32'd8451
; 
32'd163210: dataIn1 = 32'd8453
; 
32'd163211: dataIn1 = 32'd8454
; 
32'd163212: dataIn1 = 32'd8456
; 
32'd163213: dataIn1 = 32'd8479
; 
32'd163214: dataIn1 = 32'd8481
; 
32'd163215: dataIn1 = 32'd6480
; 
32'd163216: dataIn1 = 32'd8459
; 
32'd163217: dataIn1 = 32'd8460
; 
32'd163218: dataIn1 = 32'd8464
; 
32'd163219: dataIn1 = 32'd8466
; 
32'd163220: dataIn1 = 32'd8468
; 
32'd163221: dataIn1 = 32'd8469
; 
32'd163222: dataIn1 = 32'd6481
; 
32'd163223: dataIn1 = 32'd8458
; 
32'd163224: dataIn1 = 32'd8460
; 
32'd163225: dataIn1 = 32'd8462
; 
32'd163226: dataIn1 = 32'd8465
; 
32'd163227: dataIn1 = 32'd8474
; 
32'd163228: dataIn1 = 32'd8476
; 
32'd163229: dataIn1 = 32'd6482
; 
32'd163230: dataIn1 = 32'd8458
; 
32'd163231: dataIn1 = 32'd8459
; 
32'd163232: dataIn1 = 32'd8461
; 
32'd163233: dataIn1 = 32'd8463
; 
32'd163234: dataIn1 = 32'd8479
; 
32'd163235: dataIn1 = 32'd8480
; 
32'd163236: dataIn1 = 32'd6483
; 
32'd163237: dataIn1 = 32'd8467
; 
32'd163238: dataIn1 = 32'd8469
; 
32'd163239: dataIn1 = 32'd8471
; 
32'd163240: dataIn1 = 32'd8473
; 
32'd163241: dataIn1 = 32'd9163
; 
32'd163242: dataIn1 = 32'd9164
; 
32'd163243: dataIn1 = 32'd6484
; 
32'd163244: dataIn1 = 32'd8475
; 
32'd163245: dataIn1 = 32'd8476
; 
32'd163246: dataIn1 = 32'd8477
; 
32'd163247: dataIn1 = 32'd8478
; 
32'd163248: dataIn1 = 32'd9170
; 
32'd163249: dataIn1 = 32'd9171
; 
32'd163250: dataIn1 = 32'd6485
; 
32'd163251: dataIn1 = 32'd8485
; 
32'd163252: dataIn1 = 32'd8486
; 
32'd163253: dataIn1 = 32'd8490
; 
32'd163254: dataIn1 = 32'd8492
; 
32'd163255: dataIn1 = 32'd8494
; 
32'd163256: dataIn1 = 32'd8495
; 
32'd163257: dataIn1 = 32'd6486
; 
32'd163258: dataIn1 = 32'd8484
; 
32'd163259: dataIn1 = 32'd8486
; 
32'd163260: dataIn1 = 32'd8488
; 
32'd163261: dataIn1 = 32'd8491
; 
32'd163262: dataIn1 = 32'd8496
; 
32'd163263: dataIn1 = 32'd8498
; 
32'd163264: dataIn1 = 32'd6487
; 
32'd163265: dataIn1 = 32'd8484
; 
32'd163266: dataIn1 = 32'd8485
; 
32'd163267: dataIn1 = 32'd8487
; 
32'd163268: dataIn1 = 32'd8489
; 
32'd163269: dataIn1 = 32'd8501
; 
32'd163270: dataIn1 = 32'd8502
; 
32'd163271: dataIn1 = 32'd6488
; 
32'd163272: dataIn1 = 32'd8507
; 
32'd163273: dataIn1 = 32'd8508
; 
32'd163274: dataIn1 = 32'd8512
; 
32'd163275: dataIn1 = 32'd8514
; 
32'd163276: dataIn1 = 32'd8516
; 
32'd163277: dataIn1 = 32'd8517
; 
32'd163278: dataIn1 = 32'd6489
; 
32'd163279: dataIn1 = 32'd8506
; 
32'd163280: dataIn1 = 32'd8508
; 
32'd163281: dataIn1 = 32'd8510
; 
32'd163282: dataIn1 = 32'd8513
; 
32'd163283: dataIn1 = 32'd8518
; 
32'd163284: dataIn1 = 32'd8520
; 
32'd163285: dataIn1 = 32'd6490
; 
32'd163286: dataIn1 = 32'd6772
; 
32'd163287: dataIn1 = 32'd6773
; 
32'd163288: dataIn1 = 32'd8506
; 
32'd163289: dataIn1 = 32'd8507
; 
32'd163290: dataIn1 = 32'd8509
; 
32'd163291: dataIn1 = 32'd8511
; 
32'd163292: dataIn1 = 32'd6491
; 
32'd163293: dataIn1 = 32'd8518
; 
32'd163294: dataIn1 = 32'd8519
; 
32'd163295: dataIn1 = 32'd8521
; 
32'd163296: dataIn1 = 32'd8522
; 
32'd163297: dataIn1 = 32'd9172
; 
32'd163298: dataIn1 = 32'd9174
; 
32'd163299: dataIn1 = 32'd6492
; 
32'd163300: dataIn1 = 32'd8524
; 
32'd163301: dataIn1 = 32'd8525
; 
32'd163302: dataIn1 = 32'd8529
; 
32'd163303: dataIn1 = 32'd8531
; 
32'd163304: dataIn1 = 32'd8533
; 
32'd163305: dataIn1 = 32'd8534
; 
32'd163306: dataIn1 = 32'd6493
; 
32'd163307: dataIn1 = 32'd8523
; 
32'd163308: dataIn1 = 32'd8525
; 
32'd163309: dataIn1 = 32'd8527
; 
32'd163310: dataIn1 = 32'd8530
; 
32'd163311: dataIn1 = 32'd8539
; 
32'd163312: dataIn1 = 32'd8541
; 
32'd163313: dataIn1 = 32'd6494
; 
32'd163314: dataIn1 = 32'd8523
; 
32'd163315: dataIn1 = 32'd8524
; 
32'd163316: dataIn1 = 32'd8526
; 
32'd163317: dataIn1 = 32'd8528
; 
32'd163318: dataIn1 = 32'd8546
; 
32'd163319: dataIn1 = 32'd8547
; 
32'd163320: dataIn1 = 32'd6495
; 
32'd163321: dataIn1 = 32'd8532
; 
32'd163322: dataIn1 = 32'd8534
; 
32'd163323: dataIn1 = 32'd8536
; 
32'd163324: dataIn1 = 32'd8538
; 
32'd163325: dataIn1 = 32'd8601
; 
32'd163326: dataIn1 = 32'd8603
; 
32'd163327: dataIn1 = 32'd6496
; 
32'd163328: dataIn1 = 32'd8532
; 
32'd163329: dataIn1 = 32'd8533
; 
32'd163330: dataIn1 = 32'd8535
; 
32'd163331: dataIn1 = 32'd8537
; 
32'd163332: dataIn1 = 32'd8579
; 
32'd163333: dataIn1 = 32'd8580
; 
32'd163334: dataIn1 = 32'd6497
; 
32'd163335: dataIn1 = 32'd8540
; 
32'd163336: dataIn1 = 32'd8541
; 
32'd163337: dataIn1 = 32'd8544
; 
32'd163338: dataIn1 = 32'd8545
; 
32'd163339: dataIn1 = 32'd8607
; 
32'd163340: dataIn1 = 32'd8608
; 
32'd163341: dataIn1 = 32'd6498
; 
32'd163342: dataIn1 = 32'd8539
; 
32'd163343: dataIn1 = 32'd8540
; 
32'd163344: dataIn1 = 32'd8542
; 
32'd163345: dataIn1 = 32'd8543
; 
32'd163346: dataIn1 = 32'd8562
; 
32'd163347: dataIn1 = 32'd8563
; 
32'd163348: dataIn1 = 32'd6499
; 
32'd163349: dataIn1 = 32'd8547
; 
32'd163350: dataIn1 = 32'd8548
; 
32'd163351: dataIn1 = 32'd8550
; 
32'd163352: dataIn1 = 32'd8552
; 
32'd163353: dataIn1 = 32'd8590
; 
32'd163354: dataIn1 = 32'd8591
; 
32'd163355: dataIn1 = 32'd6500
; 
32'd163356: dataIn1 = 32'd8546
; 
32'd163357: dataIn1 = 32'd8548
; 
32'd163358: dataIn1 = 32'd8549
; 
32'd163359: dataIn1 = 32'd8551
; 
32'd163360: dataIn1 = 32'd8567
; 
32'd163361: dataIn1 = 32'd8569
; 
32'd163362: dataIn1 = 32'd6501
; 
32'd163363: dataIn1 = 32'd6774
; 
32'd163364: dataIn1 = 32'd6775
; 
32'd163365: dataIn1 = 32'd8554
; 
32'd163366: dataIn1 = 32'd8555
; 
32'd163367: dataIn1 = 32'd8559
; 
32'd163368: dataIn1 = 32'd8561
; 
32'd163369: dataIn1 = 32'd6502
; 
32'd163370: dataIn1 = 32'd8553
; 
32'd163371: dataIn1 = 32'd8555
; 
32'd163372: dataIn1 = 32'd8557
; 
32'd163373: dataIn1 = 32'd8560
; 
32'd163374: dataIn1 = 32'd8562
; 
32'd163375: dataIn1 = 32'd8564
; 
32'd163376: dataIn1 = 32'd6503
; 
32'd163377: dataIn1 = 32'd8553
; 
32'd163378: dataIn1 = 32'd8554
; 
32'd163379: dataIn1 = 32'd8556
; 
32'd163380: dataIn1 = 32'd8558
; 
32'd163381: dataIn1 = 32'd8567
; 
32'd163382: dataIn1 = 32'd8568
; 
32'd163383: dataIn1 = 32'd6504
; 
32'd163384: dataIn1 = 32'd8563
; 
32'd163385: dataIn1 = 32'd8564
; 
32'd163386: dataIn1 = 32'd8565
; 
32'd163387: dataIn1 = 32'd8566
; 
32'd163388: dataIn1 = 32'd9227
; 
32'd163389: dataIn1 = 32'd9228
; 
32'd163390: dataIn1 = 32'd6505
; 
32'd163391: dataIn1 = 32'd8571
; 
32'd163392: dataIn1 = 32'd8572
; 
32'd163393: dataIn1 = 32'd8576
; 
32'd163394: dataIn1 = 32'd8578
; 
32'd163395: dataIn1 = 32'd8580
; 
32'd163396: dataIn1 = 32'd8581
; 
32'd163397: dataIn1 = 32'd6506
; 
32'd163398: dataIn1 = 32'd8570
; 
32'd163399: dataIn1 = 32'd8572
; 
32'd163400: dataIn1 = 32'd8574
; 
32'd163401: dataIn1 = 32'd8577
; 
32'd163402: dataIn1 = 32'd8584
; 
32'd163403: dataIn1 = 32'd8586
; 
32'd163404: dataIn1 = 32'd6507
; 
32'd163405: dataIn1 = 32'd8570
; 
32'd163406: dataIn1 = 32'd8571
; 
32'd163407: dataIn1 = 32'd8573
; 
32'd163408: dataIn1 = 32'd8575
; 
32'd163409: dataIn1 = 32'd8589
; 
32'd163410: dataIn1 = 32'd8590
; 
32'd163411: dataIn1 = 32'd6508
; 
32'd163412: dataIn1 = 32'd8593
; 
32'd163413: dataIn1 = 32'd8594
; 
32'd163414: dataIn1 = 32'd8598
; 
32'd163415: dataIn1 = 32'd8600
; 
32'd163416: dataIn1 = 32'd8602
; 
32'd163417: dataIn1 = 32'd8603
; 
32'd163418: dataIn1 = 32'd6509
; 
32'd163419: dataIn1 = 32'd8592
; 
32'd163420: dataIn1 = 32'd8594
; 
32'd163421: dataIn1 = 32'd8596
; 
32'd163422: dataIn1 = 32'd8599
; 
32'd163423: dataIn1 = 32'd8606
; 
32'd163424: dataIn1 = 32'd8608
; 
32'd163425: dataIn1 = 32'd6510
; 
32'd163426: dataIn1 = 32'd8592
; 
32'd163427: dataIn1 = 32'd8593
; 
32'd163428: dataIn1 = 32'd8595
; 
32'd163429: dataIn1 = 32'd8597
; 
32'd163430: dataIn1 = 32'd8611
; 
32'd163431: dataIn1 = 32'd8612
; 
32'd163432: dataIn1 = 32'd6511
; 
32'd163433: dataIn1 = 32'd8606
; 
32'd163434: dataIn1 = 32'd8607
; 
32'd163435: dataIn1 = 32'd8609
; 
32'd163436: dataIn1 = 32'd8610
; 
32'd163437: dataIn1 = 32'd9217
; 
32'd163438: dataIn1 = 32'd9218
; 
32'd163439: dataIn1 = 32'd6512
; 
32'd163440: dataIn1 = 32'd8611
; 
32'd163441: dataIn1 = 32'd8613
; 
32'd163442: dataIn1 = 32'd8614
; 
32'd163443: dataIn1 = 32'd8616
; 
32'd163444: dataIn1 = 32'd9213
; 
32'd163445: dataIn1 = 32'd9215
; 
32'd163446: dataIn1 = 32'd6513
; 
32'd163447: dataIn1 = 32'd8619
; 
32'd163448: dataIn1 = 32'd8620
; 
32'd163449: dataIn1 = 32'd8624
; 
32'd163450: dataIn1 = 32'd8626
; 
32'd163451: dataIn1 = 32'd8628
; 
32'd163452: dataIn1 = 32'd8629
; 
32'd163453: dataIn1 = 32'd6514
; 
32'd163454: dataIn1 = 32'd6776
; 
32'd163455: dataIn1 = 32'd6777
; 
32'd163456: dataIn1 = 32'd8618
; 
32'd163457: dataIn1 = 32'd8620
; 
32'd163458: dataIn1 = 32'd8622
; 
32'd163459: dataIn1 = 32'd8625
; 
32'd163460: dataIn1 = 32'd6515
; 
32'd163461: dataIn1 = 32'd8618
; 
32'd163462: dataIn1 = 32'd8619
; 
32'd163463: dataIn1 = 32'd8621
; 
32'd163464: dataIn1 = 32'd8623
; 
32'd163465: dataIn1 = 32'd8634
; 
32'd163466: dataIn1 = 32'd8635
; 
32'd163467: dataIn1 = 32'd6516
; 
32'd163468: dataIn1 = 32'd8627
; 
32'd163469: dataIn1 = 32'd8629
; 
32'd163470: dataIn1 = 32'd8631
; 
32'd163471: dataIn1 = 32'd8633
; 
32'd163472: dataIn1 = 32'd8674
; 
32'd163473: dataIn1 = 32'd8676
; 
32'd163474: dataIn1 = 32'd6517
; 
32'd163475: dataIn1 = 32'd8627
; 
32'd163476: dataIn1 = 32'd8628
; 
32'd163477: dataIn1 = 32'd8630
; 
32'd163478: dataIn1 = 32'd8632
; 
32'd163479: dataIn1 = 32'd8657
; 
32'd163480: dataIn1 = 32'd8658
; 
32'd163481: dataIn1 = 32'd6518
; 
32'd163482: dataIn1 = 32'd8635
; 
32'd163483: dataIn1 = 32'd8636
; 
32'd163484: dataIn1 = 32'd8638
; 
32'd163485: dataIn1 = 32'd8640
; 
32'd163486: dataIn1 = 32'd8670
; 
32'd163487: dataIn1 = 32'd8671
; 
32'd163488: dataIn1 = 32'd6519
; 
32'd163489: dataIn1 = 32'd8634
; 
32'd163490: dataIn1 = 32'd8636
; 
32'd163491: dataIn1 = 32'd8637
; 
32'd163492: dataIn1 = 32'd8639
; 
32'd163493: dataIn1 = 32'd8641
; 
32'd163494: dataIn1 = 32'd8643
; 
32'd163495: dataIn1 = 32'd6520
; 
32'd163496: dataIn1 = 32'd8642
; 
32'd163497: dataIn1 = 32'd8643
; 
32'd163498: dataIn1 = 32'd8646
; 
32'd163499: dataIn1 = 32'd8647
; 
32'd163500: dataIn1 = 32'd8820
; 
32'd163501: dataIn1 = 32'd8821
; 
32'd163502: dataIn1 = 32'd6521
; 
32'd163503: dataIn1 = 32'd6778
; 
32'd163504: dataIn1 = 32'd6779
; 
32'd163505: dataIn1 = 32'd8641
; 
32'd163506: dataIn1 = 32'd8642
; 
32'd163507: dataIn1 = 32'd8644
; 
32'd163508: dataIn1 = 32'd8645
; 
32'd163509: dataIn1 = 32'd6522
; 
32'd163510: dataIn1 = 32'd8649
; 
32'd163511: dataIn1 = 32'd8650
; 
32'd163512: dataIn1 = 32'd8654
; 
32'd163513: dataIn1 = 32'd8656
; 
32'd163514: dataIn1 = 32'd8658
; 
32'd163515: dataIn1 = 32'd8659
; 
32'd163516: dataIn1 = 32'd6523
; 
32'd163517: dataIn1 = 32'd8648
; 
32'd163518: dataIn1 = 32'd8650
; 
32'd163519: dataIn1 = 32'd8652
; 
32'd163520: dataIn1 = 32'd8655
; 
32'd163521: dataIn1 = 32'd8662
; 
32'd163522: dataIn1 = 32'd8664
; 
32'd163523: dataIn1 = 32'd6524
; 
32'd163524: dataIn1 = 32'd8648
; 
32'd163525: dataIn1 = 32'd8649
; 
32'd163526: dataIn1 = 32'd8651
; 
32'd163527: dataIn1 = 32'd8653
; 
32'd163528: dataIn1 = 32'd8669
; 
32'd163529: dataIn1 = 32'd8670
; 
32'd163530: dataIn1 = 32'd6525
; 
32'd163531: dataIn1 = 32'd8657
; 
32'd163532: dataIn1 = 32'd8659
; 
32'd163533: dataIn1 = 32'd8660
; 
32'd163534: dataIn1 = 32'd8661
; 
32'd163535: dataIn1 = 32'd8746
; 
32'd163536: dataIn1 = 32'd8748
; 
32'd163537: dataIn1 = 32'd6526
; 
32'd163538: dataIn1 = 32'd8663
; 
32'd163539: dataIn1 = 32'd8664
; 
32'd163540: dataIn1 = 32'd8667
; 
32'd163541: dataIn1 = 32'd8668
; 
32'd163542: dataIn1 = 32'd8750
; 
32'd163543: dataIn1 = 32'd8751
; 
32'd163544: dataIn1 = 32'd6527
; 
32'd163545: dataIn1 = 32'd8662
; 
32'd163546: dataIn1 = 32'd8663
; 
32'd163547: dataIn1 = 32'd8665
; 
32'd163548: dataIn1 = 32'd8666
; 
32'd163549: dataIn1 = 32'd8836
; 
32'd163550: dataIn1 = 32'd8837
; 
32'd163551: dataIn1 = 32'd6528
; 
32'd163552: dataIn1 = 32'd8669
; 
32'd163553: dataIn1 = 32'd8671
; 
32'd163554: dataIn1 = 32'd8672
; 
32'd163555: dataIn1 = 32'd8673
; 
32'd163556: dataIn1 = 32'd8841
; 
32'd163557: dataIn1 = 32'd8843
; 
32'd163558: dataIn1 = 32'd6529
; 
32'd163559: dataIn1 = 32'd6780
; 
32'd163560: dataIn1 = 32'd6781
; 
32'd163561: dataIn1 = 32'd8675
; 
32'd163562: dataIn1 = 32'd8676
; 
32'd163563: dataIn1 = 32'd8679
; 
32'd163564: dataIn1 = 32'd8680
; 
32'd163565: dataIn1 = 32'd6530
; 
32'd163566: dataIn1 = 32'd8674
; 
32'd163567: dataIn1 = 32'd8675
; 
32'd163568: dataIn1 = 32'd8677
; 
32'd163569: dataIn1 = 32'd8678
; 
32'd163570: dataIn1 = 32'd8768
; 
32'd163571: dataIn1 = 32'd8769
; 
32'd163572: dataIn1 = 32'd6531
; 
32'd163573: dataIn1 = 32'd8682
; 
32'd163574: dataIn1 = 32'd8683
; 
32'd163575: dataIn1 = 32'd8687
; 
32'd163576: dataIn1 = 32'd8689
; 
32'd163577: dataIn1 = 32'd8691
; 
32'd163578: dataIn1 = 32'd8692
; 
32'd163579: dataIn1 = 32'd6532
; 
32'd163580: dataIn1 = 32'd8681
; 
32'd163581: dataIn1 = 32'd8683
; 
32'd163582: dataIn1 = 32'd8685
; 
32'd163583: dataIn1 = 32'd8688
; 
32'd163584: dataIn1 = 32'd8697
; 
32'd163585: dataIn1 = 32'd8699
; 
32'd163586: dataIn1 = 32'd6533
; 
32'd163587: dataIn1 = 32'd8681
; 
32'd163588: dataIn1 = 32'd8682
; 
32'd163589: dataIn1 = 32'd8684
; 
32'd163590: dataIn1 = 32'd8686
; 
32'd163591: dataIn1 = 32'd8704
; 
32'd163592: dataIn1 = 32'd8705
; 
32'd163593: dataIn1 = 32'd6534
; 
32'd163594: dataIn1 = 32'd8690
; 
32'd163595: dataIn1 = 32'd8692
; 
32'd163596: dataIn1 = 32'd8694
; 
32'd163597: dataIn1 = 32'd8696
; 
32'd163598: dataIn1 = 32'd8768
; 
32'd163599: dataIn1 = 32'd8770
; 
32'd163600: dataIn1 = 32'd6535
; 
32'd163601: dataIn1 = 32'd8690
; 
32'd163602: dataIn1 = 32'd8691
; 
32'd163603: dataIn1 = 32'd8693
; 
32'd163604: dataIn1 = 32'd8695
; 
32'd163605: dataIn1 = 32'd8746
; 
32'd163606: dataIn1 = 32'd8747
; 
32'd163607: dataIn1 = 32'd6536
; 
32'd163608: dataIn1 = 32'd8698
; 
32'd163609: dataIn1 = 32'd8699
; 
32'd163610: dataIn1 = 32'd8702
; 
32'd163611: dataIn1 = 32'd8703
; 
32'd163612: dataIn1 = 32'd8772
; 
32'd163613: dataIn1 = 32'd8773
; 
32'd163614: dataIn1 = 32'd6537
; 
32'd163615: dataIn1 = 32'd8697
; 
32'd163616: dataIn1 = 32'd8698
; 
32'd163617: dataIn1 = 32'd8700
; 
32'd163618: dataIn1 = 32'd8701
; 
32'd163619: dataIn1 = 32'd8727
; 
32'd163620: dataIn1 = 32'd8728
; 
32'd163621: dataIn1 = 32'd6538
; 
32'd163622: dataIn1 = 32'd8705
; 
32'd163623: dataIn1 = 32'd8706
; 
32'd163624: dataIn1 = 32'd8708
; 
32'd163625: dataIn1 = 32'd8710
; 
32'd163626: dataIn1 = 32'd8755
; 
32'd163627: dataIn1 = 32'd8756
; 
32'd163628: dataIn1 = 32'd6539
; 
32'd163629: dataIn1 = 32'd8704
; 
32'd163630: dataIn1 = 32'd8706
; 
32'd163631: dataIn1 = 32'd8707
; 
32'd163632: dataIn1 = 32'd8709
; 
32'd163633: dataIn1 = 32'd8732
; 
32'd163634: dataIn1 = 32'd8734
; 
32'd163635: dataIn1 = 32'd6540
; 
32'd163636: dataIn1 = 32'd8712
; 
32'd163637: dataIn1 = 32'd8713
; 
32'd163638: dataIn1 = 32'd8717
; 
32'd163639: dataIn1 = 32'd8719
; 
32'd163640: dataIn1 = 32'd8721
; 
32'd163641: dataIn1 = 32'd8722
; 
32'd163642: dataIn1 = 32'd6541
; 
32'd163643: dataIn1 = 32'd8711
; 
32'd163644: dataIn1 = 32'd8713
; 
32'd163645: dataIn1 = 32'd8715
; 
32'd163646: dataIn1 = 32'd8718
; 
32'd163647: dataIn1 = 32'd8727
; 
32'd163648: dataIn1 = 32'd8729
; 
32'd163649: dataIn1 = 32'd6542
; 
32'd163650: dataIn1 = 32'd8711
; 
32'd163651: dataIn1 = 32'd8712
; 
32'd163652: dataIn1 = 32'd8714
; 
32'd163653: dataIn1 = 32'd8716
; 
32'd163654: dataIn1 = 32'd8732
; 
32'd163655: dataIn1 = 32'd8733
; 
32'd163656: dataIn1 = 32'd6543
; 
32'd163657: dataIn1 = 32'd8720
; 
32'd163658: dataIn1 = 32'd8722
; 
32'd163659: dataIn1 = 32'd8724
; 
32'd163660: dataIn1 = 32'd8726
; 
32'd163661: dataIn1 = 32'd9213
; 
32'd163662: dataIn1 = 32'd9214
; 
32'd163663: dataIn1 = 32'd6544
; 
32'd163664: dataIn1 = 32'd8728
; 
32'd163665: dataIn1 = 32'd8729
; 
32'd163666: dataIn1 = 32'd8730
; 
32'd163667: dataIn1 = 32'd8731
; 
32'd163668: dataIn1 = 32'd9220
; 
32'd163669: dataIn1 = 32'd9221
; 
32'd163670: dataIn1 = 32'd6545
; 
32'd163671: dataIn1 = 32'd8738
; 
32'd163672: dataIn1 = 32'd8739
; 
32'd163673: dataIn1 = 32'd8743
; 
32'd163674: dataIn1 = 32'd8745
; 
32'd163675: dataIn1 = 32'd8747
; 
32'd163676: dataIn1 = 32'd8748
; 
32'd163677: dataIn1 = 32'd6546
; 
32'd163678: dataIn1 = 32'd8737
; 
32'd163679: dataIn1 = 32'd8739
; 
32'd163680: dataIn1 = 32'd8741
; 
32'd163681: dataIn1 = 32'd8744
; 
32'd163682: dataIn1 = 32'd8749
; 
32'd163683: dataIn1 = 32'd8751
; 
32'd163684: dataIn1 = 32'd6547
; 
32'd163685: dataIn1 = 32'd8737
; 
32'd163686: dataIn1 = 32'd8738
; 
32'd163687: dataIn1 = 32'd8740
; 
32'd163688: dataIn1 = 32'd8742
; 
32'd163689: dataIn1 = 32'd8754
; 
32'd163690: dataIn1 = 32'd8755
; 
32'd163691: dataIn1 = 32'd6548
; 
32'd163692: dataIn1 = 32'd8760
; 
32'd163693: dataIn1 = 32'd8761
; 
32'd163694: dataIn1 = 32'd8765
; 
32'd163695: dataIn1 = 32'd8767
; 
32'd163696: dataIn1 = 32'd8769
; 
32'd163697: dataIn1 = 32'd8770
; 
32'd163698: dataIn1 = 32'd6549
; 
32'd163699: dataIn1 = 32'd8759
; 
32'd163700: dataIn1 = 32'd8761
; 
32'd163701: dataIn1 = 32'd8763
; 
32'd163702: dataIn1 = 32'd8766
; 
32'd163703: dataIn1 = 32'd8771
; 
32'd163704: dataIn1 = 32'd8773
; 
32'd163705: dataIn1 = 32'd6550
; 
32'd163706: dataIn1 = 32'd6782
; 
32'd163707: dataIn1 = 32'd6783
; 
32'd163708: dataIn1 = 32'd8759
; 
32'd163709: dataIn1 = 32'd8760
; 
32'd163710: dataIn1 = 32'd8762
; 
32'd163711: dataIn1 = 32'd8764
; 
32'd163712: dataIn1 = 32'd6551
; 
32'd163713: dataIn1 = 32'd8771
; 
32'd163714: dataIn1 = 32'd8772
; 
32'd163715: dataIn1 = 32'd8774
; 
32'd163716: dataIn1 = 32'd8775
; 
32'd163717: dataIn1 = 32'd9222
; 
32'd163718: dataIn1 = 32'd9224
; 
32'd163719: dataIn1 = 32'd6552
; 
32'd163720: dataIn1 = 32'd8777
; 
32'd163721: dataIn1 = 32'd8778
; 
32'd163722: dataIn1 = 32'd8782
; 
32'd163723: dataIn1 = 32'd8784
; 
32'd163724: dataIn1 = 32'd8786
; 
32'd163725: dataIn1 = 32'd8787
; 
32'd163726: dataIn1 = 32'd6553
; 
32'd163727: dataIn1 = 32'd8776
; 
32'd163728: dataIn1 = 32'd8778
; 
32'd163729: dataIn1 = 32'd8780
; 
32'd163730: dataIn1 = 32'd8783
; 
32'd163731: dataIn1 = 32'd8792
; 
32'd163732: dataIn1 = 32'd8794
; 
32'd163733: dataIn1 = 32'd6554
; 
32'd163734: dataIn1 = 32'd8776
; 
32'd163735: dataIn1 = 32'd8777
; 
32'd163736: dataIn1 = 32'd8779
; 
32'd163737: dataIn1 = 32'd8781
; 
32'd163738: dataIn1 = 32'd8799
; 
32'd163739: dataIn1 = 32'd8800
; 
32'd163740: dataIn1 = 32'd6555
; 
32'd163741: dataIn1 = 32'd8785
; 
32'd163742: dataIn1 = 32'd8787
; 
32'd163743: dataIn1 = 32'd8789
; 
32'd163744: dataIn1 = 32'd8791
; 
32'd163745: dataIn1 = 32'd8853
; 
32'd163746: dataIn1 = 32'd8855
; 
32'd163747: dataIn1 = 32'd6556
; 
32'd163748: dataIn1 = 32'd8785
; 
32'd163749: dataIn1 = 32'd8786
; 
32'd163750: dataIn1 = 32'd8788
; 
32'd163751: dataIn1 = 32'd8790
; 
32'd163752: dataIn1 = 32'd8831
; 
32'd163753: dataIn1 = 32'd8832
; 
32'd163754: dataIn1 = 32'd6557
; 
32'd163755: dataIn1 = 32'd8793
; 
32'd163756: dataIn1 = 32'd8794
; 
32'd163757: dataIn1 = 32'd8797
; 
32'd163758: dataIn1 = 32'd8798
; 
32'd163759: dataIn1 = 32'd8859
; 
32'd163760: dataIn1 = 32'd8860
; 
32'd163761: dataIn1 = 32'd6558
; 
32'd163762: dataIn1 = 32'd8792
; 
32'd163763: dataIn1 = 32'd8793
; 
32'd163764: dataIn1 = 32'd8795
; 
32'd163765: dataIn1 = 32'd8796
; 
32'd163766: dataIn1 = 32'd8815
; 
32'd163767: dataIn1 = 32'd8816
; 
32'd163768: dataIn1 = 32'd6559
; 
32'd163769: dataIn1 = 32'd8800
; 
32'd163770: dataIn1 = 32'd8801
; 
32'd163771: dataIn1 = 32'd8803
; 
32'd163772: dataIn1 = 32'd8805
; 
32'd163773: dataIn1 = 32'd8842
; 
32'd163774: dataIn1 = 32'd8843
; 
32'd163775: dataIn1 = 32'd6560
; 
32'd163776: dataIn1 = 32'd8799
; 
32'd163777: dataIn1 = 32'd8801
; 
32'd163778: dataIn1 = 32'd8802
; 
32'd163779: dataIn1 = 32'd8804
; 
32'd163780: dataIn1 = 32'd8819
; 
32'd163781: dataIn1 = 32'd8821
; 
32'd163782: dataIn1 = 32'd6561
; 
32'd163783: dataIn1 = 32'd6784
; 
32'd163784: dataIn1 = 32'd6785
; 
32'd163785: dataIn1 = 32'd8807
; 
32'd163786: dataIn1 = 32'd8808
; 
32'd163787: dataIn1 = 32'd8812
; 
32'd163788: dataIn1 = 32'd8814
; 
32'd163789: dataIn1 = 32'd6562
; 
32'd163790: dataIn1 = 32'd8806
; 
32'd163791: dataIn1 = 32'd8808
; 
32'd163792: dataIn1 = 32'd8810
; 
32'd163793: dataIn1 = 32'd8813
; 
32'd163794: dataIn1 = 32'd8815
; 
32'd163795: dataIn1 = 32'd8817
; 
32'd163796: dataIn1 = 32'd6563
; 
32'd163797: dataIn1 = 32'd8806
; 
32'd163798: dataIn1 = 32'd8807
; 
32'd163799: dataIn1 = 32'd8809
; 
32'd163800: dataIn1 = 32'd8811
; 
32'd163801: dataIn1 = 32'd8819
; 
32'd163802: dataIn1 = 32'd8820
; 
32'd163803: dataIn1 = 32'd6564
; 
32'd163804: dataIn1 = 32'd8816
; 
32'd163805: dataIn1 = 32'd8817
; 
32'd163806: dataIn1 = 32'd8818
; 
32'd163807: dataIn1 = 32'd9276
; 
32'd163808: dataIn1 = 32'd9442
; 
32'd163809: dataIn1 = 32'd9443
; 
32'd163810: dataIn1 = 32'd6565
; 
32'd163811: dataIn1 = 32'd8823
; 
32'd163812: dataIn1 = 32'd8824
; 
32'd163813: dataIn1 = 32'd8828
; 
32'd163814: dataIn1 = 32'd8830
; 
32'd163815: dataIn1 = 32'd8832
; 
32'd163816: dataIn1 = 32'd8833
; 
32'd163817: dataIn1 = 32'd6566
; 
32'd163818: dataIn1 = 32'd8822
; 
32'd163819: dataIn1 = 32'd8824
; 
32'd163820: dataIn1 = 32'd8826
; 
32'd163821: dataIn1 = 32'd8829
; 
32'd163822: dataIn1 = 32'd8836
; 
32'd163823: dataIn1 = 32'd8838
; 
32'd163824: dataIn1 = 32'd6567
; 
32'd163825: dataIn1 = 32'd8822
; 
32'd163826: dataIn1 = 32'd8823
; 
32'd163827: dataIn1 = 32'd8825
; 
32'd163828: dataIn1 = 32'd8827
; 
32'd163829: dataIn1 = 32'd8841
; 
32'd163830: dataIn1 = 32'd8842
; 
32'd163831: dataIn1 = 32'd6568
; 
32'd163832: dataIn1 = 32'd8845
; 
32'd163833: dataIn1 = 32'd8846
; 
32'd163834: dataIn1 = 32'd8850
; 
32'd163835: dataIn1 = 32'd8852
; 
32'd163836: dataIn1 = 32'd8854
; 
32'd163837: dataIn1 = 32'd8855
; 
32'd163838: dataIn1 = 32'd6569
; 
32'd163839: dataIn1 = 32'd8844
; 
32'd163840: dataIn1 = 32'd8846
; 
32'd163841: dataIn1 = 32'd8848
; 
32'd163842: dataIn1 = 32'd8851
; 
32'd163843: dataIn1 = 32'd8858
; 
32'd163844: dataIn1 = 32'd8860
; 
32'd163845: dataIn1 = 32'd6570
; 
32'd163846: dataIn1 = 32'd8844
; 
32'd163847: dataIn1 = 32'd8845
; 
32'd163848: dataIn1 = 32'd8847
; 
32'd163849: dataIn1 = 32'd8849
; 
32'd163850: dataIn1 = 32'd8863
; 
32'd163851: dataIn1 = 32'd8864
; 
32'd163852: dataIn1 = 32'd6571
; 
32'd163853: dataIn1 = 32'd8858
; 
32'd163854: dataIn1 = 32'd8859
; 
32'd163855: dataIn1 = 32'd8861
; 
32'd163856: dataIn1 = 32'd8862
; 
32'd163857: dataIn1 = 32'd9428
; 
32'd163858: dataIn1 = 32'd9429
; 
32'd163859: dataIn1 = 32'd6572
; 
32'd163860: dataIn1 = 32'd8863
; 
32'd163861: dataIn1 = 32'd8865
; 
32'd163862: dataIn1 = 32'd8866
; 
32'd163863: dataIn1 = 32'd8868
; 
32'd163864: dataIn1 = 32'd9423
; 
32'd163865: dataIn1 = 32'd9425
; 
32'd163866: dataIn1 = 32'd6573
; 
32'd163867: dataIn1 = 32'd6576
; 
32'd163868: dataIn1 = 32'd6577
; 
32'd163869: dataIn1 = 32'd8871
; 
32'd163870: dataIn1 = 32'd8872
; 
32'd163871: dataIn1 = 32'd8876
; 
32'd163872: dataIn1 = 32'd8878
; 
32'd163873: dataIn1 = 32'd6574
; 
32'd163874: dataIn1 = 32'd8870
; 
32'd163875: dataIn1 = 32'd8872
; 
32'd163876: dataIn1 = 32'd8874
; 
32'd163877: dataIn1 = 32'd8877
; 
32'd163878: dataIn1 = 32'd8879
; 
32'd163879: dataIn1 = 32'd8881
; 
32'd163880: dataIn1 = 32'd6575
; 
32'd163881: dataIn1 = 32'd8870
; 
32'd163882: dataIn1 = 32'd8871
; 
32'd163883: dataIn1 = 32'd8873
; 
32'd163884: dataIn1 = 32'd8875
; 
32'd163885: dataIn1 = 32'd8886
; 
32'd163886: dataIn1 = 32'd8887
; 
32'd163887: dataIn1 = 32'd2734
; 
32'd163888: dataIn1 = 32'd5266
; 
32'd163889: dataIn1 = 32'd6573
; 
32'd163890: dataIn1 = 32'd6576
; 
32'd163891: dataIn1 = 32'd6577
; 
32'd163892: dataIn1 = 32'd6590
; 
32'd163893: dataIn1 = 32'd6593
; 
32'd163894: dataIn1 = 32'd8878
; 
32'd163895: dataIn1 = 32'd2734
; 
32'd163896: dataIn1 = 32'd5265
; 
32'd163897: dataIn1 = 32'd6573
; 
32'd163898: dataIn1 = 32'd6576
; 
32'd163899: dataIn1 = 32'd6577
; 
32'd163900: dataIn1 = 32'd6585
; 
32'd163901: dataIn1 = 32'd6588
; 
32'd163902: dataIn1 = 32'd8876
; 
32'd163903: dataIn1 = 32'd6578
; 
32'd163904: dataIn1 = 32'd8880
; 
32'd163905: dataIn1 = 32'd8881
; 
32'd163906: dataIn1 = 32'd8884
; 
32'd163907: dataIn1 = 32'd8885
; 
32'd163908: dataIn1 = 32'd8917
; 
32'd163909: dataIn1 = 32'd8918
; 
32'd163910: dataIn1 = 32'd6579
; 
32'd163911: dataIn1 = 32'd8879
; 
32'd163912: dataIn1 = 32'd8880
; 
32'd163913: dataIn1 = 32'd8882
; 
32'd163914: dataIn1 = 32'd8883
; 
32'd163915: dataIn1 = 32'd8905
; 
32'd163916: dataIn1 = 32'd8906
; 
32'd163917: dataIn1 = 32'd6580
; 
32'd163918: dataIn1 = 32'd8887
; 
32'd163919: dataIn1 = 32'd8888
; 
32'd163920: dataIn1 = 32'd8890
; 
32'd163921: dataIn1 = 32'd8892
; 
32'd163922: dataIn1 = 32'd8912
; 
32'd163923: dataIn1 = 32'd8913
; 
32'd163924: dataIn1 = 32'd6581
; 
32'd163925: dataIn1 = 32'd8886
; 
32'd163926: dataIn1 = 32'd8888
; 
32'd163927: dataIn1 = 32'd8889
; 
32'd163928: dataIn1 = 32'd8891
; 
32'd163929: dataIn1 = 32'd8908
; 
32'd163930: dataIn1 = 32'd8910
; 
32'd163931: dataIn1 = 32'd6582
; 
32'd163932: dataIn1 = 32'd8894
; 
32'd163933: dataIn1 = 32'd8895
; 
32'd163934: dataIn1 = 32'd8899
; 
32'd163935: dataIn1 = 32'd8901
; 
32'd163936: dataIn1 = 32'd8903
; 
32'd163937: dataIn1 = 32'd8904
; 
32'd163938: dataIn1 = 32'd6583
; 
32'd163939: dataIn1 = 32'd8893
; 
32'd163940: dataIn1 = 32'd8895
; 
32'd163941: dataIn1 = 32'd8897
; 
32'd163942: dataIn1 = 32'd8900
; 
32'd163943: dataIn1 = 32'd8905
; 
32'd163944: dataIn1 = 32'd8907
; 
32'd163945: dataIn1 = 32'd6584
; 
32'd163946: dataIn1 = 32'd8893
; 
32'd163947: dataIn1 = 32'd8894
; 
32'd163948: dataIn1 = 32'd8896
; 
32'd163949: dataIn1 = 32'd8898
; 
32'd163950: dataIn1 = 32'd8908
; 
32'd163951: dataIn1 = 32'd8909
; 
32'd163952: dataIn1 = 32'd5265
; 
32'd163953: dataIn1 = 32'd5267
; 
32'd163954: dataIn1 = 32'd6577
; 
32'd163955: dataIn1 = 32'd6585
; 
32'd163956: dataIn1 = 32'd6586
; 
32'd163957: dataIn1 = 32'd6587
; 
32'd163958: dataIn1 = 32'd6588
; 
32'd163959: dataIn1 = 32'd8915
; 
32'd163960: dataIn1 = 32'd3976
; 
32'd163961: dataIn1 = 32'd5267
; 
32'd163962: dataIn1 = 32'd5870
; 
32'd163963: dataIn1 = 32'd6585
; 
32'd163964: dataIn1 = 32'd6586
; 
32'd163965: dataIn1 = 32'd6587
; 
32'd163966: dataIn1 = 32'd6589
; 
32'd163967: dataIn1 = 32'd8914
; 
32'd163968: dataIn1 = 32'd6585
; 
32'd163969: dataIn1 = 32'd6586
; 
32'd163970: dataIn1 = 32'd6587
; 
32'd163971: dataIn1 = 32'd8911
; 
32'd163972: dataIn1 = 32'd8912
; 
32'd163973: dataIn1 = 32'd8914
; 
32'd163974: dataIn1 = 32'd8915
; 
32'd163975: dataIn1 = 32'd2734
; 
32'd163976: dataIn1 = 32'd5267
; 
32'd163977: dataIn1 = 32'd6577
; 
32'd163978: dataIn1 = 32'd6585
; 
32'd163979: dataIn1 = 32'd6588
; 
32'd163980: dataIn1 = 32'd6718
; 
32'd163981: dataIn1 = 32'd452
; 
32'd163982: dataIn1 = 32'd5267
; 
32'd163983: dataIn1 = 32'd5870
; 
32'd163984: dataIn1 = 32'd6586
; 
32'd163985: dataIn1 = 32'd6589
; 
32'd163986: dataIn1 = 32'd6717
; 
32'd163987: dataIn1 = 32'd5266
; 
32'd163988: dataIn1 = 32'd5268
; 
32'd163989: dataIn1 = 32'd6576
; 
32'd163990: dataIn1 = 32'd6590
; 
32'd163991: dataIn1 = 32'd6591
; 
32'd163992: dataIn1 = 32'd6592
; 
32'd163993: dataIn1 = 32'd6593
; 
32'd163994: dataIn1 = 32'd8920
; 
32'd163995: dataIn1 = 32'd6590
; 
32'd163996: dataIn1 = 32'd6591
; 
32'd163997: dataIn1 = 32'd6592
; 
32'd163998: dataIn1 = 32'd8916
; 
32'd163999: dataIn1 = 32'd8918
; 
32'd164000: dataIn1 = 32'd8919
; 
32'd164001: dataIn1 = 32'd8920
; 
32'd164002: dataIn1 = 32'd5129
; 
32'd164003: dataIn1 = 32'd5268
; 
32'd164004: dataIn1 = 32'd6131
; 
32'd164005: dataIn1 = 32'd6590
; 
32'd164006: dataIn1 = 32'd6591
; 
32'd164007: dataIn1 = 32'd6592
; 
32'd164008: dataIn1 = 32'd6594
; 
32'd164009: dataIn1 = 32'd8919
; 
32'd164010: dataIn1 = 32'd2734
; 
32'd164011: dataIn1 = 32'd5268
; 
32'd164012: dataIn1 = 32'd6576
; 
32'd164013: dataIn1 = 32'd6590
; 
32'd164014: dataIn1 = 32'd6593
; 
32'd164015: dataIn1 = 32'd6720
; 
32'd164016: dataIn1 = 32'd1119
; 
32'd164017: dataIn1 = 32'd5268
; 
32'd164018: dataIn1 = 32'd6131
; 
32'd164019: dataIn1 = 32'd6592
; 
32'd164020: dataIn1 = 32'd6594
; 
32'd164021: dataIn1 = 32'd6719
; 
32'd164022: dataIn1 = 32'd6595
; 
32'd164023: dataIn1 = 32'd8922
; 
32'd164024: dataIn1 = 32'd8923
; 
32'd164025: dataIn1 = 32'd8926
; 
32'd164026: dataIn1 = 32'd9743
; 
32'd164027: dataIn1 = 32'd9744
; 
32'd164028: dataIn1 = 32'd9746
; 
32'd164029: dataIn1 = 32'd5269
; 
32'd164030: dataIn1 = 32'd6596
; 
32'd164031: dataIn1 = 32'd6598
; 
32'd164032: dataIn1 = 32'd9742
; 
32'd164033: dataIn1 = 32'd9744
; 
32'd164034: dataIn1 = 32'd9768
; 
32'd164035: dataIn1 = 32'd9779
; 
32'd164036: dataIn1 = 32'd5269
; 
32'd164037: dataIn1 = 32'd6597
; 
32'd164038: dataIn1 = 32'd9671
; 
32'd164039: dataIn1 = 32'd9742
; 
32'd164040: dataIn1 = 32'd9743
; 
32'd164041: dataIn1 = 32'd9745
; 
32'd164042: dataIn1 = 32'd10134
; 
32'd164043: dataIn1 = 32'd2325
; 
32'd164044: dataIn1 = 32'd5269
; 
32'd164045: dataIn1 = 32'd5271
; 
32'd164046: dataIn1 = 32'd5887
; 
32'd164047: dataIn1 = 32'd6596
; 
32'd164048: dataIn1 = 32'd6598
; 
32'd164049: dataIn1 = 32'd9779
; 
32'd164050: dataIn1 = 32'd6599
; 
32'd164051: dataIn1 = 32'd8928
; 
32'd164052: dataIn1 = 32'd8929
; 
32'd164053: dataIn1 = 32'd8933
; 
32'd164054: dataIn1 = 32'd8935
; 
32'd164055: dataIn1 = 32'd9277
; 
32'd164056: dataIn1 = 32'd9278
; 
32'd164057: dataIn1 = 32'd6600
; 
32'd164058: dataIn1 = 32'd8927
; 
32'd164059: dataIn1 = 32'd8929
; 
32'd164060: dataIn1 = 32'd8931
; 
32'd164061: dataIn1 = 32'd8934
; 
32'd164062: dataIn1 = 32'd8936
; 
32'd164063: dataIn1 = 32'd8938
; 
32'd164064: dataIn1 = 32'd6601
; 
32'd164065: dataIn1 = 32'd8927
; 
32'd164066: dataIn1 = 32'd8928
; 
32'd164067: dataIn1 = 32'd8930
; 
32'd164068: dataIn1 = 32'd8932
; 
32'd164069: dataIn1 = 32'd8943
; 
32'd164070: dataIn1 = 32'd8944
; 
32'd164071: dataIn1 = 32'd6602
; 
32'd164072: dataIn1 = 32'd6610
; 
32'd164073: dataIn1 = 32'd8937
; 
32'd164074: dataIn1 = 32'd8938
; 
32'd164075: dataIn1 = 32'd8941
; 
32'd164076: dataIn1 = 32'd8942
; 
32'd164077: dataIn1 = 32'd8975
; 
32'd164078: dataIn1 = 32'd6603
; 
32'd164079: dataIn1 = 32'd8936
; 
32'd164080: dataIn1 = 32'd8937
; 
32'd164081: dataIn1 = 32'd8939
; 
32'd164082: dataIn1 = 32'd8940
; 
32'd164083: dataIn1 = 32'd8964
; 
32'd164084: dataIn1 = 32'd8965
; 
32'd164085: dataIn1 = 32'd6604
; 
32'd164086: dataIn1 = 32'd8944
; 
32'd164087: dataIn1 = 32'd8945
; 
32'd164088: dataIn1 = 32'd8947
; 
32'd164089: dataIn1 = 32'd8949
; 
32'd164090: dataIn1 = 32'd8971
; 
32'd164091: dataIn1 = 32'd8972
; 
32'd164092: dataIn1 = 32'd6605
; 
32'd164093: dataIn1 = 32'd8943
; 
32'd164094: dataIn1 = 32'd8945
; 
32'd164095: dataIn1 = 32'd8946
; 
32'd164096: dataIn1 = 32'd8948
; 
32'd164097: dataIn1 = 32'd8967
; 
32'd164098: dataIn1 = 32'd8969
; 
32'd164099: dataIn1 = 32'd6606
; 
32'd164100: dataIn1 = 32'd8951
; 
32'd164101: dataIn1 = 32'd8952
; 
32'd164102: dataIn1 = 32'd8956
; 
32'd164103: dataIn1 = 32'd8958
; 
32'd164104: dataIn1 = 32'd8960
; 
32'd164105: dataIn1 = 32'd8961
; 
32'd164106: dataIn1 = 32'd6607
; 
32'd164107: dataIn1 = 32'd8950
; 
32'd164108: dataIn1 = 32'd8952
; 
32'd164109: dataIn1 = 32'd8954
; 
32'd164110: dataIn1 = 32'd8957
; 
32'd164111: dataIn1 = 32'd8964
; 
32'd164112: dataIn1 = 32'd8966
; 
32'd164113: dataIn1 = 32'd6608
; 
32'd164114: dataIn1 = 32'd8950
; 
32'd164115: dataIn1 = 32'd8951
; 
32'd164116: dataIn1 = 32'd8953
; 
32'd164117: dataIn1 = 32'd8955
; 
32'd164118: dataIn1 = 32'd8967
; 
32'd164119: dataIn1 = 32'd8968
; 
32'd164120: dataIn1 = 32'd6609
; 
32'd164121: dataIn1 = 32'd8970
; 
32'd164122: dataIn1 = 32'd8971
; 
32'd164123: dataIn1 = 32'd8973
; 
32'd164124: dataIn1 = 32'd8974
; 
32'd164125: dataIn1 = 32'd9279
; 
32'd164126: dataIn1 = 32'd9280
; 
32'd164127: dataIn1 = 32'd5148
; 
32'd164128: dataIn1 = 32'd5276
; 
32'd164129: dataIn1 = 32'd5278
; 
32'd164130: dataIn1 = 32'd6180
; 
32'd164131: dataIn1 = 32'd6602
; 
32'd164132: dataIn1 = 32'd6610
; 
32'd164133: dataIn1 = 32'd8942
; 
32'd164134: dataIn1 = 32'd8975
; 
32'd164135: dataIn1 = 32'd6611
; 
32'd164136: dataIn1 = 32'd6786
; 
32'd164137: dataIn1 = 32'd6787
; 
32'd164138: dataIn1 = 32'd8977
; 
32'd164139: dataIn1 = 32'd8978
; 
32'd164140: dataIn1 = 32'd8982
; 
32'd164141: dataIn1 = 32'd8984
; 
32'd164142: dataIn1 = 32'd6612
; 
32'd164143: dataIn1 = 32'd8976
; 
32'd164144: dataIn1 = 32'd8978
; 
32'd164145: dataIn1 = 32'd8980
; 
32'd164146: dataIn1 = 32'd8983
; 
32'd164147: dataIn1 = 32'd8985
; 
32'd164148: dataIn1 = 32'd8987
; 
32'd164149: dataIn1 = 32'd6613
; 
32'd164150: dataIn1 = 32'd8976
; 
32'd164151: dataIn1 = 32'd8977
; 
32'd164152: dataIn1 = 32'd8979
; 
32'd164153: dataIn1 = 32'd8981
; 
32'd164154: dataIn1 = 32'd8992
; 
32'd164155: dataIn1 = 32'd8993
; 
32'd164156: dataIn1 = 32'd6614
; 
32'd164157: dataIn1 = 32'd8986
; 
32'd164158: dataIn1 = 32'd8987
; 
32'd164159: dataIn1 = 32'd8990
; 
32'd164160: dataIn1 = 32'd8991
; 
32'd164161: dataIn1 = 32'd9023
; 
32'd164162: dataIn1 = 32'd9024
; 
32'd164163: dataIn1 = 32'd6615
; 
32'd164164: dataIn1 = 32'd8985
; 
32'd164165: dataIn1 = 32'd8986
; 
32'd164166: dataIn1 = 32'd8988
; 
32'd164167: dataIn1 = 32'd8989
; 
32'd164168: dataIn1 = 32'd9011
; 
32'd164169: dataIn1 = 32'd9012
; 
32'd164170: dataIn1 = 32'd6616
; 
32'd164171: dataIn1 = 32'd8993
; 
32'd164172: dataIn1 = 32'd8994
; 
32'd164173: dataIn1 = 32'd8996
; 
32'd164174: dataIn1 = 32'd8998
; 
32'd164175: dataIn1 = 32'd9018
; 
32'd164176: dataIn1 = 32'd9019
; 
32'd164177: dataIn1 = 32'd6617
; 
32'd164178: dataIn1 = 32'd8992
; 
32'd164179: dataIn1 = 32'd8994
; 
32'd164180: dataIn1 = 32'd8995
; 
32'd164181: dataIn1 = 32'd8997
; 
32'd164182: dataIn1 = 32'd9014
; 
32'd164183: dataIn1 = 32'd9016
; 
32'd164184: dataIn1 = 32'd6618
; 
32'd164185: dataIn1 = 32'd9000
; 
32'd164186: dataIn1 = 32'd9001
; 
32'd164187: dataIn1 = 32'd9005
; 
32'd164188: dataIn1 = 32'd9007
; 
32'd164189: dataIn1 = 32'd9009
; 
32'd164190: dataIn1 = 32'd9010
; 
32'd164191: dataIn1 = 32'd6619
; 
32'd164192: dataIn1 = 32'd8999
; 
32'd164193: dataIn1 = 32'd9001
; 
32'd164194: dataIn1 = 32'd9003
; 
32'd164195: dataIn1 = 32'd9006
; 
32'd164196: dataIn1 = 32'd9011
; 
32'd164197: dataIn1 = 32'd9013
; 
32'd164198: dataIn1 = 32'd6620
; 
32'd164199: dataIn1 = 32'd8999
; 
32'd164200: dataIn1 = 32'd9000
; 
32'd164201: dataIn1 = 32'd9002
; 
32'd164202: dataIn1 = 32'd9004
; 
32'd164203: dataIn1 = 32'd9014
; 
32'd164204: dataIn1 = 32'd9015
; 
32'd164205: dataIn1 = 32'd6621
; 
32'd164206: dataIn1 = 32'd6788
; 
32'd164207: dataIn1 = 32'd6789
; 
32'd164208: dataIn1 = 32'd9017
; 
32'd164209: dataIn1 = 32'd9018
; 
32'd164210: dataIn1 = 32'd9020
; 
32'd164211: dataIn1 = 32'd9021
; 
32'd164212: dataIn1 = 32'd6622
; 
32'd164213: dataIn1 = 32'd6790
; 
32'd164214: dataIn1 = 32'd6791
; 
32'd164215: dataIn1 = 32'd9022
; 
32'd164216: dataIn1 = 32'd9024
; 
32'd164217: dataIn1 = 32'd9025
; 
32'd164218: dataIn1 = 32'd9026
; 
32'd164219: dataIn1 = 32'd6623
; 
32'd164220: dataIn1 = 32'd6626
; 
32'd164221: dataIn1 = 32'd6627
; 
32'd164222: dataIn1 = 32'd9028
; 
32'd164223: dataIn1 = 32'd9029
; 
32'd164224: dataIn1 = 32'd9033
; 
32'd164225: dataIn1 = 32'd9035
; 
32'd164226: dataIn1 = 32'd6624
; 
32'd164227: dataIn1 = 32'd9027
; 
32'd164228: dataIn1 = 32'd9029
; 
32'd164229: dataIn1 = 32'd9031
; 
32'd164230: dataIn1 = 32'd9034
; 
32'd164231: dataIn1 = 32'd9037
; 
32'd164232: dataIn1 = 32'd9039
; 
32'd164233: dataIn1 = 32'd6625
; 
32'd164234: dataIn1 = 32'd9027
; 
32'd164235: dataIn1 = 32'd9028
; 
32'd164236: dataIn1 = 32'd9030
; 
32'd164237: dataIn1 = 32'd9032
; 
32'd164238: dataIn1 = 32'd9044
; 
32'd164239: dataIn1 = 32'd9045
; 
32'd164240: dataIn1 = 32'd2749
; 
32'd164241: dataIn1 = 32'd5286
; 
32'd164242: dataIn1 = 32'd6623
; 
32'd164243: dataIn1 = 32'd6626
; 
32'd164244: dataIn1 = 32'd6627
; 
32'd164245: dataIn1 = 32'd6792
; 
32'd164246: dataIn1 = 32'd9035
; 
32'd164247: dataIn1 = 32'd9036
; 
32'd164248: dataIn1 = 32'd2749
; 
32'd164249: dataIn1 = 32'd5285
; 
32'd164250: dataIn1 = 32'd6623
; 
32'd164251: dataIn1 = 32'd6626
; 
32'd164252: dataIn1 = 32'd6627
; 
32'd164253: dataIn1 = 32'd6635
; 
32'd164254: dataIn1 = 32'd6636
; 
32'd164255: dataIn1 = 32'd9033
; 
32'd164256: dataIn1 = 32'd6628
; 
32'd164257: dataIn1 = 32'd9038
; 
32'd164258: dataIn1 = 32'd9039
; 
32'd164259: dataIn1 = 32'd9042
; 
32'd164260: dataIn1 = 32'd9043
; 
32'd164261: dataIn1 = 32'd9075
; 
32'd164262: dataIn1 = 32'd9076
; 
32'd164263: dataIn1 = 32'd6629
; 
32'd164264: dataIn1 = 32'd9037
; 
32'd164265: dataIn1 = 32'd9038
; 
32'd164266: dataIn1 = 32'd9040
; 
32'd164267: dataIn1 = 32'd9041
; 
32'd164268: dataIn1 = 32'd9063
; 
32'd164269: dataIn1 = 32'd9064
; 
32'd164270: dataIn1 = 32'd6630
; 
32'd164271: dataIn1 = 32'd9045
; 
32'd164272: dataIn1 = 32'd9046
; 
32'd164273: dataIn1 = 32'd9048
; 
32'd164274: dataIn1 = 32'd9050
; 
32'd164275: dataIn1 = 32'd9070
; 
32'd164276: dataIn1 = 32'd9071
; 
32'd164277: dataIn1 = 32'd6631
; 
32'd164278: dataIn1 = 32'd9044
; 
32'd164279: dataIn1 = 32'd9046
; 
32'd164280: dataIn1 = 32'd9047
; 
32'd164281: dataIn1 = 32'd9049
; 
32'd164282: dataIn1 = 32'd9066
; 
32'd164283: dataIn1 = 32'd9068
; 
32'd164284: dataIn1 = 32'd6632
; 
32'd164285: dataIn1 = 32'd9052
; 
32'd164286: dataIn1 = 32'd9053
; 
32'd164287: dataIn1 = 32'd9057
; 
32'd164288: dataIn1 = 32'd9059
; 
32'd164289: dataIn1 = 32'd9061
; 
32'd164290: dataIn1 = 32'd9062
; 
32'd164291: dataIn1 = 32'd6633
; 
32'd164292: dataIn1 = 32'd9051
; 
32'd164293: dataIn1 = 32'd9053
; 
32'd164294: dataIn1 = 32'd9055
; 
32'd164295: dataIn1 = 32'd9058
; 
32'd164296: dataIn1 = 32'd9063
; 
32'd164297: dataIn1 = 32'd9065
; 
32'd164298: dataIn1 = 32'd6634
; 
32'd164299: dataIn1 = 32'd9051
; 
32'd164300: dataIn1 = 32'd9052
; 
32'd164301: dataIn1 = 32'd9054
; 
32'd164302: dataIn1 = 32'd9056
; 
32'd164303: dataIn1 = 32'd9066
; 
32'd164304: dataIn1 = 32'd9067
; 
32'd164305: dataIn1 = 32'd5285
; 
32'd164306: dataIn1 = 32'd5287
; 
32'd164307: dataIn1 = 32'd6627
; 
32'd164308: dataIn1 = 32'd6635
; 
32'd164309: dataIn1 = 32'd6636
; 
32'd164310: dataIn1 = 32'd6638
; 
32'd164311: dataIn1 = 32'd6639
; 
32'd164312: dataIn1 = 32'd9073
; 
32'd164313: dataIn1 = 32'd2749
; 
32'd164314: dataIn1 = 32'd5287
; 
32'd164315: dataIn1 = 32'd6627
; 
32'd164316: dataIn1 = 32'd6635
; 
32'd164317: dataIn1 = 32'd6636
; 
32'd164318: dataIn1 = 32'd6722
; 
32'd164319: dataIn1 = 32'd1128
; 
32'd164320: dataIn1 = 32'd5287
; 
32'd164321: dataIn1 = 32'd6360
; 
32'd164322: dataIn1 = 32'd6637
; 
32'd164323: dataIn1 = 32'd6638
; 
32'd164324: dataIn1 = 32'd6721
; 
32'd164325: dataIn1 = 32'd5201
; 
32'd164326: dataIn1 = 32'd5287
; 
32'd164327: dataIn1 = 32'd6360
; 
32'd164328: dataIn1 = 32'd6635
; 
32'd164329: dataIn1 = 32'd6637
; 
32'd164330: dataIn1 = 32'd6638
; 
32'd164331: dataIn1 = 32'd6639
; 
32'd164332: dataIn1 = 32'd9072
; 
32'd164333: dataIn1 = 32'd6635
; 
32'd164334: dataIn1 = 32'd6638
; 
32'd164335: dataIn1 = 32'd6639
; 
32'd164336: dataIn1 = 32'd9069
; 
32'd164337: dataIn1 = 32'd9070
; 
32'd164338: dataIn1 = 32'd9072
; 
32'd164339: dataIn1 = 32'd9073
; 
32'd164340: dataIn1 = 32'd6640
; 
32'd164341: dataIn1 = 32'd6792
; 
32'd164342: dataIn1 = 32'd6793
; 
32'd164343: dataIn1 = 32'd9074
; 
32'd164344: dataIn1 = 32'd9076
; 
32'd164345: dataIn1 = 32'd9077
; 
32'd164346: dataIn1 = 32'd9078
; 
32'd164347: dataIn1 = 32'd6641
; 
32'd164348: dataIn1 = 32'd6644
; 
32'd164349: dataIn1 = 32'd6645
; 
32'd164350: dataIn1 = 32'd9080
; 
32'd164351: dataIn1 = 32'd9081
; 
32'd164352: dataIn1 = 32'd9085
; 
32'd164353: dataIn1 = 32'd9087
; 
32'd164354: dataIn1 = 32'd6642
; 
32'd164355: dataIn1 = 32'd9079
; 
32'd164356: dataIn1 = 32'd9081
; 
32'd164357: dataIn1 = 32'd9083
; 
32'd164358: dataIn1 = 32'd9086
; 
32'd164359: dataIn1 = 32'd9088
; 
32'd164360: dataIn1 = 32'd9090
; 
32'd164361: dataIn1 = 32'd6643
; 
32'd164362: dataIn1 = 32'd9079
; 
32'd164363: dataIn1 = 32'd9080
; 
32'd164364: dataIn1 = 32'd9082
; 
32'd164365: dataIn1 = 32'd9084
; 
32'd164366: dataIn1 = 32'd9095
; 
32'd164367: dataIn1 = 32'd9096
; 
32'd164368: dataIn1 = 32'd2750
; 
32'd164369: dataIn1 = 32'd5291
; 
32'd164370: dataIn1 = 32'd6641
; 
32'd164371: dataIn1 = 32'd6644
; 
32'd164372: dataIn1 = 32'd6645
; 
32'd164373: dataIn1 = 32'd6656
; 
32'd164374: dataIn1 = 32'd6657
; 
32'd164375: dataIn1 = 32'd9087
; 
32'd164376: dataIn1 = 32'd2750
; 
32'd164377: dataIn1 = 32'd5290
; 
32'd164378: dataIn1 = 32'd6641
; 
32'd164379: dataIn1 = 32'd6644
; 
32'd164380: dataIn1 = 32'd6645
; 
32'd164381: dataIn1 = 32'd6653
; 
32'd164382: dataIn1 = 32'd6654
; 
32'd164383: dataIn1 = 32'd9085
; 
32'd164384: dataIn1 = 32'd6646
; 
32'd164385: dataIn1 = 32'd9089
; 
32'd164386: dataIn1 = 32'd9090
; 
32'd164387: dataIn1 = 32'd9093
; 
32'd164388: dataIn1 = 32'd9094
; 
32'd164389: dataIn1 = 32'd9126
; 
32'd164390: dataIn1 = 32'd9127
; 
32'd164391: dataIn1 = 32'd6647
; 
32'd164392: dataIn1 = 32'd9088
; 
32'd164393: dataIn1 = 32'd9089
; 
32'd164394: dataIn1 = 32'd9091
; 
32'd164395: dataIn1 = 32'd9092
; 
32'd164396: dataIn1 = 32'd9114
; 
32'd164397: dataIn1 = 32'd9115
; 
32'd164398: dataIn1 = 32'd6648
; 
32'd164399: dataIn1 = 32'd9096
; 
32'd164400: dataIn1 = 32'd9097
; 
32'd164401: dataIn1 = 32'd9099
; 
32'd164402: dataIn1 = 32'd9101
; 
32'd164403: dataIn1 = 32'd9121
; 
32'd164404: dataIn1 = 32'd9122
; 
32'd164405: dataIn1 = 32'd6649
; 
32'd164406: dataIn1 = 32'd9095
; 
32'd164407: dataIn1 = 32'd9097
; 
32'd164408: dataIn1 = 32'd9098
; 
32'd164409: dataIn1 = 32'd9100
; 
32'd164410: dataIn1 = 32'd9117
; 
32'd164411: dataIn1 = 32'd9119
; 
32'd164412: dataIn1 = 32'd6650
; 
32'd164413: dataIn1 = 32'd9103
; 
32'd164414: dataIn1 = 32'd9104
; 
32'd164415: dataIn1 = 32'd9108
; 
32'd164416: dataIn1 = 32'd9110
; 
32'd164417: dataIn1 = 32'd9112
; 
32'd164418: dataIn1 = 32'd9113
; 
32'd164419: dataIn1 = 32'd6651
; 
32'd164420: dataIn1 = 32'd9102
; 
32'd164421: dataIn1 = 32'd9104
; 
32'd164422: dataIn1 = 32'd9106
; 
32'd164423: dataIn1 = 32'd9109
; 
32'd164424: dataIn1 = 32'd9114
; 
32'd164425: dataIn1 = 32'd9116
; 
32'd164426: dataIn1 = 32'd6652
; 
32'd164427: dataIn1 = 32'd9102
; 
32'd164428: dataIn1 = 32'd9103
; 
32'd164429: dataIn1 = 32'd9105
; 
32'd164430: dataIn1 = 32'd9107
; 
32'd164431: dataIn1 = 32'd9117
; 
32'd164432: dataIn1 = 32'd9118
; 
32'd164433: dataIn1 = 32'd5290
; 
32'd164434: dataIn1 = 32'd5292
; 
32'd164435: dataIn1 = 32'd6645
; 
32'd164436: dataIn1 = 32'd6653
; 
32'd164437: dataIn1 = 32'd6654
; 
32'd164438: dataIn1 = 32'd6655
; 
32'd164439: dataIn1 = 32'd6725
; 
32'd164440: dataIn1 = 32'd9124
; 
32'd164441: dataIn1 = 32'd2750
; 
32'd164442: dataIn1 = 32'd5292
; 
32'd164443: dataIn1 = 32'd6645
; 
32'd164444: dataIn1 = 32'd6653
; 
32'd164445: dataIn1 = 32'd6654
; 
32'd164446: dataIn1 = 32'd6724
; 
32'd164447: dataIn1 = 32'd6653
; 
32'd164448: dataIn1 = 32'd6655
; 
32'd164449: dataIn1 = 32'd6725
; 
32'd164450: dataIn1 = 32'd9120
; 
32'd164451: dataIn1 = 32'd9121
; 
32'd164452: dataIn1 = 32'd9123
; 
32'd164453: dataIn1 = 32'd9124
; 
32'd164454: dataIn1 = 32'd5291
; 
32'd164455: dataIn1 = 32'd5293
; 
32'd164456: dataIn1 = 32'd6644
; 
32'd164457: dataIn1 = 32'd6656
; 
32'd164458: dataIn1 = 32'd6657
; 
32'd164459: dataIn1 = 32'd6658
; 
32'd164460: dataIn1 = 32'd6660
; 
32'd164461: dataIn1 = 32'd9129
; 
32'd164462: dataIn1 = 32'd2750
; 
32'd164463: dataIn1 = 32'd5293
; 
32'd164464: dataIn1 = 32'd6644
; 
32'd164465: dataIn1 = 32'd6656
; 
32'd164466: dataIn1 = 32'd6657
; 
32'd164467: dataIn1 = 32'd6727
; 
32'd164468: dataIn1 = 32'd6656
; 
32'd164469: dataIn1 = 32'd6658
; 
32'd164470: dataIn1 = 32'd6660
; 
32'd164471: dataIn1 = 32'd9125
; 
32'd164472: dataIn1 = 32'd9127
; 
32'd164473: dataIn1 = 32'd9128
; 
32'd164474: dataIn1 = 32'd9129
; 
32'd164475: dataIn1 = 32'd1127
; 
32'd164476: dataIn1 = 32'd5293
; 
32'd164477: dataIn1 = 32'd6373
; 
32'd164478: dataIn1 = 32'd6659
; 
32'd164479: dataIn1 = 32'd6660
; 
32'd164480: dataIn1 = 32'd6726
; 
32'd164481: dataIn1 = 32'd5205
; 
32'd164482: dataIn1 = 32'd5293
; 
32'd164483: dataIn1 = 32'd6373
; 
32'd164484: dataIn1 = 32'd6656
; 
32'd164485: dataIn1 = 32'd6658
; 
32'd164486: dataIn1 = 32'd6659
; 
32'd164487: dataIn1 = 32'd6660
; 
32'd164488: dataIn1 = 32'd9128
; 
32'd164489: dataIn1 = 32'd6661
; 
32'd164490: dataIn1 = 32'd6664
; 
32'd164491: dataIn1 = 32'd6665
; 
32'd164492: dataIn1 = 32'd9131
; 
32'd164493: dataIn1 = 32'd9132
; 
32'd164494: dataIn1 = 32'd9136
; 
32'd164495: dataIn1 = 32'd9138
; 
32'd164496: dataIn1 = 32'd6662
; 
32'd164497: dataIn1 = 32'd9130
; 
32'd164498: dataIn1 = 32'd9132
; 
32'd164499: dataIn1 = 32'd9134
; 
32'd164500: dataIn1 = 32'd9137
; 
32'd164501: dataIn1 = 32'd9140
; 
32'd164502: dataIn1 = 32'd9142
; 
32'd164503: dataIn1 = 32'd6663
; 
32'd164504: dataIn1 = 32'd9130
; 
32'd164505: dataIn1 = 32'd9131
; 
32'd164506: dataIn1 = 32'd9133
; 
32'd164507: dataIn1 = 32'd9135
; 
32'd164508: dataIn1 = 32'd9147
; 
32'd164509: dataIn1 = 32'd9148
; 
32'd164510: dataIn1 = 32'd2751
; 
32'd164511: dataIn1 = 32'd5296
; 
32'd164512: dataIn1 = 32'd6661
; 
32'd164513: dataIn1 = 32'd6664
; 
32'd164514: dataIn1 = 32'd6665
; 
32'd164515: dataIn1 = 32'd6674
; 
32'd164516: dataIn1 = 32'd6677
; 
32'd164517: dataIn1 = 32'd9138
; 
32'd164518: dataIn1 = 32'd2751
; 
32'd164519: dataIn1 = 32'd5295
; 
32'd164520: dataIn1 = 32'd6661
; 
32'd164521: dataIn1 = 32'd6664
; 
32'd164522: dataIn1 = 32'd6665
; 
32'd164523: dataIn1 = 32'd6794
; 
32'd164524: dataIn1 = 32'd9136
; 
32'd164525: dataIn1 = 32'd9139
; 
32'd164526: dataIn1 = 32'd6666
; 
32'd164527: dataIn1 = 32'd9141
; 
32'd164528: dataIn1 = 32'd9142
; 
32'd164529: dataIn1 = 32'd9145
; 
32'd164530: dataIn1 = 32'd9146
; 
32'd164531: dataIn1 = 32'd9178
; 
32'd164532: dataIn1 = 32'd9179
; 
32'd164533: dataIn1 = 32'd6667
; 
32'd164534: dataIn1 = 32'd9140
; 
32'd164535: dataIn1 = 32'd9141
; 
32'd164536: dataIn1 = 32'd9143
; 
32'd164537: dataIn1 = 32'd9144
; 
32'd164538: dataIn1 = 32'd9166
; 
32'd164539: dataIn1 = 32'd9167
; 
32'd164540: dataIn1 = 32'd6668
; 
32'd164541: dataIn1 = 32'd9148
; 
32'd164542: dataIn1 = 32'd9149
; 
32'd164543: dataIn1 = 32'd9151
; 
32'd164544: dataIn1 = 32'd9153
; 
32'd164545: dataIn1 = 32'd9173
; 
32'd164546: dataIn1 = 32'd9174
; 
32'd164547: dataIn1 = 32'd6669
; 
32'd164548: dataIn1 = 32'd9147
; 
32'd164549: dataIn1 = 32'd9149
; 
32'd164550: dataIn1 = 32'd9150
; 
32'd164551: dataIn1 = 32'd9152
; 
32'd164552: dataIn1 = 32'd9169
; 
32'd164553: dataIn1 = 32'd9171
; 
32'd164554: dataIn1 = 32'd6670
; 
32'd164555: dataIn1 = 32'd9155
; 
32'd164556: dataIn1 = 32'd9156
; 
32'd164557: dataIn1 = 32'd9160
; 
32'd164558: dataIn1 = 32'd9162
; 
32'd164559: dataIn1 = 32'd9164
; 
32'd164560: dataIn1 = 32'd9165
; 
32'd164561: dataIn1 = 32'd6671
; 
32'd164562: dataIn1 = 32'd9154
; 
32'd164563: dataIn1 = 32'd9156
; 
32'd164564: dataIn1 = 32'd9158
; 
32'd164565: dataIn1 = 32'd9161
; 
32'd164566: dataIn1 = 32'd9166
; 
32'd164567: dataIn1 = 32'd9168
; 
32'd164568: dataIn1 = 32'd6672
; 
32'd164569: dataIn1 = 32'd9154
; 
32'd164570: dataIn1 = 32'd9155
; 
32'd164571: dataIn1 = 32'd9157
; 
32'd164572: dataIn1 = 32'd9159
; 
32'd164573: dataIn1 = 32'd9169
; 
32'd164574: dataIn1 = 32'd9170
; 
32'd164575: dataIn1 = 32'd6673
; 
32'd164576: dataIn1 = 32'd6794
; 
32'd164577: dataIn1 = 32'd6795
; 
32'd164578: dataIn1 = 32'd9172
; 
32'd164579: dataIn1 = 32'd9173
; 
32'd164580: dataIn1 = 32'd9175
; 
32'd164581: dataIn1 = 32'd9176
; 
32'd164582: dataIn1 = 32'd5296
; 
32'd164583: dataIn1 = 32'd5298
; 
32'd164584: dataIn1 = 32'd6664
; 
32'd164585: dataIn1 = 32'd6674
; 
32'd164586: dataIn1 = 32'd6675
; 
32'd164587: dataIn1 = 32'd6676
; 
32'd164588: dataIn1 = 32'd6677
; 
32'd164589: dataIn1 = 32'd9180
; 
32'd164590: dataIn1 = 32'd6674
; 
32'd164591: dataIn1 = 32'd6675
; 
32'd164592: dataIn1 = 32'd6676
; 
32'd164593: dataIn1 = 32'd9177
; 
32'd164594: dataIn1 = 32'd9179
; 
32'd164595: dataIn1 = 32'd9180
; 
32'd164596: dataIn1 = 32'd9285
; 
32'd164597: dataIn1 = 32'd5224
; 
32'd164598: dataIn1 = 32'd5298
; 
32'd164599: dataIn1 = 32'd6443
; 
32'd164600: dataIn1 = 32'd6674
; 
32'd164601: dataIn1 = 32'd6675
; 
32'd164602: dataIn1 = 32'd6676
; 
32'd164603: dataIn1 = 32'd6678
; 
32'd164604: dataIn1 = 32'd9285
; 
32'd164605: dataIn1 = 32'd2751
; 
32'd164606: dataIn1 = 32'd5298
; 
32'd164607: dataIn1 = 32'd6664
; 
32'd164608: dataIn1 = 32'd6674
; 
32'd164609: dataIn1 = 32'd6677
; 
32'd164610: dataIn1 = 32'd6729
; 
32'd164611: dataIn1 = 32'd1129
; 
32'd164612: dataIn1 = 32'd5298
; 
32'd164613: dataIn1 = 32'd6443
; 
32'd164614: dataIn1 = 32'd6676
; 
32'd164615: dataIn1 = 32'd6678
; 
32'd164616: dataIn1 = 32'd10222
; 
32'd164617: dataIn1 = 32'd10246
; 
32'd164618: dataIn1 = 32'd6679
; 
32'd164619: dataIn1 = 32'd6796
; 
32'd164620: dataIn1 = 32'd6797
; 
32'd164621: dataIn1 = 32'd9182
; 
32'd164622: dataIn1 = 32'd9183
; 
32'd164623: dataIn1 = 32'd9187
; 
32'd164624: dataIn1 = 32'd9189
; 
32'd164625: dataIn1 = 32'd6680
; 
32'd164626: dataIn1 = 32'd9181
; 
32'd164627: dataIn1 = 32'd9183
; 
32'd164628: dataIn1 = 32'd9185
; 
32'd164629: dataIn1 = 32'd9188
; 
32'd164630: dataIn1 = 32'd9190
; 
32'd164631: dataIn1 = 32'd9192
; 
32'd164632: dataIn1 = 32'd6681
; 
32'd164633: dataIn1 = 32'd9181
; 
32'd164634: dataIn1 = 32'd9182
; 
32'd164635: dataIn1 = 32'd9184
; 
32'd164636: dataIn1 = 32'd9186
; 
32'd164637: dataIn1 = 32'd9197
; 
32'd164638: dataIn1 = 32'd9198
; 
32'd164639: dataIn1 = 32'd6682
; 
32'd164640: dataIn1 = 32'd9191
; 
32'd164641: dataIn1 = 32'd9192
; 
32'd164642: dataIn1 = 32'd9195
; 
32'd164643: dataIn1 = 32'd9196
; 
32'd164644: dataIn1 = 32'd9228
; 
32'd164645: dataIn1 = 32'd9229
; 
32'd164646: dataIn1 = 32'd6683
; 
32'd164647: dataIn1 = 32'd9190
; 
32'd164648: dataIn1 = 32'd9191
; 
32'd164649: dataIn1 = 32'd9193
; 
32'd164650: dataIn1 = 32'd9194
; 
32'd164651: dataIn1 = 32'd9216
; 
32'd164652: dataIn1 = 32'd9217
; 
32'd164653: dataIn1 = 32'd6684
; 
32'd164654: dataIn1 = 32'd9198
; 
32'd164655: dataIn1 = 32'd9199
; 
32'd164656: dataIn1 = 32'd9201
; 
32'd164657: dataIn1 = 32'd9203
; 
32'd164658: dataIn1 = 32'd9223
; 
32'd164659: dataIn1 = 32'd9224
; 
32'd164660: dataIn1 = 32'd6685
; 
32'd164661: dataIn1 = 32'd9197
; 
32'd164662: dataIn1 = 32'd9199
; 
32'd164663: dataIn1 = 32'd9200
; 
32'd164664: dataIn1 = 32'd9202
; 
32'd164665: dataIn1 = 32'd9219
; 
32'd164666: dataIn1 = 32'd9221
; 
32'd164667: dataIn1 = 32'd6686
; 
32'd164668: dataIn1 = 32'd9205
; 
32'd164669: dataIn1 = 32'd9206
; 
32'd164670: dataIn1 = 32'd9210
; 
32'd164671: dataIn1 = 32'd9212
; 
32'd164672: dataIn1 = 32'd9214
; 
32'd164673: dataIn1 = 32'd9215
; 
32'd164674: dataIn1 = 32'd6687
; 
32'd164675: dataIn1 = 32'd9204
; 
32'd164676: dataIn1 = 32'd9206
; 
32'd164677: dataIn1 = 32'd9208
; 
32'd164678: dataIn1 = 32'd9211
; 
32'd164679: dataIn1 = 32'd9216
; 
32'd164680: dataIn1 = 32'd9218
; 
32'd164681: dataIn1 = 32'd6688
; 
32'd164682: dataIn1 = 32'd9204
; 
32'd164683: dataIn1 = 32'd9205
; 
32'd164684: dataIn1 = 32'd9207
; 
32'd164685: dataIn1 = 32'd9209
; 
32'd164686: dataIn1 = 32'd9219
; 
32'd164687: dataIn1 = 32'd9220
; 
32'd164688: dataIn1 = 32'd6689
; 
32'd164689: dataIn1 = 32'd6798
; 
32'd164690: dataIn1 = 32'd6799
; 
32'd164691: dataIn1 = 32'd9222
; 
32'd164692: dataIn1 = 32'd9223
; 
32'd164693: dataIn1 = 32'd9225
; 
32'd164694: dataIn1 = 32'd9226
; 
32'd164695: dataIn1 = 32'd6690
; 
32'd164696: dataIn1 = 32'd6800
; 
32'd164697: dataIn1 = 32'd6801
; 
32'd164698: dataIn1 = 32'd9227
; 
32'd164699: dataIn1 = 32'd9229
; 
32'd164700: dataIn1 = 32'd9230
; 
32'd164701: dataIn1 = 32'd9231
; 
32'd164702: dataIn1 = 32'd2324
; 
32'd164703: dataIn1 = 32'd2739
; 
32'd164704: dataIn1 = 32'd2741
; 
32'd164705: dataIn1 = 32'd5323
; 
32'd164706: dataIn1 = 32'd5633
; 
32'd164707: dataIn1 = 32'd6691
; 
32'd164708: dataIn1 = 32'd6692
; 
32'd164709: dataIn1 = 32'd9264
; 
32'd164710: dataIn1 = 32'd9265
; 
32'd164711: dataIn1 = 32'd9311
; 
32'd164712: dataIn1 = 32'd9313
; 
32'd164713: dataIn1 = 32'd9314
; 
32'd164714: dataIn1 = 32'd2102
; 
32'd164715: dataIn1 = 32'd6693
; 
32'd164716: dataIn1 = 32'd9262
; 
32'd164717: dataIn1 = 32'd9263
; 
32'd164718: dataIn1 = 32'd9311
; 
32'd164719: dataIn1 = 32'd9312
; 
32'd164720: dataIn1 = 32'd2104
; 
32'd164721: dataIn1 = 32'd6694
; 
32'd164722: dataIn1 = 32'd9268
; 
32'd164723: dataIn1 = 32'd9269
; 
32'd164724: dataIn1 = 32'd9315
; 
32'd164725: dataIn1 = 32'd9318
; 
32'd164726: dataIn1 = 32'd6695
; 
32'd164727: dataIn1 = 32'd9266
; 
32'd164728: dataIn1 = 32'd9267
; 
32'd164729: dataIn1 = 32'd9315
; 
32'd164730: dataIn1 = 32'd9316
; 
32'd164731: dataIn1 = 32'd9317
; 
32'd164732: dataIn1 = 32'd3920
; 
32'd164733: dataIn1 = 32'd4876
; 
32'd164734: dataIn1 = 32'd5744
; 
32'd164735: dataIn1 = 32'd6050
; 
32'd164736: dataIn1 = 32'd6696
; 
32'd164737: dataIn1 = 32'd6701
; 
32'd164738: dataIn1 = 32'd6732
; 
32'd164739: dataIn1 = 32'd1074
; 
32'd164740: dataIn1 = 32'd4868
; 
32'd164741: dataIn1 = 32'd5910
; 
32'd164742: dataIn1 = 32'd6010
; 
32'd164743: dataIn1 = 32'd6036
; 
32'd164744: dataIn1 = 32'd6697
; 
32'd164745: dataIn1 = 32'd6702
; 
32'd164746: dataIn1 = 32'd2535
; 
32'd164747: dataIn1 = 32'd4610
; 
32'd164748: dataIn1 = 32'd4642
; 
32'd164749: dataIn1 = 32'd4643
; 
32'd164750: dataIn1 = 32'd5952
; 
32'd164751: dataIn1 = 32'd6698
; 
32'd164752: dataIn1 = 32'd2546
; 
32'd164753: dataIn1 = 32'd4635
; 
32'd164754: dataIn1 = 32'd4682
; 
32'd164755: dataIn1 = 32'd4683
; 
32'd164756: dataIn1 = 32'd5982
; 
32'd164757: dataIn1 = 32'd6699
; 
32'd164758: dataIn1 = 32'd447
; 
32'd164759: dataIn1 = 32'd4865
; 
32'd164760: dataIn1 = 32'd4866
; 
32'd164761: dataIn1 = 32'd6006
; 
32'd164762: dataIn1 = 32'd6008
; 
32'd164763: dataIn1 = 32'd6700
; 
32'd164764: dataIn1 = 32'd4866
; 
32'd164765: dataIn1 = 32'd4876
; 
32'd164766: dataIn1 = 32'd6005
; 
32'd164767: dataIn1 = 32'd6048
; 
32'd164768: dataIn1 = 32'd6696
; 
32'd164769: dataIn1 = 32'd6701
; 
32'd164770: dataIn1 = 32'd6732
; 
32'd164771: dataIn1 = 32'd1074
; 
32'd164772: dataIn1 = 32'd4671
; 
32'd164773: dataIn1 = 32'd4867
; 
32'd164774: dataIn1 = 32'd6010
; 
32'd164775: dataIn1 = 32'd6697
; 
32'd164776: dataIn1 = 32'd6702
; 
32'd164777: dataIn1 = 32'd2631
; 
32'd164778: dataIn1 = 32'd4879
; 
32'd164779: dataIn1 = 32'd6045
; 
32'd164780: dataIn1 = 32'd6052
; 
32'd164781: dataIn1 = 32'd6703
; 
32'd164782: dataIn1 = 32'd7257
; 
32'd164783: dataIn1 = 32'd9232
; 
32'd164784: dataIn1 = 32'd2693
; 
32'd164785: dataIn1 = 32'd5116
; 
32'd164786: dataIn1 = 32'd5432
; 
32'd164787: dataIn1 = 32'd6081
; 
32'd164788: dataIn1 = 32'd6704
; 
32'd164789: dataIn1 = 32'd6705
; 
32'd164790: dataIn1 = 32'd6707
; 
32'd164791: dataIn1 = 32'd6734
; 
32'd164792: dataIn1 = 32'd1119
; 
32'd164793: dataIn1 = 32'd5116
; 
32'd164794: dataIn1 = 32'd5432
; 
32'd164795: dataIn1 = 32'd6079
; 
32'd164796: dataIn1 = 32'd6704
; 
32'd164797: dataIn1 = 32'd6705
; 
32'd164798: dataIn1 = 32'd6719
; 
32'd164799: dataIn1 = 32'd6733
; 
32'd164800: dataIn1 = 32'd1120
; 
32'd164801: dataIn1 = 32'd5119
; 
32'd164802: dataIn1 = 32'd5431
; 
32'd164803: dataIn1 = 32'd6096
; 
32'd164804: dataIn1 = 32'd6706
; 
32'd164805: dataIn1 = 32'd6707
; 
32'd164806: dataIn1 = 32'd9262
; 
32'd164807: dataIn1 = 32'd9312
; 
32'd164808: dataIn1 = 32'd2693
; 
32'd164809: dataIn1 = 32'd5119
; 
32'd164810: dataIn1 = 32'd5431
; 
32'd164811: dataIn1 = 32'd6094
; 
32'd164812: dataIn1 = 32'd6704
; 
32'd164813: dataIn1 = 32'd6706
; 
32'd164814: dataIn1 = 32'd6707
; 
32'd164815: dataIn1 = 32'd6734
; 
32'd164816: dataIn1 = 32'd2715
; 
32'd164817: dataIn1 = 32'd5192
; 
32'd164818: dataIn1 = 32'd5438
; 
32'd164819: dataIn1 = 32'd6321
; 
32'd164820: dataIn1 = 32'd6708
; 
32'd164821: dataIn1 = 32'd6709
; 
32'd164822: dataIn1 = 32'd6711
; 
32'd164823: dataIn1 = 32'd6736
; 
32'd164824: dataIn1 = 32'd1127
; 
32'd164825: dataIn1 = 32'd5192
; 
32'd164826: dataIn1 = 32'd5438
; 
32'd164827: dataIn1 = 32'd6319
; 
32'd164828: dataIn1 = 32'd6708
; 
32'd164829: dataIn1 = 32'd6709
; 
32'd164830: dataIn1 = 32'd6726
; 
32'd164831: dataIn1 = 32'd6735
; 
32'd164832: dataIn1 = 32'd1128
; 
32'd164833: dataIn1 = 32'd5195
; 
32'd164834: dataIn1 = 32'd5437
; 
32'd164835: dataIn1 = 32'd6337
; 
32'd164836: dataIn1 = 32'd6710
; 
32'd164837: dataIn1 = 32'd6711
; 
32'd164838: dataIn1 = 32'd6721
; 
32'd164839: dataIn1 = 32'd6737
; 
32'd164840: dataIn1 = 32'd2715
; 
32'd164841: dataIn1 = 32'd5195
; 
32'd164842: dataIn1 = 32'd5437
; 
32'd164843: dataIn1 = 32'd6335
; 
32'd164844: dataIn1 = 32'd6708
; 
32'd164845: dataIn1 = 32'd6710
; 
32'd164846: dataIn1 = 32'd6711
; 
32'd164847: dataIn1 = 32'd6736
; 
32'd164848: dataIn1 = 32'd6712
; 
32'd164849: dataIn1 = 32'd6716
; 
32'd164850: dataIn1 = 32'd6739
; 
32'd164851: dataIn1 = 32'd9748
; 
32'd164852: dataIn1 = 32'd9749
; 
32'd164853: dataIn1 = 32'd9752
; 
32'd164854: dataIn1 = 32'd9776
; 
32'd164855: dataIn1 = 32'd6713
; 
32'd164856: dataIn1 = 32'd10135
; 
32'd164857: dataIn1 = 32'd10137
; 
32'd164858: dataIn1 = 32'd10141
; 
32'd164859: dataIn1 = 32'd10143
; 
32'd164860: dataIn1 = 32'd10149
; 
32'd164861: dataIn1 = 32'd10223
; 
32'd164862: dataIn1 = 32'd5214
; 
32'd164863: dataIn1 = 32'd5215
; 
32'd164864: dataIn1 = 32'd6406
; 
32'd164865: dataIn1 = 32'd6408
; 
32'd164866: dataIn1 = 32'd6714
; 
32'd164867: dataIn1 = 32'd6764
; 
32'd164868: dataIn1 = 32'd8174
; 
32'd164869: dataIn1 = 32'd9233
; 
32'd164870: dataIn1 = 32'd1130
; 
32'd164871: dataIn1 = 32'd5214
; 
32'd164872: dataIn1 = 32'd5439
; 
32'd164873: dataIn1 = 32'd6715
; 
32'd164874: dataIn1 = 32'd6716
; 
32'd164875: dataIn1 = 32'd6723
; 
32'd164876: dataIn1 = 32'd6740
; 
32'd164877: dataIn1 = 32'd9233
; 
32'd164878: dataIn1 = 32'd2720
; 
32'd164879: dataIn1 = 32'd5214
; 
32'd164880: dataIn1 = 32'd5439
; 
32'd164881: dataIn1 = 32'd6409
; 
32'd164882: dataIn1 = 32'd6712
; 
32'd164883: dataIn1 = 32'd6715
; 
32'd164884: dataIn1 = 32'd6716
; 
32'd164885: dataIn1 = 32'd6739
; 
32'd164886: dataIn1 = 32'd9776
; 
32'd164887: dataIn1 = 32'd452
; 
32'd164888: dataIn1 = 32'd2736
; 
32'd164889: dataIn1 = 32'd3980
; 
32'd164890: dataIn1 = 32'd5267
; 
32'd164891: dataIn1 = 32'd6589
; 
32'd164892: dataIn1 = 32'd6717
; 
32'd164893: dataIn1 = 32'd6718
; 
32'd164894: dataIn1 = 32'd6742
; 
32'd164895: dataIn1 = 32'd2734
; 
32'd164896: dataIn1 = 32'd2736
; 
32'd164897: dataIn1 = 32'd5267
; 
32'd164898: dataIn1 = 32'd6588
; 
32'd164899: dataIn1 = 32'd6717
; 
32'd164900: dataIn1 = 32'd6718
; 
32'd164901: dataIn1 = 32'd6720
; 
32'd164902: dataIn1 = 32'd6741
; 
32'd164903: dataIn1 = 32'd1119
; 
32'd164904: dataIn1 = 32'd2735
; 
32'd164905: dataIn1 = 32'd5268
; 
32'd164906: dataIn1 = 32'd6594
; 
32'd164907: dataIn1 = 32'd6705
; 
32'd164908: dataIn1 = 32'd6719
; 
32'd164909: dataIn1 = 32'd6720
; 
32'd164910: dataIn1 = 32'd6733
; 
32'd164911: dataIn1 = 32'd2734
; 
32'd164912: dataIn1 = 32'd2735
; 
32'd164913: dataIn1 = 32'd5268
; 
32'd164914: dataIn1 = 32'd6593
; 
32'd164915: dataIn1 = 32'd6718
; 
32'd164916: dataIn1 = 32'd6719
; 
32'd164917: dataIn1 = 32'd6720
; 
32'd164918: dataIn1 = 32'd6741
; 
32'd164919: dataIn1 = 32'd1128
; 
32'd164920: dataIn1 = 32'd5287
; 
32'd164921: dataIn1 = 32'd5448
; 
32'd164922: dataIn1 = 32'd6637
; 
32'd164923: dataIn1 = 32'd6710
; 
32'd164924: dataIn1 = 32'd6721
; 
32'd164925: dataIn1 = 32'd6722
; 
32'd164926: dataIn1 = 32'd6737
; 
32'd164927: dataIn1 = 32'd2749
; 
32'd164928: dataIn1 = 32'd5287
; 
32'd164929: dataIn1 = 32'd5448
; 
32'd164930: dataIn1 = 32'd6636
; 
32'd164931: dataIn1 = 32'd6721
; 
32'd164932: dataIn1 = 32'd6722
; 
32'd164933: dataIn1 = 32'd9282
; 
32'd164934: dataIn1 = 32'd9323
; 
32'd164935: dataIn1 = 32'd1130
; 
32'd164936: dataIn1 = 32'd5292
; 
32'd164937: dataIn1 = 32'd5450
; 
32'd164938: dataIn1 = 32'd6715
; 
32'd164939: dataIn1 = 32'd6723
; 
32'd164940: dataIn1 = 32'd6724
; 
32'd164941: dataIn1 = 32'd6740
; 
32'd164942: dataIn1 = 32'd9234
; 
32'd164943: dataIn1 = 32'd2750
; 
32'd164944: dataIn1 = 32'd5292
; 
32'd164945: dataIn1 = 32'd5450
; 
32'd164946: dataIn1 = 32'd6654
; 
32'd164947: dataIn1 = 32'd6723
; 
32'd164948: dataIn1 = 32'd6724
; 
32'd164949: dataIn1 = 32'd6727
; 
32'd164950: dataIn1 = 32'd6743
; 
32'd164951: dataIn1 = 32'd5220
; 
32'd164952: dataIn1 = 32'd5292
; 
32'd164953: dataIn1 = 32'd6653
; 
32'd164954: dataIn1 = 32'd6655
; 
32'd164955: dataIn1 = 32'd6725
; 
32'd164956: dataIn1 = 32'd6765
; 
32'd164957: dataIn1 = 32'd9123
; 
32'd164958: dataIn1 = 32'd9234
; 
32'd164959: dataIn1 = 32'd1127
; 
32'd164960: dataIn1 = 32'd5293
; 
32'd164961: dataIn1 = 32'd5449
; 
32'd164962: dataIn1 = 32'd6659
; 
32'd164963: dataIn1 = 32'd6709
; 
32'd164964: dataIn1 = 32'd6726
; 
32'd164965: dataIn1 = 32'd6727
; 
32'd164966: dataIn1 = 32'd6735
; 
32'd164967: dataIn1 = 32'd2750
; 
32'd164968: dataIn1 = 32'd5293
; 
32'd164969: dataIn1 = 32'd5449
; 
32'd164970: dataIn1 = 32'd6657
; 
32'd164971: dataIn1 = 32'd6724
; 
32'd164972: dataIn1 = 32'd6726
; 
32'd164973: dataIn1 = 32'd6727
; 
32'd164974: dataIn1 = 32'd6743
; 
32'd164975: dataIn1 = 32'd5451
; 
32'd164976: dataIn1 = 32'd6728
; 
32'd164977: dataIn1 = 32'd6729
; 
32'd164978: dataIn1 = 32'd10222
; 
32'd164979: dataIn1 = 32'd10223
; 
32'd164980: dataIn1 = 32'd10224
; 
32'd164981: dataIn1 = 32'd10246
; 
32'd164982: dataIn1 = 32'd2751
; 
32'd164983: dataIn1 = 32'd5298
; 
32'd164984: dataIn1 = 32'd5451
; 
32'd164985: dataIn1 = 32'd6677
; 
32'd164986: dataIn1 = 32'd6728
; 
32'd164987: dataIn1 = 32'd6729
; 
32'd164988: dataIn1 = 32'd9284
; 
32'd164989: dataIn1 = 32'd9325
; 
32'd164990: dataIn1 = 32'd10246
; 
32'd164991: dataIn1 = 32'd14
; 
32'd164992: dataIn1 = 32'd2102
; 
32'd164993: dataIn1 = 32'd3457
; 
32'd164994: dataIn1 = 32'd5431
; 
32'd164995: dataIn1 = 32'd6730
; 
32'd164996: dataIn1 = 32'd9312
; 
32'd164997: dataIn1 = 32'd22
; 
32'd164998: dataIn1 = 32'd2104
; 
32'd164999: dataIn1 = 32'd2120
; 
32'd165000: dataIn1 = 32'd5444
; 
32'd165001: dataIn1 = 32'd6731
; 
32'd165002: dataIn1 = 32'd9318
; 
32'd165003: dataIn1 = 32'd447
; 
32'd165004: dataIn1 = 32'd3920
; 
32'd165005: dataIn1 = 32'd4866
; 
32'd165006: dataIn1 = 32'd6696
; 
32'd165007: dataIn1 = 32'd6701
; 
32'd165008: dataIn1 = 32'd6732
; 
32'd165009: dataIn1 = 32'd2735
; 
32'd165010: dataIn1 = 32'd5432
; 
32'd165011: dataIn1 = 32'd5513
; 
32'd165012: dataIn1 = 32'd6705
; 
32'd165013: dataIn1 = 32'd6719
; 
32'd165014: dataIn1 = 32'd6733
; 
32'd165015: dataIn1 = 32'd14
; 
32'd165016: dataIn1 = 32'd5431
; 
32'd165017: dataIn1 = 32'd5432
; 
32'd165018: dataIn1 = 32'd6704
; 
32'd165019: dataIn1 = 32'd6707
; 
32'd165020: dataIn1 = 32'd6734
; 
32'd165021: dataIn1 = 32'd5438
; 
32'd165022: dataIn1 = 32'd5449
; 
32'd165023: dataIn1 = 32'd5518
; 
32'd165024: dataIn1 = 32'd6709
; 
32'd165025: dataIn1 = 32'd6726
; 
32'd165026: dataIn1 = 32'd6735
; 
32'd165027: dataIn1 = 32'd19
; 
32'd165028: dataIn1 = 32'd5437
; 
32'd165029: dataIn1 = 32'd5438
; 
32'd165030: dataIn1 = 32'd6708
; 
32'd165031: dataIn1 = 32'd6711
; 
32'd165032: dataIn1 = 32'd6736
; 
32'd165033: dataIn1 = 32'd5437
; 
32'd165034: dataIn1 = 32'd5448
; 
32'd165035: dataIn1 = 32'd5519
; 
32'd165036: dataIn1 = 32'd6710
; 
32'd165037: dataIn1 = 32'd6721
; 
32'd165038: dataIn1 = 32'd6737
; 
32'd165039: dataIn1 = 32'd5451
; 
32'd165040: dataIn1 = 32'd6738
; 
32'd165041: dataIn1 = 32'd9672
; 
32'd165042: dataIn1 = 32'd9753
; 
32'd165043: dataIn1 = 32'd9754
; 
32'd165044: dataIn1 = 32'd10126
; 
32'd165045: dataIn1 = 32'd10146
; 
32'd165046: dataIn1 = 32'd10224
; 
32'd165047: dataIn1 = 32'd5439
; 
32'd165048: dataIn1 = 32'd5440
; 
32'd165049: dataIn1 = 32'd6712
; 
32'd165050: dataIn1 = 32'd6716
; 
32'd165051: dataIn1 = 32'd6739
; 
32'd165052: dataIn1 = 32'd9675
; 
32'd165053: dataIn1 = 32'd9752
; 
32'd165054: dataIn1 = 32'd9755
; 
32'd165055: dataIn1 = 32'd10131
; 
32'd165056: dataIn1 = 32'd5439
; 
32'd165057: dataIn1 = 32'd5450
; 
32'd165058: dataIn1 = 32'd5521
; 
32'd165059: dataIn1 = 32'd6715
; 
32'd165060: dataIn1 = 32'd6723
; 
32'd165061: dataIn1 = 32'd6740
; 
32'd165062: dataIn1 = 32'd1135
; 
32'd165063: dataIn1 = 32'd2735
; 
32'd165064: dataIn1 = 32'd2736
; 
32'd165065: dataIn1 = 32'd6718
; 
32'd165066: dataIn1 = 32'd6720
; 
32'd165067: dataIn1 = 32'd6741
; 
32'd165068: dataIn1 = 32'd2323
; 
32'd165069: dataIn1 = 32'd2736
; 
32'd165070: dataIn1 = 32'd2737
; 
32'd165071: dataIn1 = 32'd3980
; 
32'd165072: dataIn1 = 32'd6717
; 
32'd165073: dataIn1 = 32'd6742
; 
32'd165074: dataIn1 = 32'd1140
; 
32'd165075: dataIn1 = 32'd5449
; 
32'd165076: dataIn1 = 32'd5450
; 
32'd165077: dataIn1 = 32'd6724
; 
32'd165078: dataIn1 = 32'd6727
; 
32'd165079: dataIn1 = 32'd6743
; 
32'd165080: dataIn1 = 32'd2705
; 
32'd165081: dataIn1 = 32'd5152
; 
32'd165082: dataIn1 = 32'd6190
; 
32'd165083: dataIn1 = 32'd6744
; 
32'd165084: dataIn1 = 32'd6745
; 
32'd165085: dataIn1 = 32'd6748
; 
32'd165086: dataIn1 = 32'd7363
; 
32'd165087: dataIn1 = 32'd9236
; 
32'd165088: dataIn1 = 32'd2705
; 
32'd165089: dataIn1 = 32'd5150
; 
32'd165090: dataIn1 = 32'd6190
; 
32'd165091: dataIn1 = 32'd6744
; 
32'd165092: dataIn1 = 32'd6745
; 
32'd165093: dataIn1 = 32'd6747
; 
32'd165094: dataIn1 = 32'd7360
; 
32'd165095: dataIn1 = 32'd9235
; 
32'd165096: dataIn1 = 32'd5153
; 
32'd165097: dataIn1 = 32'd5154
; 
32'd165098: dataIn1 = 32'd6197
; 
32'd165099: dataIn1 = 32'd6746
; 
32'd165100: dataIn1 = 32'd6747
; 
32'd165101: dataIn1 = 32'd6753
; 
32'd165102: dataIn1 = 32'd7383
; 
32'd165103: dataIn1 = 32'd9237
; 
32'd165104: dataIn1 = 32'd5150
; 
32'd165105: dataIn1 = 32'd5154
; 
32'd165106: dataIn1 = 32'd6197
; 
32'd165107: dataIn1 = 32'd6745
; 
32'd165108: dataIn1 = 32'd6746
; 
32'd165109: dataIn1 = 32'd6747
; 
32'd165110: dataIn1 = 32'd7382
; 
32'd165111: dataIn1 = 32'd9235
; 
32'd165112: dataIn1 = 32'd5152
; 
32'd165113: dataIn1 = 32'd5157
; 
32'd165114: dataIn1 = 32'd6205
; 
32'd165115: dataIn1 = 32'd6744
; 
32'd165116: dataIn1 = 32'd6748
; 
32'd165117: dataIn1 = 32'd6749
; 
32'd165118: dataIn1 = 32'd7418
; 
32'd165119: dataIn1 = 32'd9236
; 
32'd165120: dataIn1 = 32'd5157
; 
32'd165121: dataIn1 = 32'd5158
; 
32'd165122: dataIn1 = 32'd6205
; 
32'd165123: dataIn1 = 32'd6748
; 
32'd165124: dataIn1 = 32'd6749
; 
32'd165125: dataIn1 = 32'd6750
; 
32'd165126: dataIn1 = 32'd7417
; 
32'd165127: dataIn1 = 32'd9238
; 
32'd165128: dataIn1 = 32'd1124
; 
32'd165129: dataIn1 = 32'd5158
; 
32'd165130: dataIn1 = 32'd6226
; 
32'd165131: dataIn1 = 32'd6749
; 
32'd165132: dataIn1 = 32'd6750
; 
32'd165133: dataIn1 = 32'd6751
; 
32'd165134: dataIn1 = 32'd7500
; 
32'd165135: dataIn1 = 32'd9238
; 
32'd165136: dataIn1 = 32'd1124
; 
32'd165137: dataIn1 = 32'd5163
; 
32'd165138: dataIn1 = 32'd6226
; 
32'd165139: dataIn1 = 32'd6750
; 
32'd165140: dataIn1 = 32'd6751
; 
32'd165141: dataIn1 = 32'd7498
; 
32'd165142: dataIn1 = 32'd9280
; 
32'd165143: dataIn1 = 32'd9322
; 
32'd165144: dataIn1 = 32'd1123
; 
32'd165145: dataIn1 = 32'd5167
; 
32'd165146: dataIn1 = 32'd6237
; 
32'd165147: dataIn1 = 32'd6752
; 
32'd165148: dataIn1 = 32'd6753
; 
32'd165149: dataIn1 = 32'd6791
; 
32'd165150: dataIn1 = 32'd7550
; 
32'd165151: dataIn1 = 32'd9239
; 
32'd165152: dataIn1 = 32'd1123
; 
32'd165153: dataIn1 = 32'd5153
; 
32'd165154: dataIn1 = 32'd6237
; 
32'd165155: dataIn1 = 32'd6746
; 
32'd165156: dataIn1 = 32'd6752
; 
32'd165157: dataIn1 = 32'd6753
; 
32'd165158: dataIn1 = 32'd7548
; 
32'd165159: dataIn1 = 32'd9237
; 
32'd165160: dataIn1 = 32'd2710
; 
32'd165161: dataIn1 = 32'd5171
; 
32'd165162: dataIn1 = 32'd6250
; 
32'd165163: dataIn1 = 32'd6754
; 
32'd165164: dataIn1 = 32'd6755
; 
32'd165165: dataIn1 = 32'd6758
; 
32'd165166: dataIn1 = 32'd7614
; 
32'd165167: dataIn1 = 32'd9241
; 
32'd165168: dataIn1 = 32'd2710
; 
32'd165169: dataIn1 = 32'd5169
; 
32'd165170: dataIn1 = 32'd6250
; 
32'd165171: dataIn1 = 32'd6754
; 
32'd165172: dataIn1 = 32'd6755
; 
32'd165173: dataIn1 = 32'd6757
; 
32'd165174: dataIn1 = 32'd7611
; 
32'd165175: dataIn1 = 32'd9240
; 
32'd165176: dataIn1 = 32'd5172
; 
32'd165177: dataIn1 = 32'd5173
; 
32'd165178: dataIn1 = 32'd6257
; 
32'd165179: dataIn1 = 32'd6756
; 
32'd165180: dataIn1 = 32'd6757
; 
32'd165181: dataIn1 = 32'd6763
; 
32'd165182: dataIn1 = 32'd7634
; 
32'd165183: dataIn1 = 32'd9242
; 
32'd165184: dataIn1 = 32'd5169
; 
32'd165185: dataIn1 = 32'd5173
; 
32'd165186: dataIn1 = 32'd6257
; 
32'd165187: dataIn1 = 32'd6755
; 
32'd165188: dataIn1 = 32'd6756
; 
32'd165189: dataIn1 = 32'd6757
; 
32'd165190: dataIn1 = 32'd7633
; 
32'd165191: dataIn1 = 32'd9240
; 
32'd165192: dataIn1 = 32'd5171
; 
32'd165193: dataIn1 = 32'd5176
; 
32'd165194: dataIn1 = 32'd6265
; 
32'd165195: dataIn1 = 32'd6754
; 
32'd165196: dataIn1 = 32'd6758
; 
32'd165197: dataIn1 = 32'd6759
; 
32'd165198: dataIn1 = 32'd7669
; 
32'd165199: dataIn1 = 32'd9241
; 
32'd165200: dataIn1 = 32'd5176
; 
32'd165201: dataIn1 = 32'd5177
; 
32'd165202: dataIn1 = 32'd6265
; 
32'd165203: dataIn1 = 32'd6758
; 
32'd165204: dataIn1 = 32'd6759
; 
32'd165205: dataIn1 = 32'd6760
; 
32'd165206: dataIn1 = 32'd7668
; 
32'd165207: dataIn1 = 32'd9243
; 
32'd165208: dataIn1 = 32'd1126
; 
32'd165209: dataIn1 = 32'd5177
; 
32'd165210: dataIn1 = 32'd6286
; 
32'd165211: dataIn1 = 32'd6759
; 
32'd165212: dataIn1 = 32'd6760
; 
32'd165213: dataIn1 = 32'd6761
; 
32'd165214: dataIn1 = 32'd7753
; 
32'd165215: dataIn1 = 32'd9243
; 
32'd165216: dataIn1 = 32'd1126
; 
32'd165217: dataIn1 = 32'd5182
; 
32'd165218: dataIn1 = 32'd6286
; 
32'd165219: dataIn1 = 32'd6760
; 
32'd165220: dataIn1 = 32'd6761
; 
32'd165221: dataIn1 = 32'd6789
; 
32'd165222: dataIn1 = 32'd7751
; 
32'd165223: dataIn1 = 32'd9244
; 
32'd165224: dataIn1 = 32'd1125
; 
32'd165225: dataIn1 = 32'd5186
; 
32'd165226: dataIn1 = 32'd6297
; 
32'd165227: dataIn1 = 32'd6762
; 
32'd165228: dataIn1 = 32'd6763
; 
32'd165229: dataIn1 = 32'd6793
; 
32'd165230: dataIn1 = 32'd7803
; 
32'd165231: dataIn1 = 32'd9245
; 
32'd165232: dataIn1 = 32'd1125
; 
32'd165233: dataIn1 = 32'd5172
; 
32'd165234: dataIn1 = 32'd6297
; 
32'd165235: dataIn1 = 32'd6756
; 
32'd165236: dataIn1 = 32'd6762
; 
32'd165237: dataIn1 = 32'd6763
; 
32'd165238: dataIn1 = 32'd7801
; 
32'd165239: dataIn1 = 32'd9242
; 
32'd165240: dataIn1 = 32'd1130
; 
32'd165241: dataIn1 = 32'd5215
; 
32'd165242: dataIn1 = 32'd6429
; 
32'd165243: dataIn1 = 32'd6714
; 
32'd165244: dataIn1 = 32'd6764
; 
32'd165245: dataIn1 = 32'd6765
; 
32'd165246: dataIn1 = 32'd8259
; 
32'd165247: dataIn1 = 32'd9233
; 
32'd165248: dataIn1 = 32'd1130
; 
32'd165249: dataIn1 = 32'd5220
; 
32'd165250: dataIn1 = 32'd6429
; 
32'd165251: dataIn1 = 32'd6725
; 
32'd165252: dataIn1 = 32'd6764
; 
32'd165253: dataIn1 = 32'd6765
; 
32'd165254: dataIn1 = 32'd8257
; 
32'd165255: dataIn1 = 32'd9234
; 
32'd165256: dataIn1 = 32'd2725
; 
32'd165257: dataIn1 = 32'd5228
; 
32'd165258: dataIn1 = 32'd6454
; 
32'd165259: dataIn1 = 32'd6766
; 
32'd165260: dataIn1 = 32'd6767
; 
32'd165261: dataIn1 = 32'd6770
; 
32'd165262: dataIn1 = 32'd8372
; 
32'd165263: dataIn1 = 32'd9247
; 
32'd165264: dataIn1 = 32'd2725
; 
32'd165265: dataIn1 = 32'd5226
; 
32'd165266: dataIn1 = 32'd6454
; 
32'd165267: dataIn1 = 32'd6766
; 
32'd165268: dataIn1 = 32'd6767
; 
32'd165269: dataIn1 = 32'd6769
; 
32'd165270: dataIn1 = 32'd8369
; 
32'd165271: dataIn1 = 32'd9246
; 
32'd165272: dataIn1 = 32'd5229
; 
32'd165273: dataIn1 = 32'd5230
; 
32'd165274: dataIn1 = 32'd6461
; 
32'd165275: dataIn1 = 32'd6768
; 
32'd165276: dataIn1 = 32'd6769
; 
32'd165277: dataIn1 = 32'd6775
; 
32'd165278: dataIn1 = 32'd8392
; 
32'd165279: dataIn1 = 32'd9248
; 
32'd165280: dataIn1 = 32'd5226
; 
32'd165281: dataIn1 = 32'd5230
; 
32'd165282: dataIn1 = 32'd6461
; 
32'd165283: dataIn1 = 32'd6767
; 
32'd165284: dataIn1 = 32'd6768
; 
32'd165285: dataIn1 = 32'd6769
; 
32'd165286: dataIn1 = 32'd8391
; 
32'd165287: dataIn1 = 32'd9246
; 
32'd165288: dataIn1 = 32'd5228
; 
32'd165289: dataIn1 = 32'd5233
; 
32'd165290: dataIn1 = 32'd6469
; 
32'd165291: dataIn1 = 32'd6766
; 
32'd165292: dataIn1 = 32'd6770
; 
32'd165293: dataIn1 = 32'd6771
; 
32'd165294: dataIn1 = 32'd8427
; 
32'd165295: dataIn1 = 32'd9247
; 
32'd165296: dataIn1 = 32'd5233
; 
32'd165297: dataIn1 = 32'd5234
; 
32'd165298: dataIn1 = 32'd6469
; 
32'd165299: dataIn1 = 32'd6770
; 
32'd165300: dataIn1 = 32'd6771
; 
32'd165301: dataIn1 = 32'd6772
; 
32'd165302: dataIn1 = 32'd8426
; 
32'd165303: dataIn1 = 32'd9249
; 
32'd165304: dataIn1 = 32'd1132
; 
32'd165305: dataIn1 = 32'd5234
; 
32'd165306: dataIn1 = 32'd6490
; 
32'd165307: dataIn1 = 32'd6771
; 
32'd165308: dataIn1 = 32'd6772
; 
32'd165309: dataIn1 = 32'd6773
; 
32'd165310: dataIn1 = 32'd8511
; 
32'd165311: dataIn1 = 32'd9249
; 
32'd165312: dataIn1 = 32'd1132
; 
32'd165313: dataIn1 = 32'd5239
; 
32'd165314: dataIn1 = 32'd6490
; 
32'd165315: dataIn1 = 32'd6772
; 
32'd165316: dataIn1 = 32'd6773
; 
32'd165317: dataIn1 = 32'd6795
; 
32'd165318: dataIn1 = 32'd8509
; 
32'd165319: dataIn1 = 32'd9250
; 
32'd165320: dataIn1 = 32'd1131
; 
32'd165321: dataIn1 = 32'd5243
; 
32'd165322: dataIn1 = 32'd6501
; 
32'd165323: dataIn1 = 32'd6774
; 
32'd165324: dataIn1 = 32'd6775
; 
32'd165325: dataIn1 = 32'd6801
; 
32'd165326: dataIn1 = 32'd8561
; 
32'd165327: dataIn1 = 32'd9251
; 
32'd165328: dataIn1 = 32'd1131
; 
32'd165329: dataIn1 = 32'd5229
; 
32'd165330: dataIn1 = 32'd6501
; 
32'd165331: dataIn1 = 32'd6768
; 
32'd165332: dataIn1 = 32'd6774
; 
32'd165333: dataIn1 = 32'd6775
; 
32'd165334: dataIn1 = 32'd8559
; 
32'd165335: dataIn1 = 32'd9248
; 
32'd165336: dataIn1 = 32'd2730
; 
32'd165337: dataIn1 = 32'd5247
; 
32'd165338: dataIn1 = 32'd6514
; 
32'd165339: dataIn1 = 32'd6776
; 
32'd165340: dataIn1 = 32'd6777
; 
32'd165341: dataIn1 = 32'd6780
; 
32'd165342: dataIn1 = 32'd8625
; 
32'd165343: dataIn1 = 32'd9253
; 
32'd165344: dataIn1 = 32'd2730
; 
32'd165345: dataIn1 = 32'd5245
; 
32'd165346: dataIn1 = 32'd6514
; 
32'd165347: dataIn1 = 32'd6776
; 
32'd165348: dataIn1 = 32'd6777
; 
32'd165349: dataIn1 = 32'd6779
; 
32'd165350: dataIn1 = 32'd8622
; 
32'd165351: dataIn1 = 32'd9252
; 
32'd165352: dataIn1 = 32'd5248
; 
32'd165353: dataIn1 = 32'd5249
; 
32'd165354: dataIn1 = 32'd6521
; 
32'd165355: dataIn1 = 32'd6778
; 
32'd165356: dataIn1 = 32'd6779
; 
32'd165357: dataIn1 = 32'd6785
; 
32'd165358: dataIn1 = 32'd8645
; 
32'd165359: dataIn1 = 32'd9254
; 
32'd165360: dataIn1 = 32'd5245
; 
32'd165361: dataIn1 = 32'd5249
; 
32'd165362: dataIn1 = 32'd6521
; 
32'd165363: dataIn1 = 32'd6777
; 
32'd165364: dataIn1 = 32'd6778
; 
32'd165365: dataIn1 = 32'd6779
; 
32'd165366: dataIn1 = 32'd8644
; 
32'd165367: dataIn1 = 32'd9252
; 
32'd165368: dataIn1 = 32'd5247
; 
32'd165369: dataIn1 = 32'd5252
; 
32'd165370: dataIn1 = 32'd6529
; 
32'd165371: dataIn1 = 32'd6776
; 
32'd165372: dataIn1 = 32'd6780
; 
32'd165373: dataIn1 = 32'd6781
; 
32'd165374: dataIn1 = 32'd8680
; 
32'd165375: dataIn1 = 32'd9253
; 
32'd165376: dataIn1 = 32'd5252
; 
32'd165377: dataIn1 = 32'd5253
; 
32'd165378: dataIn1 = 32'd6529
; 
32'd165379: dataIn1 = 32'd6780
; 
32'd165380: dataIn1 = 32'd6781
; 
32'd165381: dataIn1 = 32'd6782
; 
32'd165382: dataIn1 = 32'd8679
; 
32'd165383: dataIn1 = 32'd9255
; 
32'd165384: dataIn1 = 32'd1134
; 
32'd165385: dataIn1 = 32'd5253
; 
32'd165386: dataIn1 = 32'd6550
; 
32'd165387: dataIn1 = 32'd6781
; 
32'd165388: dataIn1 = 32'd6782
; 
32'd165389: dataIn1 = 32'd6783
; 
32'd165390: dataIn1 = 32'd8764
; 
32'd165391: dataIn1 = 32'd9255
; 
32'd165392: dataIn1 = 32'd1134
; 
32'd165393: dataIn1 = 32'd5258
; 
32'd165394: dataIn1 = 32'd6550
; 
32'd165395: dataIn1 = 32'd6782
; 
32'd165396: dataIn1 = 32'd6783
; 
32'd165397: dataIn1 = 32'd6799
; 
32'd165398: dataIn1 = 32'd8762
; 
32'd165399: dataIn1 = 32'd9256
; 
32'd165400: dataIn1 = 32'd1133
; 
32'd165401: dataIn1 = 32'd5262
; 
32'd165402: dataIn1 = 32'd6561
; 
32'd165403: dataIn1 = 32'd6784
; 
32'd165404: dataIn1 = 32'd6785
; 
32'd165405: dataIn1 = 32'd6849
; 
32'd165406: dataIn1 = 32'd8814
; 
32'd165407: dataIn1 = 32'd9257
; 
32'd165408: dataIn1 = 32'd1133
; 
32'd165409: dataIn1 = 32'd5248
; 
32'd165410: dataIn1 = 32'd6561
; 
32'd165411: dataIn1 = 32'd6778
; 
32'd165412: dataIn1 = 32'd6784
; 
32'd165413: dataIn1 = 32'd6785
; 
32'd165414: dataIn1 = 32'd8812
; 
32'd165415: dataIn1 = 32'd9254
; 
32'd165416: dataIn1 = 32'd2747
; 
32'd165417: dataIn1 = 32'd5281
; 
32'd165418: dataIn1 = 32'd6611
; 
32'd165419: dataIn1 = 32'd6786
; 
32'd165420: dataIn1 = 32'd6787
; 
32'd165421: dataIn1 = 32'd6790
; 
32'd165422: dataIn1 = 32'd8984
; 
32'd165423: dataIn1 = 32'd9259
; 
32'd165424: dataIn1 = 32'd2747
; 
32'd165425: dataIn1 = 32'd5280
; 
32'd165426: dataIn1 = 32'd6611
; 
32'd165427: dataIn1 = 32'd6786
; 
32'd165428: dataIn1 = 32'd6787
; 
32'd165429: dataIn1 = 32'd6788
; 
32'd165430: dataIn1 = 32'd8982
; 
32'd165431: dataIn1 = 32'd9258
; 
32'd165432: dataIn1 = 32'd5280
; 
32'd165433: dataIn1 = 32'd5282
; 
32'd165434: dataIn1 = 32'd6621
; 
32'd165435: dataIn1 = 32'd6787
; 
32'd165436: dataIn1 = 32'd6788
; 
32'd165437: dataIn1 = 32'd6789
; 
32'd165438: dataIn1 = 32'd9021
; 
32'd165439: dataIn1 = 32'd9258
; 
32'd165440: dataIn1 = 32'd5182
; 
32'd165441: dataIn1 = 32'd5282
; 
32'd165442: dataIn1 = 32'd6621
; 
32'd165443: dataIn1 = 32'd6761
; 
32'd165444: dataIn1 = 32'd6788
; 
32'd165445: dataIn1 = 32'd6789
; 
32'd165446: dataIn1 = 32'd9020
; 
32'd165447: dataIn1 = 32'd9244
; 
32'd165448: dataIn1 = 32'd5281
; 
32'd165449: dataIn1 = 32'd5283
; 
32'd165450: dataIn1 = 32'd6622
; 
32'd165451: dataIn1 = 32'd6786
; 
32'd165452: dataIn1 = 32'd6790
; 
32'd165453: dataIn1 = 32'd6791
; 
32'd165454: dataIn1 = 32'd9026
; 
32'd165455: dataIn1 = 32'd9259
; 
32'd165456: dataIn1 = 32'd5167
; 
32'd165457: dataIn1 = 32'd5283
; 
32'd165458: dataIn1 = 32'd6622
; 
32'd165459: dataIn1 = 32'd6752
; 
32'd165460: dataIn1 = 32'd6790
; 
32'd165461: dataIn1 = 32'd6791
; 
32'd165462: dataIn1 = 32'd9025
; 
32'd165463: dataIn1 = 32'd9239
; 
32'd165464: dataIn1 = 32'd5286
; 
32'd165465: dataIn1 = 32'd5288
; 
32'd165466: dataIn1 = 32'd6626
; 
32'd165467: dataIn1 = 32'd6640
; 
32'd165468: dataIn1 = 32'd6792
; 
32'd165469: dataIn1 = 32'd6793
; 
32'd165470: dataIn1 = 32'd9036
; 
32'd165471: dataIn1 = 32'd9078
; 
32'd165472: dataIn1 = 32'd5186
; 
32'd165473: dataIn1 = 32'd5288
; 
32'd165474: dataIn1 = 32'd6640
; 
32'd165475: dataIn1 = 32'd6762
; 
32'd165476: dataIn1 = 32'd6792
; 
32'd165477: dataIn1 = 32'd6793
; 
32'd165478: dataIn1 = 32'd9077
; 
32'd165479: dataIn1 = 32'd9245
; 
32'd165480: dataIn1 = 32'd5295
; 
32'd165481: dataIn1 = 32'd5297
; 
32'd165482: dataIn1 = 32'd6665
; 
32'd165483: dataIn1 = 32'd6673
; 
32'd165484: dataIn1 = 32'd6794
; 
32'd165485: dataIn1 = 32'd6795
; 
32'd165486: dataIn1 = 32'd9139
; 
32'd165487: dataIn1 = 32'd9176
; 
32'd165488: dataIn1 = 32'd5239
; 
32'd165489: dataIn1 = 32'd5297
; 
32'd165490: dataIn1 = 32'd6673
; 
32'd165491: dataIn1 = 32'd6773
; 
32'd165492: dataIn1 = 32'd6794
; 
32'd165493: dataIn1 = 32'd6795
; 
32'd165494: dataIn1 = 32'd9175
; 
32'd165495: dataIn1 = 32'd9250
; 
32'd165496: dataIn1 = 32'd2752
; 
32'd165497: dataIn1 = 32'd5301
; 
32'd165498: dataIn1 = 32'd6679
; 
32'd165499: dataIn1 = 32'd6796
; 
32'd165500: dataIn1 = 32'd6797
; 
32'd165501: dataIn1 = 32'd6800
; 
32'd165502: dataIn1 = 32'd9189
; 
32'd165503: dataIn1 = 32'd9261
; 
32'd165504: dataIn1 = 32'd2752
; 
32'd165505: dataIn1 = 32'd5300
; 
32'd165506: dataIn1 = 32'd6679
; 
32'd165507: dataIn1 = 32'd6796
; 
32'd165508: dataIn1 = 32'd6797
; 
32'd165509: dataIn1 = 32'd6798
; 
32'd165510: dataIn1 = 32'd9187
; 
32'd165511: dataIn1 = 32'd9260
; 
32'd165512: dataIn1 = 32'd5300
; 
32'd165513: dataIn1 = 32'd5302
; 
32'd165514: dataIn1 = 32'd6689
; 
32'd165515: dataIn1 = 32'd6797
; 
32'd165516: dataIn1 = 32'd6798
; 
32'd165517: dataIn1 = 32'd6799
; 
32'd165518: dataIn1 = 32'd9226
; 
32'd165519: dataIn1 = 32'd9260
; 
32'd165520: dataIn1 = 32'd5258
; 
32'd165521: dataIn1 = 32'd5302
; 
32'd165522: dataIn1 = 32'd6689
; 
32'd165523: dataIn1 = 32'd6783
; 
32'd165524: dataIn1 = 32'd6798
; 
32'd165525: dataIn1 = 32'd6799
; 
32'd165526: dataIn1 = 32'd9225
; 
32'd165527: dataIn1 = 32'd9256
; 
32'd165528: dataIn1 = 32'd5301
; 
32'd165529: dataIn1 = 32'd5303
; 
32'd165530: dataIn1 = 32'd6690
; 
32'd165531: dataIn1 = 32'd6796
; 
32'd165532: dataIn1 = 32'd6800
; 
32'd165533: dataIn1 = 32'd6801
; 
32'd165534: dataIn1 = 32'd9231
; 
32'd165535: dataIn1 = 32'd9261
; 
32'd165536: dataIn1 = 32'd5243
; 
32'd165537: dataIn1 = 32'd5303
; 
32'd165538: dataIn1 = 32'd6690
; 
32'd165539: dataIn1 = 32'd6774
; 
32'd165540: dataIn1 = 32'd6800
; 
32'd165541: dataIn1 = 32'd6801
; 
32'd165542: dataIn1 = 32'd9230
; 
32'd165543: dataIn1 = 32'd9251
; 
32'd165544: dataIn1 = 32'd6802
; 
32'd165545: dataIn1 = 32'd6805
; 
32'd165546: dataIn1 = 32'd9341
; 
32'd165547: dataIn1 = 32'd9342
; 
32'd165548: dataIn1 = 32'd9346
; 
32'd165549: dataIn1 = 32'd9348
; 
32'd165550: dataIn1 = 32'd6803
; 
32'd165551: dataIn1 = 32'd9340
; 
32'd165552: dataIn1 = 32'd9342
; 
32'd165553: dataIn1 = 32'd9344
; 
32'd165554: dataIn1 = 32'd9347
; 
32'd165555: dataIn1 = 32'd9349
; 
32'd165556: dataIn1 = 32'd9351
; 
32'd165557: dataIn1 = 32'd6804
; 
32'd165558: dataIn1 = 32'd9340
; 
32'd165559: dataIn1 = 32'd9341
; 
32'd165560: dataIn1 = 32'd9343
; 
32'd165561: dataIn1 = 32'd9345
; 
32'd165562: dataIn1 = 32'd9356
; 
32'd165563: dataIn1 = 32'd9357
; 
32'd165564: dataIn1 = 32'd3583
; 
32'd165565: dataIn1 = 32'd6802
; 
32'd165566: dataIn1 = 32'd6805
; 
32'd165567: dataIn1 = 32'd6806
; 
32'd165568: dataIn1 = 32'd6821
; 
32'd165569: dataIn1 = 32'd6824
; 
32'd165570: dataIn1 = 32'd9346
; 
32'd165571: dataIn1 = 32'd9348
; 
32'd165572: dataIn1 = 32'd3583
; 
32'd165573: dataIn1 = 32'd5636
; 
32'd165574: dataIn1 = 32'd6805
; 
32'd165575: dataIn1 = 32'd6806
; 
32'd165576: dataIn1 = 32'd6816
; 
32'd165577: dataIn1 = 32'd6819
; 
32'd165578: dataIn1 = 32'd9346
; 
32'd165579: dataIn1 = 32'd9383
; 
32'd165580: dataIn1 = 32'd6807
; 
32'd165581: dataIn1 = 32'd9350
; 
32'd165582: dataIn1 = 32'd9351
; 
32'd165583: dataIn1 = 32'd9354
; 
32'd165584: dataIn1 = 32'd9355
; 
32'd165585: dataIn1 = 32'd9385
; 
32'd165586: dataIn1 = 32'd9386
; 
32'd165587: dataIn1 = 32'd6808
; 
32'd165588: dataIn1 = 32'd9349
; 
32'd165589: dataIn1 = 32'd9350
; 
32'd165590: dataIn1 = 32'd9352
; 
32'd165591: dataIn1 = 32'd9353
; 
32'd165592: dataIn1 = 32'd9372
; 
32'd165593: dataIn1 = 32'd9373
; 
32'd165594: dataIn1 = 32'd6809
; 
32'd165595: dataIn1 = 32'd9357
; 
32'd165596: dataIn1 = 32'd9358
; 
32'd165597: dataIn1 = 32'd9360
; 
32'd165598: dataIn1 = 32'd9362
; 
32'd165599: dataIn1 = 32'd9381
; 
32'd165600: dataIn1 = 32'd9382
; 
32'd165601: dataIn1 = 32'd6810
; 
32'd165602: dataIn1 = 32'd9356
; 
32'd165603: dataIn1 = 32'd9358
; 
32'd165604: dataIn1 = 32'd9359
; 
32'd165605: dataIn1 = 32'd9361
; 
32'd165606: dataIn1 = 32'd9377
; 
32'd165607: dataIn1 = 32'd9379
; 
32'd165608: dataIn1 = 32'd6811
; 
32'd165609: dataIn1 = 32'd9364
; 
32'd165610: dataIn1 = 32'd9365
; 
32'd165611: dataIn1 = 32'd9369
; 
32'd165612: dataIn1 = 32'd9371
; 
32'd165613: dataIn1 = 32'd9808
; 
32'd165614: dataIn1 = 32'd9809
; 
32'd165615: dataIn1 = 32'd6812
; 
32'd165616: dataIn1 = 32'd9363
; 
32'd165617: dataIn1 = 32'd9365
; 
32'd165618: dataIn1 = 32'd9367
; 
32'd165619: dataIn1 = 32'd9370
; 
32'd165620: dataIn1 = 32'd9372
; 
32'd165621: dataIn1 = 32'd9374
; 
32'd165622: dataIn1 = 32'd6813
; 
32'd165623: dataIn1 = 32'd9363
; 
32'd165624: dataIn1 = 32'd9364
; 
32'd165625: dataIn1 = 32'd9366
; 
32'd165626: dataIn1 = 32'd9368
; 
32'd165627: dataIn1 = 32'd9377
; 
32'd165628: dataIn1 = 32'd9378
; 
32'd165629: dataIn1 = 32'd6814
; 
32'd165630: dataIn1 = 32'd9756
; 
32'd165631: dataIn1 = 32'd9757
; 
32'd165632: dataIn1 = 32'd9809
; 
32'd165633: dataIn1 = 32'd9810
; 
32'd165634: dataIn1 = 32'd6815
; 
32'd165635: dataIn1 = 32'd9373
; 
32'd165636: dataIn1 = 32'd9374
; 
32'd165637: dataIn1 = 32'd9375
; 
32'd165638: dataIn1 = 32'd9376
; 
32'd165639: dataIn1 = 32'd5639
; 
32'd165640: dataIn1 = 32'd6806
; 
32'd165641: dataIn1 = 32'd6816
; 
32'd165642: dataIn1 = 32'd6817
; 
32'd165643: dataIn1 = 32'd6818
; 
32'd165644: dataIn1 = 32'd6819
; 
32'd165645: dataIn1 = 32'd9383
; 
32'd165646: dataIn1 = 32'd9446
; 
32'd165647: dataIn1 = 32'd5125
; 
32'd165648: dataIn1 = 32'd5639
; 
32'd165649: dataIn1 = 32'd6118
; 
32'd165650: dataIn1 = 32'd6816
; 
32'd165651: dataIn1 = 32'd6817
; 
32'd165652: dataIn1 = 32'd6820
; 
32'd165653: dataIn1 = 32'd9446
; 
32'd165654: dataIn1 = 32'd6816
; 
32'd165655: dataIn1 = 32'd6818
; 
32'd165656: dataIn1 = 32'd9380
; 
32'd165657: dataIn1 = 32'd9381
; 
32'd165658: dataIn1 = 32'd9383
; 
32'd165659: dataIn1 = 32'd9446
; 
32'd165660: dataIn1 = 32'd3583
; 
32'd165661: dataIn1 = 32'd5639
; 
32'd165662: dataIn1 = 32'd6806
; 
32'd165663: dataIn1 = 32'd6816
; 
32'd165664: dataIn1 = 32'd6819
; 
32'd165665: dataIn1 = 32'd9263
; 
32'd165666: dataIn1 = 32'd9265
; 
32'd165667: dataIn1 = 32'd1120
; 
32'd165668: dataIn1 = 32'd5639
; 
32'd165669: dataIn1 = 32'd6118
; 
32'd165670: dataIn1 = 32'd6817
; 
32'd165671: dataIn1 = 32'd6820
; 
32'd165672: dataIn1 = 32'd9262
; 
32'd165673: dataIn1 = 32'd9263
; 
32'd165674: dataIn1 = 32'd5637
; 
32'd165675: dataIn1 = 32'd5641
; 
32'd165676: dataIn1 = 32'd6805
; 
32'd165677: dataIn1 = 32'd6821
; 
32'd165678: dataIn1 = 32'd6823
; 
32'd165679: dataIn1 = 32'd6824
; 
32'd165680: dataIn1 = 32'd9348
; 
32'd165681: dataIn1 = 32'd9390
; 
32'd165682: dataIn1 = 32'd6822
; 
32'd165683: dataIn1 = 32'd6823
; 
32'd165684: dataIn1 = 32'd9384
; 
32'd165685: dataIn1 = 32'd9386
; 
32'd165686: dataIn1 = 32'd9388
; 
32'd165687: dataIn1 = 32'd9390
; 
32'd165688: dataIn1 = 32'd5641
; 
32'd165689: dataIn1 = 32'd6821
; 
32'd165690: dataIn1 = 32'd6822
; 
32'd165691: dataIn1 = 32'd6823
; 
32'd165692: dataIn1 = 32'd6826
; 
32'd165693: dataIn1 = 32'd6827
; 
32'd165694: dataIn1 = 32'd9388
; 
32'd165695: dataIn1 = 32'd9390
; 
32'd165696: dataIn1 = 32'd3583
; 
32'd165697: dataIn1 = 32'd5641
; 
32'd165698: dataIn1 = 32'd6805
; 
32'd165699: dataIn1 = 32'd6821
; 
32'd165700: dataIn1 = 32'd6824
; 
32'd165701: dataIn1 = 32'd9264
; 
32'd165702: dataIn1 = 32'd9265
; 
32'd165703: dataIn1 = 32'd6825
; 
32'd165704: dataIn1 = 32'd9384
; 
32'd165705: dataIn1 = 32'd9385
; 
32'd165706: dataIn1 = 32'd9387
; 
32'd165707: dataIn1 = 32'd9389
; 
32'd165708: dataIn1 = 32'd2103
; 
32'd165709: dataIn1 = 32'd5641
; 
32'd165710: dataIn1 = 32'd6823
; 
32'd165711: dataIn1 = 32'd6826
; 
32'd165712: dataIn1 = 32'd6827
; 
32'd165713: dataIn1 = 32'd9264
; 
32'd165714: dataIn1 = 32'd10286
; 
32'd165715: dataIn1 = 32'd2103
; 
32'd165716: dataIn1 = 32'd5640
; 
32'd165717: dataIn1 = 32'd6823
; 
32'd165718: dataIn1 = 32'd6826
; 
32'd165719: dataIn1 = 32'd6827
; 
32'd165720: dataIn1 = 32'd9388
; 
32'd165721: dataIn1 = 32'd6828
; 
32'd165722: dataIn1 = 32'd6832
; 
32'd165723: dataIn1 = 32'd9392
; 
32'd165724: dataIn1 = 32'd9393
; 
32'd165725: dataIn1 = 32'd9397
; 
32'd165726: dataIn1 = 32'd9399
; 
32'd165727: dataIn1 = 32'd6829
; 
32'd165728: dataIn1 = 32'd9391
; 
32'd165729: dataIn1 = 32'd9393
; 
32'd165730: dataIn1 = 32'd9395
; 
32'd165731: dataIn1 = 32'd9398
; 
32'd165732: dataIn1 = 32'd9400
; 
32'd165733: dataIn1 = 32'd9402
; 
32'd165734: dataIn1 = 32'd6830
; 
32'd165735: dataIn1 = 32'd9391
; 
32'd165736: dataIn1 = 32'd9392
; 
32'd165737: dataIn1 = 32'd9394
; 
32'd165738: dataIn1 = 32'd9396
; 
32'd165739: dataIn1 = 32'd9407
; 
32'd165740: dataIn1 = 32'd9408
; 
32'd165741: dataIn1 = 32'd3585
; 
32'd165742: dataIn1 = 32'd5644
; 
32'd165743: dataIn1 = 32'd6831
; 
32'd165744: dataIn1 = 32'd6832
; 
32'd165745: dataIn1 = 32'd6847
; 
32'd165746: dataIn1 = 32'd6850
; 
32'd165747: dataIn1 = 32'd9399
; 
32'd165748: dataIn1 = 32'd9445
; 
32'd165749: dataIn1 = 32'd3585
; 
32'd165750: dataIn1 = 32'd6828
; 
32'd165751: dataIn1 = 32'd6831
; 
32'd165752: dataIn1 = 32'd6832
; 
32'd165753: dataIn1 = 32'd6842
; 
32'd165754: dataIn1 = 32'd6845
; 
32'd165755: dataIn1 = 32'd9397
; 
32'd165756: dataIn1 = 32'd9399
; 
32'd165757: dataIn1 = 32'd6833
; 
32'd165758: dataIn1 = 32'd9401
; 
32'd165759: dataIn1 = 32'd9402
; 
32'd165760: dataIn1 = 32'd9405
; 
32'd165761: dataIn1 = 32'd9406
; 
32'd165762: dataIn1 = 32'd9443
; 
32'd165763: dataIn1 = 32'd9444
; 
32'd165764: dataIn1 = 32'd6834
; 
32'd165765: dataIn1 = 32'd9400
; 
32'd165766: dataIn1 = 32'd9401
; 
32'd165767: dataIn1 = 32'd9403
; 
32'd165768: dataIn1 = 32'd9404
; 
32'd165769: dataIn1 = 32'd9427
; 
32'd165770: dataIn1 = 32'd9428
; 
32'd165771: dataIn1 = 32'd6835
; 
32'd165772: dataIn1 = 32'd9408
; 
32'd165773: dataIn1 = 32'd9409
; 
32'd165774: dataIn1 = 32'd9411
; 
32'd165775: dataIn1 = 32'd9413
; 
32'd165776: dataIn1 = 32'd9436
; 
32'd165777: dataIn1 = 32'd9437
; 
32'd165778: dataIn1 = 32'd6836
; 
32'd165779: dataIn1 = 32'd9407
; 
32'd165780: dataIn1 = 32'd9409
; 
32'd165781: dataIn1 = 32'd9410
; 
32'd165782: dataIn1 = 32'd9412
; 
32'd165783: dataIn1 = 32'd9430
; 
32'd165784: dataIn1 = 32'd9432
; 
32'd165785: dataIn1 = 32'd6837
; 
32'd165786: dataIn1 = 32'd9415
; 
32'd165787: dataIn1 = 32'd9416
; 
32'd165788: dataIn1 = 32'd9420
; 
32'd165789: dataIn1 = 32'd9422
; 
32'd165790: dataIn1 = 32'd9424
; 
32'd165791: dataIn1 = 32'd9425
; 
32'd165792: dataIn1 = 32'd6838
; 
32'd165793: dataIn1 = 32'd9414
; 
32'd165794: dataIn1 = 32'd9416
; 
32'd165795: dataIn1 = 32'd9418
; 
32'd165796: dataIn1 = 32'd9421
; 
32'd165797: dataIn1 = 32'd9427
; 
32'd165798: dataIn1 = 32'd9429
; 
32'd165799: dataIn1 = 32'd6839
; 
32'd165800: dataIn1 = 32'd9414
; 
32'd165801: dataIn1 = 32'd9415
; 
32'd165802: dataIn1 = 32'd9417
; 
32'd165803: dataIn1 = 32'd9419
; 
32'd165804: dataIn1 = 32'd9430
; 
32'd165805: dataIn1 = 32'd9431
; 
32'd165806: dataIn1 = 32'd6840
; 
32'd165807: dataIn1 = 32'd9423
; 
32'd165808: dataIn1 = 32'd9424
; 
32'd165809: dataIn1 = 32'd9426
; 
32'd165810: dataIn1 = 32'd9448
; 
32'd165811: dataIn1 = 32'd6841
; 
32'd165812: dataIn1 = 32'd9431
; 
32'd165813: dataIn1 = 32'd9432
; 
32'd165814: dataIn1 = 32'd9433
; 
32'd165815: dataIn1 = 32'd9434
; 
32'd165816: dataIn1 = 32'd5643
; 
32'd165817: dataIn1 = 32'd5647
; 
32'd165818: dataIn1 = 32'd6832
; 
32'd165819: dataIn1 = 32'd6842
; 
32'd165820: dataIn1 = 32'd6843
; 
32'd165821: dataIn1 = 32'd6845
; 
32'd165822: dataIn1 = 32'd9397
; 
32'd165823: dataIn1 = 32'd9440
; 
32'd165824: dataIn1 = 32'd2105
; 
32'd165825: dataIn1 = 32'd5647
; 
32'd165826: dataIn1 = 32'd6842
; 
32'd165827: dataIn1 = 32'd6843
; 
32'd165828: dataIn1 = 32'd6844
; 
32'd165829: dataIn1 = 32'd9438
; 
32'd165830: dataIn1 = 32'd9440
; 
32'd165831: dataIn1 = 32'd10291
; 
32'd165832: dataIn1 = 32'd6843
; 
32'd165833: dataIn1 = 32'd6844
; 
32'd165834: dataIn1 = 32'd9435
; 
32'd165835: dataIn1 = 32'd9436
; 
32'd165836: dataIn1 = 32'd9438
; 
32'd165837: dataIn1 = 32'd9440
; 
32'd165838: dataIn1 = 32'd3585
; 
32'd165839: dataIn1 = 32'd5647
; 
32'd165840: dataIn1 = 32'd6832
; 
32'd165841: dataIn1 = 32'd6842
; 
32'd165842: dataIn1 = 32'd6845
; 
32'd165843: dataIn1 = 32'd9266
; 
32'd165844: dataIn1 = 32'd9267
; 
32'd165845: dataIn1 = 32'd6846
; 
32'd165846: dataIn1 = 32'd9435
; 
32'd165847: dataIn1 = 32'd9437
; 
32'd165848: dataIn1 = 32'd9439
; 
32'd165849: dataIn1 = 32'd9441
; 
32'd165850: dataIn1 = 32'd5648
; 
32'd165851: dataIn1 = 32'd6831
; 
32'd165852: dataIn1 = 32'd6847
; 
32'd165853: dataIn1 = 32'd6848
; 
32'd165854: dataIn1 = 32'd6849
; 
32'd165855: dataIn1 = 32'd6850
; 
32'd165856: dataIn1 = 32'd9445
; 
32'd165857: dataIn1 = 32'd9447
; 
32'd165858: dataIn1 = 32'd6847
; 
32'd165859: dataIn1 = 32'd6848
; 
32'd165860: dataIn1 = 32'd9442
; 
32'd165861: dataIn1 = 32'd9444
; 
32'd165862: dataIn1 = 32'd9445
; 
32'd165863: dataIn1 = 32'd9447
; 
32'd165864: dataIn1 = 32'd5262
; 
32'd165865: dataIn1 = 32'd5648
; 
32'd165866: dataIn1 = 32'd6784
; 
32'd165867: dataIn1 = 32'd6847
; 
32'd165868: dataIn1 = 32'd6849
; 
32'd165869: dataIn1 = 32'd9257
; 
32'd165870: dataIn1 = 32'd9447
; 
32'd165871: dataIn1 = 32'd3585
; 
32'd165872: dataIn1 = 32'd5648
; 
32'd165873: dataIn1 = 32'd6831
; 
32'd165874: dataIn1 = 32'd6847
; 
32'd165875: dataIn1 = 32'd6850
; 
32'd165876: dataIn1 = 32'd9267
; 
32'd165877: dataIn1 = 32'd9269
; 
32'd165878: dataIn1 = 32'd5828
; 
32'd165879: dataIn1 = 32'd5829
; 
32'd165880: dataIn1 = 32'd6851
; 
32'd165881: dataIn1 = 32'd6852
; 
32'd165882: dataIn1 = 32'd6853
; 
32'd165883: dataIn1 = 32'd6854
; 
32'd165884: dataIn1 = 32'd6855
; 
32'd165885: dataIn1 = 32'd5827
; 
32'd165886: dataIn1 = 32'd5829
; 
32'd165887: dataIn1 = 32'd6851
; 
32'd165888: dataIn1 = 32'd6852
; 
32'd165889: dataIn1 = 32'd6853
; 
32'd165890: dataIn1 = 32'd6856
; 
32'd165891: dataIn1 = 32'd6857
; 
32'd165892: dataIn1 = 32'd5827
; 
32'd165893: dataIn1 = 32'd5828
; 
32'd165894: dataIn1 = 32'd6851
; 
32'd165895: dataIn1 = 32'd6852
; 
32'd165896: dataIn1 = 32'd6853
; 
32'd165897: dataIn1 = 32'd6858
; 
32'd165898: dataIn1 = 32'd6859
; 
32'd165899: dataIn1 = 32'd3963
; 
32'd165900: dataIn1 = 32'd5829
; 
32'd165901: dataIn1 = 32'd6851
; 
32'd165902: dataIn1 = 32'd6854
; 
32'd165903: dataIn1 = 32'd6855
; 
32'd165904: dataIn1 = 32'd6867
; 
32'd165905: dataIn1 = 32'd6870
; 
32'd165906: dataIn1 = 32'd3963
; 
32'd165907: dataIn1 = 32'd5828
; 
32'd165908: dataIn1 = 32'd6851
; 
32'd165909: dataIn1 = 32'd6854
; 
32'd165910: dataIn1 = 32'd6855
; 
32'd165911: dataIn1 = 32'd9271
; 
32'd165912: dataIn1 = 32'd3964
; 
32'd165913: dataIn1 = 32'd5829
; 
32'd165914: dataIn1 = 32'd6852
; 
32'd165915: dataIn1 = 32'd6856
; 
32'd165916: dataIn1 = 32'd6857
; 
32'd165917: dataIn1 = 32'd6868
; 
32'd165918: dataIn1 = 32'd6871
; 
32'd165919: dataIn1 = 32'd3964
; 
32'd165920: dataIn1 = 32'd5827
; 
32'd165921: dataIn1 = 32'd6852
; 
32'd165922: dataIn1 = 32'd6856
; 
32'd165923: dataIn1 = 32'd6857
; 
32'd165924: dataIn1 = 32'd6861
; 
32'd165925: dataIn1 = 32'd6865
; 
32'd165926: dataIn1 = 32'd3965
; 
32'd165927: dataIn1 = 32'd5828
; 
32'd165928: dataIn1 = 32'd6853
; 
32'd165929: dataIn1 = 32'd6858
; 
32'd165930: dataIn1 = 32'd6859
; 
32'd165931: dataIn1 = 32'd9270
; 
32'd165932: dataIn1 = 32'd3965
; 
32'd165933: dataIn1 = 32'd5827
; 
32'd165934: dataIn1 = 32'd6853
; 
32'd165935: dataIn1 = 32'd6858
; 
32'd165936: dataIn1 = 32'd6859
; 
32'd165937: dataIn1 = 32'd6862
; 
32'd165938: dataIn1 = 32'd6866
; 
32'd165939: dataIn1 = 32'd5830
; 
32'd165940: dataIn1 = 32'd5831
; 
32'd165941: dataIn1 = 32'd6860
; 
32'd165942: dataIn1 = 32'd6861
; 
32'd165943: dataIn1 = 32'd6862
; 
32'd165944: dataIn1 = 32'd6863
; 
32'd165945: dataIn1 = 32'd6864
; 
32'd165946: dataIn1 = 32'd5827
; 
32'd165947: dataIn1 = 32'd5831
; 
32'd165948: dataIn1 = 32'd6857
; 
32'd165949: dataIn1 = 32'd6860
; 
32'd165950: dataIn1 = 32'd6861
; 
32'd165951: dataIn1 = 32'd6862
; 
32'd165952: dataIn1 = 32'd6865
; 
32'd165953: dataIn1 = 32'd5827
; 
32'd165954: dataIn1 = 32'd5830
; 
32'd165955: dataIn1 = 32'd6859
; 
32'd165956: dataIn1 = 32'd6860
; 
32'd165957: dataIn1 = 32'd6861
; 
32'd165958: dataIn1 = 32'd6862
; 
32'd165959: dataIn1 = 32'd6866
; 
32'd165960: dataIn1 = 32'd2319
; 
32'd165961: dataIn1 = 32'd5831
; 
32'd165962: dataIn1 = 32'd6860
; 
32'd165963: dataIn1 = 32'd6863
; 
32'd165964: dataIn1 = 32'd6864
; 
32'd165965: dataIn1 = 32'd6883
; 
32'd165966: dataIn1 = 32'd6886
; 
32'd165967: dataIn1 = 32'd2319
; 
32'd165968: dataIn1 = 32'd5830
; 
32'd165969: dataIn1 = 32'd6860
; 
32'd165970: dataIn1 = 32'd6863
; 
32'd165971: dataIn1 = 32'd6864
; 
32'd165972: dataIn1 = 32'd6900
; 
32'd165973: dataIn1 = 32'd6903
; 
32'd165974: dataIn1 = 32'd3964
; 
32'd165975: dataIn1 = 32'd5831
; 
32'd165976: dataIn1 = 32'd6857
; 
32'd165977: dataIn1 = 32'd6861
; 
32'd165978: dataIn1 = 32'd6865
; 
32'd165979: dataIn1 = 32'd6880
; 
32'd165980: dataIn1 = 32'd6884
; 
32'd165981: dataIn1 = 32'd3965
; 
32'd165982: dataIn1 = 32'd5830
; 
32'd165983: dataIn1 = 32'd6859
; 
32'd165984: dataIn1 = 32'd6862
; 
32'd165985: dataIn1 = 32'd6866
; 
32'd165986: dataIn1 = 32'd6902
; 
32'd165987: dataIn1 = 32'd6906
; 
32'd165988: dataIn1 = 32'd5829
; 
32'd165989: dataIn1 = 32'd5833
; 
32'd165990: dataIn1 = 32'd6854
; 
32'd165991: dataIn1 = 32'd6867
; 
32'd165992: dataIn1 = 32'd6868
; 
32'd165993: dataIn1 = 32'd6869
; 
32'd165994: dataIn1 = 32'd6870
; 
32'd165995: dataIn1 = 32'd5829
; 
32'd165996: dataIn1 = 32'd5832
; 
32'd165997: dataIn1 = 32'd6856
; 
32'd165998: dataIn1 = 32'd6867
; 
32'd165999: dataIn1 = 32'd6868
; 
32'd166000: dataIn1 = 32'd6869
; 
32'd166001: dataIn1 = 32'd6871
; 
32'd166002: dataIn1 = 32'd5832
; 
32'd166003: dataIn1 = 32'd5833
; 
32'd166004: dataIn1 = 32'd6867
; 
32'd166005: dataIn1 = 32'd6868
; 
32'd166006: dataIn1 = 32'd6869
; 
32'd166007: dataIn1 = 32'd6872
; 
32'd166008: dataIn1 = 32'd6873
; 
32'd166009: dataIn1 = 32'd3963
; 
32'd166010: dataIn1 = 32'd5833
; 
32'd166011: dataIn1 = 32'd5835
; 
32'd166012: dataIn1 = 32'd6854
; 
32'd166013: dataIn1 = 32'd6867
; 
32'd166014: dataIn1 = 32'd6870
; 
32'd166015: dataIn1 = 32'd3964
; 
32'd166016: dataIn1 = 32'd5832
; 
32'd166017: dataIn1 = 32'd6856
; 
32'd166018: dataIn1 = 32'd6868
; 
32'd166019: dataIn1 = 32'd6871
; 
32'd166020: dataIn1 = 32'd6879
; 
32'd166021: dataIn1 = 32'd6896
; 
32'd166022: dataIn1 = 32'd2321
; 
32'd166023: dataIn1 = 32'd5833
; 
32'd166024: dataIn1 = 32'd5834
; 
32'd166025: dataIn1 = 32'd6869
; 
32'd166026: dataIn1 = 32'd6872
; 
32'd166027: dataIn1 = 32'd6873
; 
32'd166028: dataIn1 = 32'd2321
; 
32'd166029: dataIn1 = 32'd5832
; 
32'd166030: dataIn1 = 32'd6869
; 
32'd166031: dataIn1 = 32'd6872
; 
32'd166032: dataIn1 = 32'd6873
; 
32'd166033: dataIn1 = 32'd6897
; 
32'd166034: dataIn1 = 32'd6899
; 
32'd166035: dataIn1 = 32'd5837
; 
32'd166036: dataIn1 = 32'd5838
; 
32'd166037: dataIn1 = 32'd6874
; 
32'd166038: dataIn1 = 32'd6875
; 
32'd166039: dataIn1 = 32'd6876
; 
32'd166040: dataIn1 = 32'd6877
; 
32'd166041: dataIn1 = 32'd6878
; 
32'd166042: dataIn1 = 32'd5836
; 
32'd166043: dataIn1 = 32'd5838
; 
32'd166044: dataIn1 = 32'd6874
; 
32'd166045: dataIn1 = 32'd6875
; 
32'd166046: dataIn1 = 32'd6876
; 
32'd166047: dataIn1 = 32'd6879
; 
32'd166048: dataIn1 = 32'd6880
; 
32'd166049: dataIn1 = 32'd5836
; 
32'd166050: dataIn1 = 32'd5837
; 
32'd166051: dataIn1 = 32'd6874
; 
32'd166052: dataIn1 = 32'd6875
; 
32'd166053: dataIn1 = 32'd6876
; 
32'd166054: dataIn1 = 32'd6881
; 
32'd166055: dataIn1 = 32'd6882
; 
32'd166056: dataIn1 = 32'd3968
; 
32'd166057: dataIn1 = 32'd5838
; 
32'd166058: dataIn1 = 32'd6874
; 
32'd166059: dataIn1 = 32'd6877
; 
32'd166060: dataIn1 = 32'd6878
; 
32'd166061: dataIn1 = 32'd6895
; 
32'd166062: dataIn1 = 32'd6898
; 
32'd166063: dataIn1 = 32'd3968
; 
32'd166064: dataIn1 = 32'd5837
; 
32'd166065: dataIn1 = 32'd6874
; 
32'd166066: dataIn1 = 32'd6877
; 
32'd166067: dataIn1 = 32'd6878
; 
32'd166068: dataIn1 = 32'd6888
; 
32'd166069: dataIn1 = 32'd6891
; 
32'd166070: dataIn1 = 32'd3964
; 
32'd166071: dataIn1 = 32'd5838
; 
32'd166072: dataIn1 = 32'd6871
; 
32'd166073: dataIn1 = 32'd6875
; 
32'd166074: dataIn1 = 32'd6879
; 
32'd166075: dataIn1 = 32'd6880
; 
32'd166076: dataIn1 = 32'd6896
; 
32'd166077: dataIn1 = 32'd3964
; 
32'd166078: dataIn1 = 32'd5836
; 
32'd166079: dataIn1 = 32'd6865
; 
32'd166080: dataIn1 = 32'd6875
; 
32'd166081: dataIn1 = 32'd6879
; 
32'd166082: dataIn1 = 32'd6880
; 
32'd166083: dataIn1 = 32'd6884
; 
32'd166084: dataIn1 = 32'd3969
; 
32'd166085: dataIn1 = 32'd5837
; 
32'd166086: dataIn1 = 32'd6876
; 
32'd166087: dataIn1 = 32'd6881
; 
32'd166088: dataIn1 = 32'd6882
; 
32'd166089: dataIn1 = 32'd6890
; 
32'd166090: dataIn1 = 32'd6894
; 
32'd166091: dataIn1 = 32'd3969
; 
32'd166092: dataIn1 = 32'd5836
; 
32'd166093: dataIn1 = 32'd6876
; 
32'd166094: dataIn1 = 32'd6881
; 
32'd166095: dataIn1 = 32'd6882
; 
32'd166096: dataIn1 = 32'd6885
; 
32'd166097: dataIn1 = 32'd6887
; 
32'd166098: dataIn1 = 32'd5831
; 
32'd166099: dataIn1 = 32'd5839
; 
32'd166100: dataIn1 = 32'd6863
; 
32'd166101: dataIn1 = 32'd6883
; 
32'd166102: dataIn1 = 32'd6884
; 
32'd166103: dataIn1 = 32'd6885
; 
32'd166104: dataIn1 = 32'd6886
; 
32'd166105: dataIn1 = 32'd5831
; 
32'd166106: dataIn1 = 32'd5836
; 
32'd166107: dataIn1 = 32'd6865
; 
32'd166108: dataIn1 = 32'd6880
; 
32'd166109: dataIn1 = 32'd6883
; 
32'd166110: dataIn1 = 32'd6884
; 
32'd166111: dataIn1 = 32'd6885
; 
32'd166112: dataIn1 = 32'd5836
; 
32'd166113: dataIn1 = 32'd5839
; 
32'd166114: dataIn1 = 32'd6882
; 
32'd166115: dataIn1 = 32'd6883
; 
32'd166116: dataIn1 = 32'd6884
; 
32'd166117: dataIn1 = 32'd6885
; 
32'd166118: dataIn1 = 32'd6887
; 
32'd166119: dataIn1 = 32'd2319
; 
32'd166120: dataIn1 = 32'd5839
; 
32'd166121: dataIn1 = 32'd6863
; 
32'd166122: dataIn1 = 32'd6883
; 
32'd166123: dataIn1 = 32'd6886
; 
32'd166124: dataIn1 = 32'd6919
; 
32'd166125: dataIn1 = 32'd6961
; 
32'd166126: dataIn1 = 32'd3969
; 
32'd166127: dataIn1 = 32'd5839
; 
32'd166128: dataIn1 = 32'd6882
; 
32'd166129: dataIn1 = 32'd6885
; 
32'd166130: dataIn1 = 32'd6887
; 
32'd166131: dataIn1 = 32'd6960
; 
32'd166132: dataIn1 = 32'd6963
; 
32'd166133: dataIn1 = 32'd5837
; 
32'd166134: dataIn1 = 32'd5841
; 
32'd166135: dataIn1 = 32'd6878
; 
32'd166136: dataIn1 = 32'd6888
; 
32'd166137: dataIn1 = 32'd6889
; 
32'd166138: dataIn1 = 32'd6890
; 
32'd166139: dataIn1 = 32'd6891
; 
32'd166140: dataIn1 = 32'd5840
; 
32'd166141: dataIn1 = 32'd5841
; 
32'd166142: dataIn1 = 32'd6888
; 
32'd166143: dataIn1 = 32'd6889
; 
32'd166144: dataIn1 = 32'd6890
; 
32'd166145: dataIn1 = 32'd6892
; 
32'd166146: dataIn1 = 32'd6893
; 
32'd166147: dataIn1 = 32'd5837
; 
32'd166148: dataIn1 = 32'd5840
; 
32'd166149: dataIn1 = 32'd6881
; 
32'd166150: dataIn1 = 32'd6888
; 
32'd166151: dataIn1 = 32'd6889
; 
32'd166152: dataIn1 = 32'd6890
; 
32'd166153: dataIn1 = 32'd6894
; 
32'd166154: dataIn1 = 32'd3968
; 
32'd166155: dataIn1 = 32'd5841
; 
32'd166156: dataIn1 = 32'd6878
; 
32'd166157: dataIn1 = 32'd6888
; 
32'd166158: dataIn1 = 32'd6891
; 
32'd166159: dataIn1 = 32'd7021
; 
32'd166160: dataIn1 = 32'd7029
; 
32'd166161: dataIn1 = 32'd127
; 
32'd166162: dataIn1 = 32'd5787
; 
32'd166163: dataIn1 = 32'd5841
; 
32'd166164: dataIn1 = 32'd6889
; 
32'd166165: dataIn1 = 32'd6892
; 
32'd166166: dataIn1 = 32'd6893
; 
32'd166167: dataIn1 = 32'd7030
; 
32'd166168: dataIn1 = 32'd127
; 
32'd166169: dataIn1 = 32'd5840
; 
32'd166170: dataIn1 = 32'd5944
; 
32'd166171: dataIn1 = 32'd6889
; 
32'd166172: dataIn1 = 32'd6892
; 
32'd166173: dataIn1 = 32'd6893
; 
32'd166174: dataIn1 = 32'd6965
; 
32'd166175: dataIn1 = 32'd3969
; 
32'd166176: dataIn1 = 32'd5840
; 
32'd166177: dataIn1 = 32'd6881
; 
32'd166178: dataIn1 = 32'd6890
; 
32'd166179: dataIn1 = 32'd6894
; 
32'd166180: dataIn1 = 32'd6959
; 
32'd166181: dataIn1 = 32'd6966
; 
32'd166182: dataIn1 = 32'd5838
; 
32'd166183: dataIn1 = 32'd5842
; 
32'd166184: dataIn1 = 32'd6877
; 
32'd166185: dataIn1 = 32'd6895
; 
32'd166186: dataIn1 = 32'd6896
; 
32'd166187: dataIn1 = 32'd6897
; 
32'd166188: dataIn1 = 32'd6898
; 
32'd166189: dataIn1 = 32'd5832
; 
32'd166190: dataIn1 = 32'd5838
; 
32'd166191: dataIn1 = 32'd6871
; 
32'd166192: dataIn1 = 32'd6879
; 
32'd166193: dataIn1 = 32'd6895
; 
32'd166194: dataIn1 = 32'd6896
; 
32'd166195: dataIn1 = 32'd6897
; 
32'd166196: dataIn1 = 32'd5832
; 
32'd166197: dataIn1 = 32'd5842
; 
32'd166198: dataIn1 = 32'd6873
; 
32'd166199: dataIn1 = 32'd6895
; 
32'd166200: dataIn1 = 32'd6896
; 
32'd166201: dataIn1 = 32'd6897
; 
32'd166202: dataIn1 = 32'd6899
; 
32'd166203: dataIn1 = 32'd3968
; 
32'd166204: dataIn1 = 32'd5842
; 
32'd166205: dataIn1 = 32'd6877
; 
32'd166206: dataIn1 = 32'd6895
; 
32'd166207: dataIn1 = 32'd6898
; 
32'd166208: dataIn1 = 32'd7020
; 
32'd166209: dataIn1 = 32'd7032
; 
32'd166210: dataIn1 = 32'd2321
; 
32'd166211: dataIn1 = 32'd5842
; 
32'd166212: dataIn1 = 32'd6873
; 
32'd166213: dataIn1 = 32'd6897
; 
32'd166214: dataIn1 = 32'd6899
; 
32'd166215: dataIn1 = 32'd7016
; 
32'd166216: dataIn1 = 32'd7034
; 
32'd166217: dataIn1 = 32'd5830
; 
32'd166218: dataIn1 = 32'd5846
; 
32'd166219: dataIn1 = 32'd6864
; 
32'd166220: dataIn1 = 32'd6900
; 
32'd166221: dataIn1 = 32'd6901
; 
32'd166222: dataIn1 = 32'd6902
; 
32'd166223: dataIn1 = 32'd6903
; 
32'd166224: dataIn1 = 32'd5843
; 
32'd166225: dataIn1 = 32'd5846
; 
32'd166226: dataIn1 = 32'd6900
; 
32'd166227: dataIn1 = 32'd6901
; 
32'd166228: dataIn1 = 32'd6902
; 
32'd166229: dataIn1 = 32'd6904
; 
32'd166230: dataIn1 = 32'd6905
; 
32'd166231: dataIn1 = 32'd5830
; 
32'd166232: dataIn1 = 32'd5843
; 
32'd166233: dataIn1 = 32'd6866
; 
32'd166234: dataIn1 = 32'd6900
; 
32'd166235: dataIn1 = 32'd6901
; 
32'd166236: dataIn1 = 32'd6902
; 
32'd166237: dataIn1 = 32'd6906
; 
32'd166238: dataIn1 = 32'd2319
; 
32'd166239: dataIn1 = 32'd5846
; 
32'd166240: dataIn1 = 32'd6864
; 
32'd166241: dataIn1 = 32'd6900
; 
32'd166242: dataIn1 = 32'd6903
; 
32'd166243: dataIn1 = 32'd6920
; 
32'd166244: dataIn1 = 32'd6981
; 
32'd166245: dataIn1 = 32'd3971
; 
32'd166246: dataIn1 = 32'd5846
; 
32'd166247: dataIn1 = 32'd6901
; 
32'd166248: dataIn1 = 32'd6904
; 
32'd166249: dataIn1 = 32'd6905
; 
32'd166250: dataIn1 = 32'd6978
; 
32'd166251: dataIn1 = 32'd6982
; 
32'd166252: dataIn1 = 32'd3971
; 
32'd166253: dataIn1 = 32'd5843
; 
32'd166254: dataIn1 = 32'd5845
; 
32'd166255: dataIn1 = 32'd6901
; 
32'd166256: dataIn1 = 32'd6904
; 
32'd166257: dataIn1 = 32'd6905
; 
32'd166258: dataIn1 = 32'd3965
; 
32'd166259: dataIn1 = 32'd5843
; 
32'd166260: dataIn1 = 32'd5844
; 
32'd166261: dataIn1 = 32'd6866
; 
32'd166262: dataIn1 = 32'd6902
; 
32'd166263: dataIn1 = 32'd6906
; 
32'd166264: dataIn1 = 32'd5850
; 
32'd166265: dataIn1 = 32'd5851
; 
32'd166266: dataIn1 = 32'd6907
; 
32'd166267: dataIn1 = 32'd6908
; 
32'd166268: dataIn1 = 32'd6909
; 
32'd166269: dataIn1 = 32'd6910
; 
32'd166270: dataIn1 = 32'd6911
; 
32'd166271: dataIn1 = 32'd5849
; 
32'd166272: dataIn1 = 32'd5851
; 
32'd166273: dataIn1 = 32'd6907
; 
32'd166274: dataIn1 = 32'd6908
; 
32'd166275: dataIn1 = 32'd6909
; 
32'd166276: dataIn1 = 32'd6912
; 
32'd166277: dataIn1 = 32'd6913
; 
32'd166278: dataIn1 = 32'd5849
; 
32'd166279: dataIn1 = 32'd5850
; 
32'd166280: dataIn1 = 32'd6907
; 
32'd166281: dataIn1 = 32'd6908
; 
32'd166282: dataIn1 = 32'd6909
; 
32'd166283: dataIn1 = 32'd6914
; 
32'd166284: dataIn1 = 32'd6915
; 
32'd166285: dataIn1 = 32'd3972
; 
32'd166286: dataIn1 = 32'd5851
; 
32'd166287: dataIn1 = 32'd6907
; 
32'd166288: dataIn1 = 32'd6910
; 
32'd166289: dataIn1 = 32'd6911
; 
32'd166290: dataIn1 = 32'd6930
; 
32'd166291: dataIn1 = 32'd6933
; 
32'd166292: dataIn1 = 32'd3972
; 
32'd166293: dataIn1 = 32'd5850
; 
32'd166294: dataIn1 = 32'd6907
; 
32'd166295: dataIn1 = 32'd6910
; 
32'd166296: dataIn1 = 32'd6911
; 
32'd166297: dataIn1 = 32'd6923
; 
32'd166298: dataIn1 = 32'd6926
; 
32'd166299: dataIn1 = 32'd3973
; 
32'd166300: dataIn1 = 32'd5851
; 
32'd166301: dataIn1 = 32'd6908
; 
32'd166302: dataIn1 = 32'd6912
; 
32'd166303: dataIn1 = 32'd6913
; 
32'd166304: dataIn1 = 32'd6931
; 
32'd166305: dataIn1 = 32'd6934
; 
32'd166306: dataIn1 = 32'd3973
; 
32'd166307: dataIn1 = 32'd5849
; 
32'd166308: dataIn1 = 32'd6908
; 
32'd166309: dataIn1 = 32'd6912
; 
32'd166310: dataIn1 = 32'd6913
; 
32'd166311: dataIn1 = 32'd6917
; 
32'd166312: dataIn1 = 32'd6921
; 
32'd166313: dataIn1 = 32'd3974
; 
32'd166314: dataIn1 = 32'd5850
; 
32'd166315: dataIn1 = 32'd6909
; 
32'd166316: dataIn1 = 32'd6914
; 
32'd166317: dataIn1 = 32'd6915
; 
32'd166318: dataIn1 = 32'd6925
; 
32'd166319: dataIn1 = 32'd6929
; 
32'd166320: dataIn1 = 32'd3974
; 
32'd166321: dataIn1 = 32'd5849
; 
32'd166322: dataIn1 = 32'd6909
; 
32'd166323: dataIn1 = 32'd6914
; 
32'd166324: dataIn1 = 32'd6915
; 
32'd166325: dataIn1 = 32'd6918
; 
32'd166326: dataIn1 = 32'd6922
; 
32'd166327: dataIn1 = 32'd5852
; 
32'd166328: dataIn1 = 32'd5853
; 
32'd166329: dataIn1 = 32'd6916
; 
32'd166330: dataIn1 = 32'd6917
; 
32'd166331: dataIn1 = 32'd6918
; 
32'd166332: dataIn1 = 32'd6919
; 
32'd166333: dataIn1 = 32'd6920
; 
32'd166334: dataIn1 = 32'd5849
; 
32'd166335: dataIn1 = 32'd5853
; 
32'd166336: dataIn1 = 32'd6913
; 
32'd166337: dataIn1 = 32'd6916
; 
32'd166338: dataIn1 = 32'd6917
; 
32'd166339: dataIn1 = 32'd6918
; 
32'd166340: dataIn1 = 32'd6921
; 
32'd166341: dataIn1 = 32'd5849
; 
32'd166342: dataIn1 = 32'd5852
; 
32'd166343: dataIn1 = 32'd6915
; 
32'd166344: dataIn1 = 32'd6916
; 
32'd166345: dataIn1 = 32'd6917
; 
32'd166346: dataIn1 = 32'd6918
; 
32'd166347: dataIn1 = 32'd6922
; 
32'd166348: dataIn1 = 32'd2319
; 
32'd166349: dataIn1 = 32'd5853
; 
32'd166350: dataIn1 = 32'd6886
; 
32'd166351: dataIn1 = 32'd6916
; 
32'd166352: dataIn1 = 32'd6919
; 
32'd166353: dataIn1 = 32'd6920
; 
32'd166354: dataIn1 = 32'd6961
; 
32'd166355: dataIn1 = 32'd2319
; 
32'd166356: dataIn1 = 32'd5852
; 
32'd166357: dataIn1 = 32'd6903
; 
32'd166358: dataIn1 = 32'd6916
; 
32'd166359: dataIn1 = 32'd6919
; 
32'd166360: dataIn1 = 32'd6920
; 
32'd166361: dataIn1 = 32'd6981
; 
32'd166362: dataIn1 = 32'd3973
; 
32'd166363: dataIn1 = 32'd5853
; 
32'd166364: dataIn1 = 32'd6913
; 
32'd166365: dataIn1 = 32'd6917
; 
32'd166366: dataIn1 = 32'd6921
; 
32'd166367: dataIn1 = 32'd6958
; 
32'd166368: dataIn1 = 32'd6962
; 
32'd166369: dataIn1 = 32'd3974
; 
32'd166370: dataIn1 = 32'd5852
; 
32'd166371: dataIn1 = 32'd6915
; 
32'd166372: dataIn1 = 32'd6918
; 
32'd166373: dataIn1 = 32'd6922
; 
32'd166374: dataIn1 = 32'd6980
; 
32'd166375: dataIn1 = 32'd6983
; 
32'd166376: dataIn1 = 32'd5850
; 
32'd166377: dataIn1 = 32'd5855
; 
32'd166378: dataIn1 = 32'd6911
; 
32'd166379: dataIn1 = 32'd6923
; 
32'd166380: dataIn1 = 32'd6924
; 
32'd166381: dataIn1 = 32'd6925
; 
32'd166382: dataIn1 = 32'd6926
; 
32'd166383: dataIn1 = 32'd5854
; 
32'd166384: dataIn1 = 32'd5855
; 
32'd166385: dataIn1 = 32'd6923
; 
32'd166386: dataIn1 = 32'd6924
; 
32'd166387: dataIn1 = 32'd6925
; 
32'd166388: dataIn1 = 32'd6927
; 
32'd166389: dataIn1 = 32'd6928
; 
32'd166390: dataIn1 = 32'd5850
; 
32'd166391: dataIn1 = 32'd5854
; 
32'd166392: dataIn1 = 32'd6914
; 
32'd166393: dataIn1 = 32'd6923
; 
32'd166394: dataIn1 = 32'd6924
; 
32'd166395: dataIn1 = 32'd6925
; 
32'd166396: dataIn1 = 32'd6929
; 
32'd166397: dataIn1 = 32'd3972
; 
32'd166398: dataIn1 = 32'd5855
; 
32'd166399: dataIn1 = 32'd6911
; 
32'd166400: dataIn1 = 32'd6923
; 
32'd166401: dataIn1 = 32'd6926
; 
32'd166402: dataIn1 = 32'd6941
; 
32'd166403: dataIn1 = 32'd6946
; 
32'd166404: dataIn1 = 32'd2322
; 
32'd166405: dataIn1 = 32'd5855
; 
32'd166406: dataIn1 = 32'd6924
; 
32'd166407: dataIn1 = 32'd6927
; 
32'd166408: dataIn1 = 32'd6928
; 
32'd166409: dataIn1 = 32'd6947
; 
32'd166410: dataIn1 = 32'd6949
; 
32'd166411: dataIn1 = 32'd2322
; 
32'd166412: dataIn1 = 32'd5854
; 
32'd166413: dataIn1 = 32'd6924
; 
32'd166414: dataIn1 = 32'd6927
; 
32'd166415: dataIn1 = 32'd6928
; 
32'd166416: dataIn1 = 32'd6985
; 
32'd166417: dataIn1 = 32'd6988
; 
32'd166418: dataIn1 = 32'd3974
; 
32'd166419: dataIn1 = 32'd5854
; 
32'd166420: dataIn1 = 32'd6914
; 
32'd166421: dataIn1 = 32'd6925
; 
32'd166422: dataIn1 = 32'd6929
; 
32'd166423: dataIn1 = 32'd6979
; 
32'd166424: dataIn1 = 32'd6986
; 
32'd166425: dataIn1 = 32'd5851
; 
32'd166426: dataIn1 = 32'd5857
; 
32'd166427: dataIn1 = 32'd6910
; 
32'd166428: dataIn1 = 32'd6930
; 
32'd166429: dataIn1 = 32'd6931
; 
32'd166430: dataIn1 = 32'd6932
; 
32'd166431: dataIn1 = 32'd6933
; 
32'd166432: dataIn1 = 32'd5851
; 
32'd166433: dataIn1 = 32'd5856
; 
32'd166434: dataIn1 = 32'd6912
; 
32'd166435: dataIn1 = 32'd6930
; 
32'd166436: dataIn1 = 32'd6931
; 
32'd166437: dataIn1 = 32'd6932
; 
32'd166438: dataIn1 = 32'd6934
; 
32'd166439: dataIn1 = 32'd5856
; 
32'd166440: dataIn1 = 32'd5857
; 
32'd166441: dataIn1 = 32'd6930
; 
32'd166442: dataIn1 = 32'd6931
; 
32'd166443: dataIn1 = 32'd6932
; 
32'd166444: dataIn1 = 32'd6935
; 
32'd166445: dataIn1 = 32'd6936
; 
32'd166446: dataIn1 = 32'd3972
; 
32'd166447: dataIn1 = 32'd5857
; 
32'd166448: dataIn1 = 32'd6910
; 
32'd166449: dataIn1 = 32'd6930
; 
32'd166450: dataIn1 = 32'd6933
; 
32'd166451: dataIn1 = 32'd6940
; 
32'd166452: dataIn1 = 32'd6951
; 
32'd166453: dataIn1 = 32'd3973
; 
32'd166454: dataIn1 = 32'd5856
; 
32'd166455: dataIn1 = 32'd6912
; 
32'd166456: dataIn1 = 32'd6931
; 
32'd166457: dataIn1 = 32'd6934
; 
32'd166458: dataIn1 = 32'd6957
; 
32'd166459: dataIn1 = 32'd6968
; 
32'd166460: dataIn1 = 32'd1104
; 
32'd166461: dataIn1 = 32'd4837
; 
32'd166462: dataIn1 = 32'd5857
; 
32'd166463: dataIn1 = 32'd6932
; 
32'd166464: dataIn1 = 32'd6935
; 
32'd166465: dataIn1 = 32'd6936
; 
32'd166466: dataIn1 = 32'd1104
; 
32'd166467: dataIn1 = 32'd5856
; 
32'd166468: dataIn1 = 32'd6932
; 
32'd166469: dataIn1 = 32'd6935
; 
32'd166470: dataIn1 = 32'd6936
; 
32'd166471: dataIn1 = 32'd6969
; 
32'd166472: dataIn1 = 32'd6971
; 
32'd166473: dataIn1 = 32'd5859
; 
32'd166474: dataIn1 = 32'd5860
; 
32'd166475: dataIn1 = 32'd6937
; 
32'd166476: dataIn1 = 32'd6938
; 
32'd166477: dataIn1 = 32'd6939
; 
32'd166478: dataIn1 = 32'd6940
; 
32'd166479: dataIn1 = 32'd6941
; 
32'd166480: dataIn1 = 32'd2621
; 
32'd166481: dataIn1 = 32'd5858
; 
32'd166482: dataIn1 = 32'd5860
; 
32'd166483: dataIn1 = 32'd6937
; 
32'd166484: dataIn1 = 32'd6938
; 
32'd166485: dataIn1 = 32'd6939
; 
32'd166486: dataIn1 = 32'd5858
; 
32'd166487: dataIn1 = 32'd5859
; 
32'd166488: dataIn1 = 32'd6937
; 
32'd166489: dataIn1 = 32'd6938
; 
32'd166490: dataIn1 = 32'd6939
; 
32'd166491: dataIn1 = 32'd6942
; 
32'd166492: dataIn1 = 32'd6943
; 
32'd166493: dataIn1 = 32'd3972
; 
32'd166494: dataIn1 = 32'd5860
; 
32'd166495: dataIn1 = 32'd6933
; 
32'd166496: dataIn1 = 32'd6937
; 
32'd166497: dataIn1 = 32'd6940
; 
32'd166498: dataIn1 = 32'd6941
; 
32'd166499: dataIn1 = 32'd6951
; 
32'd166500: dataIn1 = 32'd3972
; 
32'd166501: dataIn1 = 32'd5859
; 
32'd166502: dataIn1 = 32'd6926
; 
32'd166503: dataIn1 = 32'd6937
; 
32'd166504: dataIn1 = 32'd6940
; 
32'd166505: dataIn1 = 32'd6941
; 
32'd166506: dataIn1 = 32'd6946
; 
32'd166507: dataIn1 = 32'd3975
; 
32'd166508: dataIn1 = 32'd5859
; 
32'd166509: dataIn1 = 32'd6939
; 
32'd166510: dataIn1 = 32'd6942
; 
32'd166511: dataIn1 = 32'd6943
; 
32'd166512: dataIn1 = 32'd6948
; 
32'd166513: dataIn1 = 32'd6950
; 
32'd166514: dataIn1 = 32'd3975
; 
32'd166515: dataIn1 = 32'd5858
; 
32'd166516: dataIn1 = 32'd6939
; 
32'd166517: dataIn1 = 32'd6942
; 
32'd166518: dataIn1 = 32'd6943
; 
32'd166519: dataIn1 = 32'd6944
; 
32'd166520: dataIn1 = 32'd6945
; 
32'd166521: dataIn1 = 32'd3975
; 
32'd166522: dataIn1 = 32'd5861
; 
32'd166523: dataIn1 = 32'd6943
; 
32'd166524: dataIn1 = 32'd6944
; 
32'd166525: dataIn1 = 32'd6945
; 
32'd166526: dataIn1 = 32'd8899
; 
32'd166527: dataIn1 = 32'd8903
; 
32'd166528: dataIn1 = 32'd4836
; 
32'd166529: dataIn1 = 32'd5858
; 
32'd166530: dataIn1 = 32'd5861
; 
32'd166531: dataIn1 = 32'd6943
; 
32'd166532: dataIn1 = 32'd6944
; 
32'd166533: dataIn1 = 32'd6945
; 
32'd166534: dataIn1 = 32'd5855
; 
32'd166535: dataIn1 = 32'd5859
; 
32'd166536: dataIn1 = 32'd6926
; 
32'd166537: dataIn1 = 32'd6941
; 
32'd166538: dataIn1 = 32'd6946
; 
32'd166539: dataIn1 = 32'd6947
; 
32'd166540: dataIn1 = 32'd6948
; 
32'd166541: dataIn1 = 32'd5855
; 
32'd166542: dataIn1 = 32'd5862
; 
32'd166543: dataIn1 = 32'd6927
; 
32'd166544: dataIn1 = 32'd6946
; 
32'd166545: dataIn1 = 32'd6947
; 
32'd166546: dataIn1 = 32'd6948
; 
32'd166547: dataIn1 = 32'd6949
; 
32'd166548: dataIn1 = 32'd5859
; 
32'd166549: dataIn1 = 32'd5862
; 
32'd166550: dataIn1 = 32'd6942
; 
32'd166551: dataIn1 = 32'd6946
; 
32'd166552: dataIn1 = 32'd6947
; 
32'd166553: dataIn1 = 32'd6948
; 
32'd166554: dataIn1 = 32'd6950
; 
32'd166555: dataIn1 = 32'd2322
; 
32'd166556: dataIn1 = 32'd5862
; 
32'd166557: dataIn1 = 32'd6927
; 
32'd166558: dataIn1 = 32'd6947
; 
32'd166559: dataIn1 = 32'd6949
; 
32'd166560: dataIn1 = 32'd8891
; 
32'd166561: dataIn1 = 32'd8910
; 
32'd166562: dataIn1 = 32'd3975
; 
32'd166563: dataIn1 = 32'd5862
; 
32'd166564: dataIn1 = 32'd6942
; 
32'd166565: dataIn1 = 32'd6948
; 
32'd166566: dataIn1 = 32'd6950
; 
32'd166567: dataIn1 = 32'd8898
; 
32'd166568: dataIn1 = 32'd8909
; 
32'd166569: dataIn1 = 32'd4837
; 
32'd166570: dataIn1 = 32'd5857
; 
32'd166571: dataIn1 = 32'd5860
; 
32'd166572: dataIn1 = 32'd6933
; 
32'd166573: dataIn1 = 32'd6940
; 
32'd166574: dataIn1 = 32'd6951
; 
32'd166575: dataIn1 = 32'd5864
; 
32'd166576: dataIn1 = 32'd5865
; 
32'd166577: dataIn1 = 32'd6952
; 
32'd166578: dataIn1 = 32'd6953
; 
32'd166579: dataIn1 = 32'd6954
; 
32'd166580: dataIn1 = 32'd6955
; 
32'd166581: dataIn1 = 32'd6956
; 
32'd166582: dataIn1 = 32'd5863
; 
32'd166583: dataIn1 = 32'd5865
; 
32'd166584: dataIn1 = 32'd6952
; 
32'd166585: dataIn1 = 32'd6953
; 
32'd166586: dataIn1 = 32'd6954
; 
32'd166587: dataIn1 = 32'd6957
; 
32'd166588: dataIn1 = 32'd6958
; 
32'd166589: dataIn1 = 32'd5863
; 
32'd166590: dataIn1 = 32'd5864
; 
32'd166591: dataIn1 = 32'd6952
; 
32'd166592: dataIn1 = 32'd6953
; 
32'd166593: dataIn1 = 32'd6954
; 
32'd166594: dataIn1 = 32'd6959
; 
32'd166595: dataIn1 = 32'd6960
; 
32'd166596: dataIn1 = 32'd2620
; 
32'd166597: dataIn1 = 32'd5865
; 
32'd166598: dataIn1 = 32'd6952
; 
32'd166599: dataIn1 = 32'd6955
; 
32'd166600: dataIn1 = 32'd6956
; 
32'd166601: dataIn1 = 32'd6967
; 
32'd166602: dataIn1 = 32'd6970
; 
32'd166603: dataIn1 = 32'd2620
; 
32'd166604: dataIn1 = 32'd5864
; 
32'd166605: dataIn1 = 32'd5945
; 
32'd166606: dataIn1 = 32'd6952
; 
32'd166607: dataIn1 = 32'd6955
; 
32'd166608: dataIn1 = 32'd6956
; 
32'd166609: dataIn1 = 32'd6964
; 
32'd166610: dataIn1 = 32'd3973
; 
32'd166611: dataIn1 = 32'd5865
; 
32'd166612: dataIn1 = 32'd6934
; 
32'd166613: dataIn1 = 32'd6953
; 
32'd166614: dataIn1 = 32'd6957
; 
32'd166615: dataIn1 = 32'd6958
; 
32'd166616: dataIn1 = 32'd6968
; 
32'd166617: dataIn1 = 32'd3973
; 
32'd166618: dataIn1 = 32'd5863
; 
32'd166619: dataIn1 = 32'd6921
; 
32'd166620: dataIn1 = 32'd6953
; 
32'd166621: dataIn1 = 32'd6957
; 
32'd166622: dataIn1 = 32'd6958
; 
32'd166623: dataIn1 = 32'd6962
; 
32'd166624: dataIn1 = 32'd3969
; 
32'd166625: dataIn1 = 32'd5864
; 
32'd166626: dataIn1 = 32'd6894
; 
32'd166627: dataIn1 = 32'd6954
; 
32'd166628: dataIn1 = 32'd6959
; 
32'd166629: dataIn1 = 32'd6960
; 
32'd166630: dataIn1 = 32'd6966
; 
32'd166631: dataIn1 = 32'd3969
; 
32'd166632: dataIn1 = 32'd5863
; 
32'd166633: dataIn1 = 32'd6887
; 
32'd166634: dataIn1 = 32'd6954
; 
32'd166635: dataIn1 = 32'd6959
; 
32'd166636: dataIn1 = 32'd6960
; 
32'd166637: dataIn1 = 32'd6963
; 
32'd166638: dataIn1 = 32'd5839
; 
32'd166639: dataIn1 = 32'd5853
; 
32'd166640: dataIn1 = 32'd6886
; 
32'd166641: dataIn1 = 32'd6919
; 
32'd166642: dataIn1 = 32'd6961
; 
32'd166643: dataIn1 = 32'd6962
; 
32'd166644: dataIn1 = 32'd6963
; 
32'd166645: dataIn1 = 32'd5853
; 
32'd166646: dataIn1 = 32'd5863
; 
32'd166647: dataIn1 = 32'd6921
; 
32'd166648: dataIn1 = 32'd6958
; 
32'd166649: dataIn1 = 32'd6961
; 
32'd166650: dataIn1 = 32'd6962
; 
32'd166651: dataIn1 = 32'd6963
; 
32'd166652: dataIn1 = 32'd5839
; 
32'd166653: dataIn1 = 32'd5863
; 
32'd166654: dataIn1 = 32'd6887
; 
32'd166655: dataIn1 = 32'd6960
; 
32'd166656: dataIn1 = 32'd6961
; 
32'd166657: dataIn1 = 32'd6962
; 
32'd166658: dataIn1 = 32'd6963
; 
32'd166659: dataIn1 = 32'd4830
; 
32'd166660: dataIn1 = 32'd5864
; 
32'd166661: dataIn1 = 32'd5945
; 
32'd166662: dataIn1 = 32'd6956
; 
32'd166663: dataIn1 = 32'd6964
; 
32'd166664: dataIn1 = 32'd6965
; 
32'd166665: dataIn1 = 32'd6966
; 
32'd166666: dataIn1 = 32'd4830
; 
32'd166667: dataIn1 = 32'd5840
; 
32'd166668: dataIn1 = 32'd5944
; 
32'd166669: dataIn1 = 32'd6893
; 
32'd166670: dataIn1 = 32'd6964
; 
32'd166671: dataIn1 = 32'd6965
; 
32'd166672: dataIn1 = 32'd6966
; 
32'd166673: dataIn1 = 32'd5840
; 
32'd166674: dataIn1 = 32'd5864
; 
32'd166675: dataIn1 = 32'd6894
; 
32'd166676: dataIn1 = 32'd6959
; 
32'd166677: dataIn1 = 32'd6964
; 
32'd166678: dataIn1 = 32'd6965
; 
32'd166679: dataIn1 = 32'd6966
; 
32'd166680: dataIn1 = 32'd4831
; 
32'd166681: dataIn1 = 32'd5865
; 
32'd166682: dataIn1 = 32'd6955
; 
32'd166683: dataIn1 = 32'd6967
; 
32'd166684: dataIn1 = 32'd6968
; 
32'd166685: dataIn1 = 32'd6969
; 
32'd166686: dataIn1 = 32'd6970
; 
32'd166687: dataIn1 = 32'd5856
; 
32'd166688: dataIn1 = 32'd5865
; 
32'd166689: dataIn1 = 32'd6934
; 
32'd166690: dataIn1 = 32'd6957
; 
32'd166691: dataIn1 = 32'd6967
; 
32'd166692: dataIn1 = 32'd6968
; 
32'd166693: dataIn1 = 32'd6969
; 
32'd166694: dataIn1 = 32'd4831
; 
32'd166695: dataIn1 = 32'd5856
; 
32'd166696: dataIn1 = 32'd6936
; 
32'd166697: dataIn1 = 32'd6967
; 
32'd166698: dataIn1 = 32'd6968
; 
32'd166699: dataIn1 = 32'd6969
; 
32'd166700: dataIn1 = 32'd6971
; 
32'd166701: dataIn1 = 32'd2620
; 
32'd166702: dataIn1 = 32'd4829
; 
32'd166703: dataIn1 = 32'd4831
; 
32'd166704: dataIn1 = 32'd6955
; 
32'd166705: dataIn1 = 32'd6967
; 
32'd166706: dataIn1 = 32'd6970
; 
32'd166707: dataIn1 = 32'd1104
; 
32'd166708: dataIn1 = 32'd4826
; 
32'd166709: dataIn1 = 32'd4831
; 
32'd166710: dataIn1 = 32'd6936
; 
32'd166711: dataIn1 = 32'd6969
; 
32'd166712: dataIn1 = 32'd6971
; 
32'd166713: dataIn1 = 32'd5867
; 
32'd166714: dataIn1 = 32'd5868
; 
32'd166715: dataIn1 = 32'd6972
; 
32'd166716: dataIn1 = 32'd6973
; 
32'd166717: dataIn1 = 32'd6974
; 
32'd166718: dataIn1 = 32'd6975
; 
32'd166719: dataIn1 = 32'd6976
; 
32'd166720: dataIn1 = 32'd5866
; 
32'd166721: dataIn1 = 32'd5868
; 
32'd166722: dataIn1 = 32'd6972
; 
32'd166723: dataIn1 = 32'd6973
; 
32'd166724: dataIn1 = 32'd6974
; 
32'd166725: dataIn1 = 32'd6977
; 
32'd166726: dataIn1 = 32'd6978
; 
32'd166727: dataIn1 = 32'd5866
; 
32'd166728: dataIn1 = 32'd5867
; 
32'd166729: dataIn1 = 32'd6972
; 
32'd166730: dataIn1 = 32'd6973
; 
32'd166731: dataIn1 = 32'd6974
; 
32'd166732: dataIn1 = 32'd6979
; 
32'd166733: dataIn1 = 32'd6980
; 
32'd166734: dataIn1 = 32'd3976
; 
32'd166735: dataIn1 = 32'd5868
; 
32'd166736: dataIn1 = 32'd5870
; 
32'd166737: dataIn1 = 32'd6972
; 
32'd166738: dataIn1 = 32'd6975
; 
32'd166739: dataIn1 = 32'd6976
; 
32'd166740: dataIn1 = 32'd3976
; 
32'd166741: dataIn1 = 32'd5867
; 
32'd166742: dataIn1 = 32'd6972
; 
32'd166743: dataIn1 = 32'd6975
; 
32'd166744: dataIn1 = 32'd6976
; 
32'd166745: dataIn1 = 32'd6984
; 
32'd166746: dataIn1 = 32'd6987
; 
32'd166747: dataIn1 = 32'd3971
; 
32'd166748: dataIn1 = 32'd5847
; 
32'd166749: dataIn1 = 32'd5868
; 
32'd166750: dataIn1 = 32'd6973
; 
32'd166751: dataIn1 = 32'd6977
; 
32'd166752: dataIn1 = 32'd6978
; 
32'd166753: dataIn1 = 32'd3971
; 
32'd166754: dataIn1 = 32'd5866
; 
32'd166755: dataIn1 = 32'd6904
; 
32'd166756: dataIn1 = 32'd6973
; 
32'd166757: dataIn1 = 32'd6977
; 
32'd166758: dataIn1 = 32'd6978
; 
32'd166759: dataIn1 = 32'd6982
; 
32'd166760: dataIn1 = 32'd3974
; 
32'd166761: dataIn1 = 32'd5867
; 
32'd166762: dataIn1 = 32'd6929
; 
32'd166763: dataIn1 = 32'd6974
; 
32'd166764: dataIn1 = 32'd6979
; 
32'd166765: dataIn1 = 32'd6980
; 
32'd166766: dataIn1 = 32'd6986
; 
32'd166767: dataIn1 = 32'd3974
; 
32'd166768: dataIn1 = 32'd5866
; 
32'd166769: dataIn1 = 32'd6922
; 
32'd166770: dataIn1 = 32'd6974
; 
32'd166771: dataIn1 = 32'd6979
; 
32'd166772: dataIn1 = 32'd6980
; 
32'd166773: dataIn1 = 32'd6983
; 
32'd166774: dataIn1 = 32'd5846
; 
32'd166775: dataIn1 = 32'd5852
; 
32'd166776: dataIn1 = 32'd6903
; 
32'd166777: dataIn1 = 32'd6920
; 
32'd166778: dataIn1 = 32'd6981
; 
32'd166779: dataIn1 = 32'd6982
; 
32'd166780: dataIn1 = 32'd6983
; 
32'd166781: dataIn1 = 32'd5846
; 
32'd166782: dataIn1 = 32'd5866
; 
32'd166783: dataIn1 = 32'd6904
; 
32'd166784: dataIn1 = 32'd6978
; 
32'd166785: dataIn1 = 32'd6981
; 
32'd166786: dataIn1 = 32'd6982
; 
32'd166787: dataIn1 = 32'd6983
; 
32'd166788: dataIn1 = 32'd5852
; 
32'd166789: dataIn1 = 32'd5866
; 
32'd166790: dataIn1 = 32'd6922
; 
32'd166791: dataIn1 = 32'd6980
; 
32'd166792: dataIn1 = 32'd6981
; 
32'd166793: dataIn1 = 32'd6982
; 
32'd166794: dataIn1 = 32'd6983
; 
32'd166795: dataIn1 = 32'd5867
; 
32'd166796: dataIn1 = 32'd5869
; 
32'd166797: dataIn1 = 32'd6976
; 
32'd166798: dataIn1 = 32'd6984
; 
32'd166799: dataIn1 = 32'd6985
; 
32'd166800: dataIn1 = 32'd6986
; 
32'd166801: dataIn1 = 32'd6987
; 
32'd166802: dataIn1 = 32'd5854
; 
32'd166803: dataIn1 = 32'd5869
; 
32'd166804: dataIn1 = 32'd6928
; 
32'd166805: dataIn1 = 32'd6984
; 
32'd166806: dataIn1 = 32'd6985
; 
32'd166807: dataIn1 = 32'd6986
; 
32'd166808: dataIn1 = 32'd6988
; 
32'd166809: dataIn1 = 32'd5854
; 
32'd166810: dataIn1 = 32'd5867
; 
32'd166811: dataIn1 = 32'd6929
; 
32'd166812: dataIn1 = 32'd6979
; 
32'd166813: dataIn1 = 32'd6984
; 
32'd166814: dataIn1 = 32'd6985
; 
32'd166815: dataIn1 = 32'd6986
; 
32'd166816: dataIn1 = 32'd3976
; 
32'd166817: dataIn1 = 32'd5869
; 
32'd166818: dataIn1 = 32'd6976
; 
32'd166819: dataIn1 = 32'd6984
; 
32'd166820: dataIn1 = 32'd6987
; 
32'd166821: dataIn1 = 32'd8911
; 
32'd166822: dataIn1 = 32'd8914
; 
32'd166823: dataIn1 = 32'd2322
; 
32'd166824: dataIn1 = 32'd5869
; 
32'd166825: dataIn1 = 32'd6928
; 
32'd166826: dataIn1 = 32'd6985
; 
32'd166827: dataIn1 = 32'd6988
; 
32'd166828: dataIn1 = 32'd8892
; 
32'd166829: dataIn1 = 32'd8913
; 
32'd166830: dataIn1 = 32'd5872
; 
32'd166831: dataIn1 = 32'd5873
; 
32'd166832: dataIn1 = 32'd6989
; 
32'd166833: dataIn1 = 32'd6990
; 
32'd166834: dataIn1 = 32'd6991
; 
32'd166835: dataIn1 = 32'd6992
; 
32'd166836: dataIn1 = 32'd6993
; 
32'd166837: dataIn1 = 32'd5871
; 
32'd166838: dataIn1 = 32'd5873
; 
32'd166839: dataIn1 = 32'd6989
; 
32'd166840: dataIn1 = 32'd6990
; 
32'd166841: dataIn1 = 32'd6991
; 
32'd166842: dataIn1 = 32'd6994
; 
32'd166843: dataIn1 = 32'd6995
; 
32'd166844: dataIn1 = 32'd5871
; 
32'd166845: dataIn1 = 32'd5872
; 
32'd166846: dataIn1 = 32'd6989
; 
32'd166847: dataIn1 = 32'd6990
; 
32'd166848: dataIn1 = 32'd6991
; 
32'd166849: dataIn1 = 32'd6996
; 
32'd166850: dataIn1 = 32'd6997
; 
32'd166851: dataIn1 = 32'd3981
; 
32'd166852: dataIn1 = 32'd5873
; 
32'd166853: dataIn1 = 32'd6989
; 
32'd166854: dataIn1 = 32'd6992
; 
32'd166855: dataIn1 = 32'd6993
; 
32'd166856: dataIn1 = 32'd7010
; 
32'd166857: dataIn1 = 32'd7013
; 
32'd166858: dataIn1 = 32'd3981
; 
32'd166859: dataIn1 = 32'd5872
; 
32'd166860: dataIn1 = 32'd6989
; 
32'd166861: dataIn1 = 32'd6992
; 
32'd166862: dataIn1 = 32'd6993
; 
32'd166863: dataIn1 = 32'd7005
; 
32'd166864: dataIn1 = 32'd7008
; 
32'd166865: dataIn1 = 32'd3982
; 
32'd166866: dataIn1 = 32'd5873
; 
32'd166867: dataIn1 = 32'd6990
; 
32'd166868: dataIn1 = 32'd6994
; 
32'd166869: dataIn1 = 32'd6995
; 
32'd166870: dataIn1 = 32'd7011
; 
32'd166871: dataIn1 = 32'd7014
; 
32'd166872: dataIn1 = 32'd3982
; 
32'd166873: dataIn1 = 32'd5871
; 
32'd166874: dataIn1 = 32'd6990
; 
32'd166875: dataIn1 = 32'd6994
; 
32'd166876: dataIn1 = 32'd6995
; 
32'd166877: dataIn1 = 32'd6999
; 
32'd166878: dataIn1 = 32'd7003
; 
32'd166879: dataIn1 = 32'd3983
; 
32'd166880: dataIn1 = 32'd5872
; 
32'd166881: dataIn1 = 32'd6991
; 
32'd166882: dataIn1 = 32'd6996
; 
32'd166883: dataIn1 = 32'd6997
; 
32'd166884: dataIn1 = 32'd7007
; 
32'd166885: dataIn1 = 32'd7009
; 
32'd166886: dataIn1 = 32'd3983
; 
32'd166887: dataIn1 = 32'd5871
; 
32'd166888: dataIn1 = 32'd6991
; 
32'd166889: dataIn1 = 32'd6996
; 
32'd166890: dataIn1 = 32'd6997
; 
32'd166891: dataIn1 = 32'd7000
; 
32'd166892: dataIn1 = 32'd7004
; 
32'd166893: dataIn1 = 32'd5874
; 
32'd166894: dataIn1 = 32'd5875
; 
32'd166895: dataIn1 = 32'd6998
; 
32'd166896: dataIn1 = 32'd6999
; 
32'd166897: dataIn1 = 32'd7000
; 
32'd166898: dataIn1 = 32'd7001
; 
32'd166899: dataIn1 = 32'd7002
; 
32'd166900: dataIn1 = 32'd5871
; 
32'd166901: dataIn1 = 32'd5875
; 
32'd166902: dataIn1 = 32'd6995
; 
32'd166903: dataIn1 = 32'd6998
; 
32'd166904: dataIn1 = 32'd6999
; 
32'd166905: dataIn1 = 32'd7000
; 
32'd166906: dataIn1 = 32'd7003
; 
32'd166907: dataIn1 = 32'd5871
; 
32'd166908: dataIn1 = 32'd5874
; 
32'd166909: dataIn1 = 32'd6997
; 
32'd166910: dataIn1 = 32'd6998
; 
32'd166911: dataIn1 = 32'd6999
; 
32'd166912: dataIn1 = 32'd7000
; 
32'd166913: dataIn1 = 32'd7004
; 
32'd166914: dataIn1 = 32'd449
; 
32'd166915: dataIn1 = 32'd5793
; 
32'd166916: dataIn1 = 32'd5875
; 
32'd166917: dataIn1 = 32'd6998
; 
32'd166918: dataIn1 = 32'd7001
; 
32'd166919: dataIn1 = 32'd7002
; 
32'd166920: dataIn1 = 32'd7026
; 
32'd166921: dataIn1 = 32'd449
; 
32'd166922: dataIn1 = 32'd5821
; 
32'd166923: dataIn1 = 32'd5874
; 
32'd166924: dataIn1 = 32'd6998
; 
32'd166925: dataIn1 = 32'd7001
; 
32'd166926: dataIn1 = 32'd7002
; 
32'd166927: dataIn1 = 32'd7044
; 
32'd166928: dataIn1 = 32'd3982
; 
32'd166929: dataIn1 = 32'd5875
; 
32'd166930: dataIn1 = 32'd6995
; 
32'd166931: dataIn1 = 32'd6999
; 
32'd166932: dataIn1 = 32'd7003
; 
32'd166933: dataIn1 = 32'd7023
; 
32'd166934: dataIn1 = 32'd7027
; 
32'd166935: dataIn1 = 32'd3983
; 
32'd166936: dataIn1 = 32'd5874
; 
32'd166937: dataIn1 = 32'd6997
; 
32'd166938: dataIn1 = 32'd7000
; 
32'd166939: dataIn1 = 32'd7004
; 
32'd166940: dataIn1 = 32'd7043
; 
32'd166941: dataIn1 = 32'd7046
; 
32'd166942: dataIn1 = 32'd5872
; 
32'd166943: dataIn1 = 32'd5877
; 
32'd166944: dataIn1 = 32'd6993
; 
32'd166945: dataIn1 = 32'd7005
; 
32'd166946: dataIn1 = 32'd7006
; 
32'd166947: dataIn1 = 32'd7007
; 
32'd166948: dataIn1 = 32'd7008
; 
32'd166949: dataIn1 = 32'd2325
; 
32'd166950: dataIn1 = 32'd5876
; 
32'd166951: dataIn1 = 32'd5877
; 
32'd166952: dataIn1 = 32'd7005
; 
32'd166953: dataIn1 = 32'd7006
; 
32'd166954: dataIn1 = 32'd7007
; 
32'd166955: dataIn1 = 32'd5872
; 
32'd166956: dataIn1 = 32'd5876
; 
32'd166957: dataIn1 = 32'd6996
; 
32'd166958: dataIn1 = 32'd7005
; 
32'd166959: dataIn1 = 32'd7006
; 
32'd166960: dataIn1 = 32'd7007
; 
32'd166961: dataIn1 = 32'd7009
; 
32'd166962: dataIn1 = 32'd3981
; 
32'd166963: dataIn1 = 32'd5877
; 
32'd166964: dataIn1 = 32'd6993
; 
32'd166965: dataIn1 = 32'd7005
; 
32'd166966: dataIn1 = 32'd7008
; 
32'd166967: dataIn1 = 32'd9273
; 
32'd166968: dataIn1 = 32'd3983
; 
32'd166969: dataIn1 = 32'd5876
; 
32'd166970: dataIn1 = 32'd6996
; 
32'd166971: dataIn1 = 32'd7007
; 
32'd166972: dataIn1 = 32'd7009
; 
32'd166973: dataIn1 = 32'd7042
; 
32'd166974: dataIn1 = 32'd7049
; 
32'd166975: dataIn1 = 32'd5873
; 
32'd166976: dataIn1 = 32'd5879
; 
32'd166977: dataIn1 = 32'd6992
; 
32'd166978: dataIn1 = 32'd7010
; 
32'd166979: dataIn1 = 32'd7011
; 
32'd166980: dataIn1 = 32'd7012
; 
32'd166981: dataIn1 = 32'd7013
; 
32'd166982: dataIn1 = 32'd5873
; 
32'd166983: dataIn1 = 32'd5878
; 
32'd166984: dataIn1 = 32'd6994
; 
32'd166985: dataIn1 = 32'd7010
; 
32'd166986: dataIn1 = 32'd7011
; 
32'd166987: dataIn1 = 32'd7012
; 
32'd166988: dataIn1 = 32'd7014
; 
32'd166989: dataIn1 = 32'd5878
; 
32'd166990: dataIn1 = 32'd5879
; 
32'd166991: dataIn1 = 32'd7010
; 
32'd166992: dataIn1 = 32'd7011
; 
32'd166993: dataIn1 = 32'd7012
; 
32'd166994: dataIn1 = 32'd7015
; 
32'd166995: dataIn1 = 32'd7016
; 
32'd166996: dataIn1 = 32'd3981
; 
32'd166997: dataIn1 = 32'd5879
; 
32'd166998: dataIn1 = 32'd5880
; 
32'd166999: dataIn1 = 32'd6992
; 
32'd167000: dataIn1 = 32'd7010
; 
32'd167001: dataIn1 = 32'd7013
; 
32'd167002: dataIn1 = 32'd3982
; 
32'd167003: dataIn1 = 32'd5878
; 
32'd167004: dataIn1 = 32'd6994
; 
32'd167005: dataIn1 = 32'd7011
; 
32'd167006: dataIn1 = 32'd7014
; 
32'd167007: dataIn1 = 32'd7022
; 
32'd167008: dataIn1 = 32'd7033
; 
32'd167009: dataIn1 = 32'd2321
; 
32'd167010: dataIn1 = 32'd5834
; 
32'd167011: dataIn1 = 32'd5879
; 
32'd167012: dataIn1 = 32'd7012
; 
32'd167013: dataIn1 = 32'd7015
; 
32'd167014: dataIn1 = 32'd7016
; 
32'd167015: dataIn1 = 32'd2321
; 
32'd167016: dataIn1 = 32'd5878
; 
32'd167017: dataIn1 = 32'd6899
; 
32'd167018: dataIn1 = 32'd7012
; 
32'd167019: dataIn1 = 32'd7015
; 
32'd167020: dataIn1 = 32'd7016
; 
32'd167021: dataIn1 = 32'd7034
; 
32'd167022: dataIn1 = 32'd5882
; 
32'd167023: dataIn1 = 32'd5883
; 
32'd167024: dataIn1 = 32'd7017
; 
32'd167025: dataIn1 = 32'd7018
; 
32'd167026: dataIn1 = 32'd7019
; 
32'd167027: dataIn1 = 32'd7020
; 
32'd167028: dataIn1 = 32'd7021
; 
32'd167029: dataIn1 = 32'd5881
; 
32'd167030: dataIn1 = 32'd5883
; 
32'd167031: dataIn1 = 32'd7017
; 
32'd167032: dataIn1 = 32'd7018
; 
32'd167033: dataIn1 = 32'd7019
; 
32'd167034: dataIn1 = 32'd7022
; 
32'd167035: dataIn1 = 32'd7023
; 
32'd167036: dataIn1 = 32'd5881
; 
32'd167037: dataIn1 = 32'd5882
; 
32'd167038: dataIn1 = 32'd7017
; 
32'd167039: dataIn1 = 32'd7018
; 
32'd167040: dataIn1 = 32'd7019
; 
32'd167041: dataIn1 = 32'd7024
; 
32'd167042: dataIn1 = 32'd7025
; 
32'd167043: dataIn1 = 32'd3968
; 
32'd167044: dataIn1 = 32'd5883
; 
32'd167045: dataIn1 = 32'd6898
; 
32'd167046: dataIn1 = 32'd7017
; 
32'd167047: dataIn1 = 32'd7020
; 
32'd167048: dataIn1 = 32'd7021
; 
32'd167049: dataIn1 = 32'd7032
; 
32'd167050: dataIn1 = 32'd3968
; 
32'd167051: dataIn1 = 32'd5882
; 
32'd167052: dataIn1 = 32'd6891
; 
32'd167053: dataIn1 = 32'd7017
; 
32'd167054: dataIn1 = 32'd7020
; 
32'd167055: dataIn1 = 32'd7021
; 
32'd167056: dataIn1 = 32'd7029
; 
32'd167057: dataIn1 = 32'd3982
; 
32'd167058: dataIn1 = 32'd5883
; 
32'd167059: dataIn1 = 32'd7014
; 
32'd167060: dataIn1 = 32'd7018
; 
32'd167061: dataIn1 = 32'd7022
; 
32'd167062: dataIn1 = 32'd7023
; 
32'd167063: dataIn1 = 32'd7033
; 
32'd167064: dataIn1 = 32'd3982
; 
32'd167065: dataIn1 = 32'd5881
; 
32'd167066: dataIn1 = 32'd7003
; 
32'd167067: dataIn1 = 32'd7018
; 
32'd167068: dataIn1 = 32'd7022
; 
32'd167069: dataIn1 = 32'd7023
; 
32'd167070: dataIn1 = 32'd7027
; 
32'd167071: dataIn1 = 32'd2315
; 
32'd167072: dataIn1 = 32'd5789
; 
32'd167073: dataIn1 = 32'd5882
; 
32'd167074: dataIn1 = 32'd7019
; 
32'd167075: dataIn1 = 32'd7024
; 
32'd167076: dataIn1 = 32'd7025
; 
32'd167077: dataIn1 = 32'd7031
; 
32'd167078: dataIn1 = 32'd2315
; 
32'd167079: dataIn1 = 32'd5794
; 
32'd167080: dataIn1 = 32'd5881
; 
32'd167081: dataIn1 = 32'd7019
; 
32'd167082: dataIn1 = 32'd7024
; 
32'd167083: dataIn1 = 32'd7025
; 
32'd167084: dataIn1 = 32'd7028
; 
32'd167085: dataIn1 = 32'd3947
; 
32'd167086: dataIn1 = 32'd5793
; 
32'd167087: dataIn1 = 32'd5875
; 
32'd167088: dataIn1 = 32'd7001
; 
32'd167089: dataIn1 = 32'd7026
; 
32'd167090: dataIn1 = 32'd7027
; 
32'd167091: dataIn1 = 32'd7028
; 
32'd167092: dataIn1 = 32'd5875
; 
32'd167093: dataIn1 = 32'd5881
; 
32'd167094: dataIn1 = 32'd7003
; 
32'd167095: dataIn1 = 32'd7023
; 
32'd167096: dataIn1 = 32'd7026
; 
32'd167097: dataIn1 = 32'd7027
; 
32'd167098: dataIn1 = 32'd7028
; 
32'd167099: dataIn1 = 32'd3947
; 
32'd167100: dataIn1 = 32'd5794
; 
32'd167101: dataIn1 = 32'd5881
; 
32'd167102: dataIn1 = 32'd7025
; 
32'd167103: dataIn1 = 32'd7026
; 
32'd167104: dataIn1 = 32'd7027
; 
32'd167105: dataIn1 = 32'd7028
; 
32'd167106: dataIn1 = 32'd5841
; 
32'd167107: dataIn1 = 32'd5882
; 
32'd167108: dataIn1 = 32'd6891
; 
32'd167109: dataIn1 = 32'd7021
; 
32'd167110: dataIn1 = 32'd7029
; 
32'd167111: dataIn1 = 32'd7030
; 
32'd167112: dataIn1 = 32'd7031
; 
32'd167113: dataIn1 = 32'd3946
; 
32'd167114: dataIn1 = 32'd5787
; 
32'd167115: dataIn1 = 32'd5841
; 
32'd167116: dataIn1 = 32'd6892
; 
32'd167117: dataIn1 = 32'd7029
; 
32'd167118: dataIn1 = 32'd7030
; 
32'd167119: dataIn1 = 32'd7031
; 
32'd167120: dataIn1 = 32'd3946
; 
32'd167121: dataIn1 = 32'd5789
; 
32'd167122: dataIn1 = 32'd5882
; 
32'd167123: dataIn1 = 32'd7024
; 
32'd167124: dataIn1 = 32'd7029
; 
32'd167125: dataIn1 = 32'd7030
; 
32'd167126: dataIn1 = 32'd7031
; 
32'd167127: dataIn1 = 32'd5842
; 
32'd167128: dataIn1 = 32'd5883
; 
32'd167129: dataIn1 = 32'd6898
; 
32'd167130: dataIn1 = 32'd7020
; 
32'd167131: dataIn1 = 32'd7032
; 
32'd167132: dataIn1 = 32'd7033
; 
32'd167133: dataIn1 = 32'd7034
; 
32'd167134: dataIn1 = 32'd5878
; 
32'd167135: dataIn1 = 32'd5883
; 
32'd167136: dataIn1 = 32'd7014
; 
32'd167137: dataIn1 = 32'd7022
; 
32'd167138: dataIn1 = 32'd7032
; 
32'd167139: dataIn1 = 32'd7033
; 
32'd167140: dataIn1 = 32'd7034
; 
32'd167141: dataIn1 = 32'd5842
; 
32'd167142: dataIn1 = 32'd5878
; 
32'd167143: dataIn1 = 32'd6899
; 
32'd167144: dataIn1 = 32'd7016
; 
32'd167145: dataIn1 = 32'd7032
; 
32'd167146: dataIn1 = 32'd7033
; 
32'd167147: dataIn1 = 32'd7034
; 
32'd167148: dataIn1 = 32'd5885
; 
32'd167149: dataIn1 = 32'd5886
; 
32'd167150: dataIn1 = 32'd7035
; 
32'd167151: dataIn1 = 32'd7036
; 
32'd167152: dataIn1 = 32'd7037
; 
32'd167153: dataIn1 = 32'd7038
; 
32'd167154: dataIn1 = 32'd7039
; 
32'd167155: dataIn1 = 32'd5884
; 
32'd167156: dataIn1 = 32'd5886
; 
32'd167157: dataIn1 = 32'd7035
; 
32'd167158: dataIn1 = 32'd7036
; 
32'd167159: dataIn1 = 32'd7037
; 
32'd167160: dataIn1 = 32'd7040
; 
32'd167161: dataIn1 = 32'd7041
; 
32'd167162: dataIn1 = 32'd5884
; 
32'd167163: dataIn1 = 32'd5885
; 
32'd167164: dataIn1 = 32'd7035
; 
32'd167165: dataIn1 = 32'd7036
; 
32'd167166: dataIn1 = 32'd7037
; 
32'd167167: dataIn1 = 32'd7042
; 
32'd167168: dataIn1 = 32'd7043
; 
32'd167169: dataIn1 = 32'd3985
; 
32'd167170: dataIn1 = 32'd5886
; 
32'd167171: dataIn1 = 32'd7035
; 
32'd167172: dataIn1 = 32'd7038
; 
32'd167173: dataIn1 = 32'd7039
; 
32'd167174: dataIn1 = 32'd7051
; 
32'd167175: dataIn1 = 32'd7054
; 
32'd167176: dataIn1 = 32'd3985
; 
32'd167177: dataIn1 = 32'd5885
; 
32'd167178: dataIn1 = 32'd7035
; 
32'd167179: dataIn1 = 32'd7038
; 
32'd167180: dataIn1 = 32'd7039
; 
32'd167181: dataIn1 = 32'd7047
; 
32'd167182: dataIn1 = 32'd7050
; 
32'd167183: dataIn1 = 32'd2316
; 
32'd167184: dataIn1 = 32'd5825
; 
32'd167185: dataIn1 = 32'd5886
; 
32'd167186: dataIn1 = 32'd7036
; 
32'd167187: dataIn1 = 32'd7040
; 
32'd167188: dataIn1 = 32'd7041
; 
32'd167189: dataIn1 = 32'd7052
; 
32'd167190: dataIn1 = 32'd2316
; 
32'd167191: dataIn1 = 32'd5820
; 
32'd167192: dataIn1 = 32'd5884
; 
32'd167193: dataIn1 = 32'd7036
; 
32'd167194: dataIn1 = 32'd7040
; 
32'd167195: dataIn1 = 32'd7041
; 
32'd167196: dataIn1 = 32'd7045
; 
32'd167197: dataIn1 = 32'd3983
; 
32'd167198: dataIn1 = 32'd5885
; 
32'd167199: dataIn1 = 32'd7009
; 
32'd167200: dataIn1 = 32'd7037
; 
32'd167201: dataIn1 = 32'd7042
; 
32'd167202: dataIn1 = 32'd7043
; 
32'd167203: dataIn1 = 32'd7049
; 
32'd167204: dataIn1 = 32'd3983
; 
32'd167205: dataIn1 = 32'd5884
; 
32'd167206: dataIn1 = 32'd7004
; 
32'd167207: dataIn1 = 32'd7037
; 
32'd167208: dataIn1 = 32'd7042
; 
32'd167209: dataIn1 = 32'd7043
; 
32'd167210: dataIn1 = 32'd7046
; 
32'd167211: dataIn1 = 32'd3954
; 
32'd167212: dataIn1 = 32'd5821
; 
32'd167213: dataIn1 = 32'd5874
; 
32'd167214: dataIn1 = 32'd7002
; 
32'd167215: dataIn1 = 32'd7044
; 
32'd167216: dataIn1 = 32'd7045
; 
32'd167217: dataIn1 = 32'd7046
; 
32'd167218: dataIn1 = 32'd3954
; 
32'd167219: dataIn1 = 32'd5820
; 
32'd167220: dataIn1 = 32'd5884
; 
32'd167221: dataIn1 = 32'd7041
; 
32'd167222: dataIn1 = 32'd7044
; 
32'd167223: dataIn1 = 32'd7045
; 
32'd167224: dataIn1 = 32'd7046
; 
32'd167225: dataIn1 = 32'd5874
; 
32'd167226: dataIn1 = 32'd5884
; 
32'd167227: dataIn1 = 32'd7004
; 
32'd167228: dataIn1 = 32'd7043
; 
32'd167229: dataIn1 = 32'd7044
; 
32'd167230: dataIn1 = 32'd7045
; 
32'd167231: dataIn1 = 32'd7046
; 
32'd167232: dataIn1 = 32'd5885
; 
32'd167233: dataIn1 = 32'd5887
; 
32'd167234: dataIn1 = 32'd7039
; 
32'd167235: dataIn1 = 32'd7047
; 
32'd167236: dataIn1 = 32'd7048
; 
32'd167237: dataIn1 = 32'd7049
; 
32'd167238: dataIn1 = 32'd7050
; 
32'd167239: dataIn1 = 32'd2325
; 
32'd167240: dataIn1 = 32'd5876
; 
32'd167241: dataIn1 = 32'd5887
; 
32'd167242: dataIn1 = 32'd7047
; 
32'd167243: dataIn1 = 32'd7048
; 
32'd167244: dataIn1 = 32'd7049
; 
32'd167245: dataIn1 = 32'd5876
; 
32'd167246: dataIn1 = 32'd5885
; 
32'd167247: dataIn1 = 32'd7009
; 
32'd167248: dataIn1 = 32'd7042
; 
32'd167249: dataIn1 = 32'd7047
; 
32'd167250: dataIn1 = 32'd7048
; 
32'd167251: dataIn1 = 32'd7049
; 
32'd167252: dataIn1 = 32'd3985
; 
32'd167253: dataIn1 = 32'd5887
; 
32'd167254: dataIn1 = 32'd7039
; 
32'd167255: dataIn1 = 32'd7047
; 
32'd167256: dataIn1 = 32'd7050
; 
32'd167257: dataIn1 = 32'd9768
; 
32'd167258: dataIn1 = 32'd9779
; 
32'd167259: dataIn1 = 32'd5886
; 
32'd167260: dataIn1 = 32'd5888
; 
32'd167261: dataIn1 = 32'd7038
; 
32'd167262: dataIn1 = 32'd7051
; 
32'd167263: dataIn1 = 32'd7052
; 
32'd167264: dataIn1 = 32'd7053
; 
32'd167265: dataIn1 = 32'd7054
; 
32'd167266: dataIn1 = 32'd3955
; 
32'd167267: dataIn1 = 32'd5825
; 
32'd167268: dataIn1 = 32'd5886
; 
32'd167269: dataIn1 = 32'd7040
; 
32'd167270: dataIn1 = 32'd7051
; 
32'd167271: dataIn1 = 32'd7052
; 
32'd167272: dataIn1 = 32'd7053
; 
32'd167273: dataIn1 = 32'd3955
; 
32'd167274: dataIn1 = 32'd5826
; 
32'd167275: dataIn1 = 32'd5888
; 
32'd167276: dataIn1 = 32'd7051
; 
32'd167277: dataIn1 = 32'd7052
; 
32'd167278: dataIn1 = 32'd7053
; 
32'd167279: dataIn1 = 32'd8925
; 
32'd167280: dataIn1 = 32'd3985
; 
32'd167281: dataIn1 = 32'd5888
; 
32'd167282: dataIn1 = 32'd7038
; 
32'd167283: dataIn1 = 32'd7051
; 
32'd167284: dataIn1 = 32'd7054
; 
32'd167285: dataIn1 = 32'd8923
; 
32'd167286: dataIn1 = 32'd8926
; 
32'd167287: dataIn1 = 32'd6068
; 
32'd167288: dataIn1 = 32'd6069
; 
32'd167289: dataIn1 = 32'd7055
; 
32'd167290: dataIn1 = 32'd7056
; 
32'd167291: dataIn1 = 32'd7057
; 
32'd167292: dataIn1 = 32'd7058
; 
32'd167293: dataIn1 = 32'd7059
; 
32'd167294: dataIn1 = 32'd6067
; 
32'd167295: dataIn1 = 32'd6069
; 
32'd167296: dataIn1 = 32'd7055
; 
32'd167297: dataIn1 = 32'd7056
; 
32'd167298: dataIn1 = 32'd7057
; 
32'd167299: dataIn1 = 32'd7060
; 
32'd167300: dataIn1 = 32'd7061
; 
32'd167301: dataIn1 = 32'd6067
; 
32'd167302: dataIn1 = 32'd6068
; 
32'd167303: dataIn1 = 32'd7055
; 
32'd167304: dataIn1 = 32'd7056
; 
32'd167305: dataIn1 = 32'd7057
; 
32'd167306: dataIn1 = 32'd7062
; 
32'd167307: dataIn1 = 32'd7063
; 
32'd167308: dataIn1 = 32'd5112
; 
32'd167309: dataIn1 = 32'd6069
; 
32'd167310: dataIn1 = 32'd7055
; 
32'd167311: dataIn1 = 32'd7058
; 
32'd167312: dataIn1 = 32'd7059
; 
32'd167313: dataIn1 = 32'd7071
; 
32'd167314: dataIn1 = 32'd7074
; 
32'd167315: dataIn1 = 32'd5112
; 
32'd167316: dataIn1 = 32'd6068
; 
32'd167317: dataIn1 = 32'd6073
; 
32'd167318: dataIn1 = 32'd7055
; 
32'd167319: dataIn1 = 32'd7058
; 
32'd167320: dataIn1 = 32'd7059
; 
32'd167321: dataIn1 = 32'd5113
; 
32'd167322: dataIn1 = 32'd6069
; 
32'd167323: dataIn1 = 32'd7056
; 
32'd167324: dataIn1 = 32'd7060
; 
32'd167325: dataIn1 = 32'd7061
; 
32'd167326: dataIn1 = 32'd7072
; 
32'd167327: dataIn1 = 32'd7075
; 
32'd167328: dataIn1 = 32'd5113
; 
32'd167329: dataIn1 = 32'd6067
; 
32'd167330: dataIn1 = 32'd7056
; 
32'd167331: dataIn1 = 32'd7060
; 
32'd167332: dataIn1 = 32'd7061
; 
32'd167333: dataIn1 = 32'd7065
; 
32'd167334: dataIn1 = 32'd7069
; 
32'd167335: dataIn1 = 32'd5114
; 
32'd167336: dataIn1 = 32'd6068
; 
32'd167337: dataIn1 = 32'd6072
; 
32'd167338: dataIn1 = 32'd7057
; 
32'd167339: dataIn1 = 32'd7062
; 
32'd167340: dataIn1 = 32'd7063
; 
32'd167341: dataIn1 = 32'd5114
; 
32'd167342: dataIn1 = 32'd6067
; 
32'd167343: dataIn1 = 32'd7057
; 
32'd167344: dataIn1 = 32'd7062
; 
32'd167345: dataIn1 = 32'd7063
; 
32'd167346: dataIn1 = 32'd7066
; 
32'd167347: dataIn1 = 32'd7070
; 
32'd167348: dataIn1 = 32'd6070
; 
32'd167349: dataIn1 = 32'd6071
; 
32'd167350: dataIn1 = 32'd7064
; 
32'd167351: dataIn1 = 32'd7065
; 
32'd167352: dataIn1 = 32'd7066
; 
32'd167353: dataIn1 = 32'd7067
; 
32'd167354: dataIn1 = 32'd7068
; 
32'd167355: dataIn1 = 32'd6067
; 
32'd167356: dataIn1 = 32'd6071
; 
32'd167357: dataIn1 = 32'd7061
; 
32'd167358: dataIn1 = 32'd7064
; 
32'd167359: dataIn1 = 32'd7065
; 
32'd167360: dataIn1 = 32'd7066
; 
32'd167361: dataIn1 = 32'd7069
; 
32'd167362: dataIn1 = 32'd6067
; 
32'd167363: dataIn1 = 32'd6070
; 
32'd167364: dataIn1 = 32'd7063
; 
32'd167365: dataIn1 = 32'd7064
; 
32'd167366: dataIn1 = 32'd7065
; 
32'd167367: dataIn1 = 32'd7066
; 
32'd167368: dataIn1 = 32'd7070
; 
32'd167369: dataIn1 = 32'd2692
; 
32'd167370: dataIn1 = 32'd6071
; 
32'd167371: dataIn1 = 32'd7064
; 
32'd167372: dataIn1 = 32'd7067
; 
32'd167373: dataIn1 = 32'd7068
; 
32'd167374: dataIn1 = 32'd7094
; 
32'd167375: dataIn1 = 32'd7097
; 
32'd167376: dataIn1 = 32'd2692
; 
32'd167377: dataIn1 = 32'd6070
; 
32'd167378: dataIn1 = 32'd7064
; 
32'd167379: dataIn1 = 32'd7067
; 
32'd167380: dataIn1 = 32'd7068
; 
32'd167381: dataIn1 = 32'd7104
; 
32'd167382: dataIn1 = 32'd7107
; 
32'd167383: dataIn1 = 32'd5113
; 
32'd167384: dataIn1 = 32'd6071
; 
32'd167385: dataIn1 = 32'd7061
; 
32'd167386: dataIn1 = 32'd7065
; 
32'd167387: dataIn1 = 32'd7069
; 
32'd167388: dataIn1 = 32'd7091
; 
32'd167389: dataIn1 = 32'd7095
; 
32'd167390: dataIn1 = 32'd5114
; 
32'd167391: dataIn1 = 32'd6070
; 
32'd167392: dataIn1 = 32'd7063
; 
32'd167393: dataIn1 = 32'd7066
; 
32'd167394: dataIn1 = 32'd7070
; 
32'd167395: dataIn1 = 32'd7106
; 
32'd167396: dataIn1 = 32'd7110
; 
32'd167397: dataIn1 = 32'd6069
; 
32'd167398: dataIn1 = 32'd6075
; 
32'd167399: dataIn1 = 32'd7058
; 
32'd167400: dataIn1 = 32'd7071
; 
32'd167401: dataIn1 = 32'd7072
; 
32'd167402: dataIn1 = 32'd7073
; 
32'd167403: dataIn1 = 32'd7074
; 
32'd167404: dataIn1 = 32'd6069
; 
32'd167405: dataIn1 = 32'd6074
; 
32'd167406: dataIn1 = 32'd7060
; 
32'd167407: dataIn1 = 32'd7071
; 
32'd167408: dataIn1 = 32'd7072
; 
32'd167409: dataIn1 = 32'd7073
; 
32'd167410: dataIn1 = 32'd7075
; 
32'd167411: dataIn1 = 32'd6074
; 
32'd167412: dataIn1 = 32'd6075
; 
32'd167413: dataIn1 = 32'd7071
; 
32'd167414: dataIn1 = 32'd7072
; 
32'd167415: dataIn1 = 32'd7073
; 
32'd167416: dataIn1 = 32'd7076
; 
32'd167417: dataIn1 = 32'd7077
; 
32'd167418: dataIn1 = 32'd5112
; 
32'd167419: dataIn1 = 32'd6075
; 
32'd167420: dataIn1 = 32'd7058
; 
32'd167421: dataIn1 = 32'd7071
; 
32'd167422: dataIn1 = 32'd7074
; 
32'd167423: dataIn1 = 32'd7078
; 
32'd167424: dataIn1 = 32'd7081
; 
32'd167425: dataIn1 = 32'd5113
; 
32'd167426: dataIn1 = 32'd6074
; 
32'd167427: dataIn1 = 32'd7060
; 
32'd167428: dataIn1 = 32'd7072
; 
32'd167429: dataIn1 = 32'd7075
; 
32'd167430: dataIn1 = 32'd7090
; 
32'd167431: dataIn1 = 32'd7100
; 
32'd167432: dataIn1 = 32'd2694
; 
32'd167433: dataIn1 = 32'd6075
; 
32'd167434: dataIn1 = 32'd7073
; 
32'd167435: dataIn1 = 32'd7076
; 
32'd167436: dataIn1 = 32'd7077
; 
32'd167437: dataIn1 = 32'd7080
; 
32'd167438: dataIn1 = 32'd7084
; 
32'd167439: dataIn1 = 32'd2694
; 
32'd167440: dataIn1 = 32'd6074
; 
32'd167441: dataIn1 = 32'd7073
; 
32'd167442: dataIn1 = 32'd7076
; 
32'd167443: dataIn1 = 32'd7077
; 
32'd167444: dataIn1 = 32'd7101
; 
32'd167445: dataIn1 = 32'd7103
; 
32'd167446: dataIn1 = 32'd6075
; 
32'd167447: dataIn1 = 32'd6078
; 
32'd167448: dataIn1 = 32'd7074
; 
32'd167449: dataIn1 = 32'd7078
; 
32'd167450: dataIn1 = 32'd7079
; 
32'd167451: dataIn1 = 32'd7080
; 
32'd167452: dataIn1 = 32'd7081
; 
32'd167453: dataIn1 = 32'd6078
; 
32'd167454: dataIn1 = 32'd6082
; 
32'd167455: dataIn1 = 32'd7078
; 
32'd167456: dataIn1 = 32'd7079
; 
32'd167457: dataIn1 = 32'd7080
; 
32'd167458: dataIn1 = 32'd7082
; 
32'd167459: dataIn1 = 32'd7083
; 
32'd167460: dataIn1 = 32'd6075
; 
32'd167461: dataIn1 = 32'd6082
; 
32'd167462: dataIn1 = 32'd7076
; 
32'd167463: dataIn1 = 32'd7078
; 
32'd167464: dataIn1 = 32'd7079
; 
32'd167465: dataIn1 = 32'd7080
; 
32'd167466: dataIn1 = 32'd7084
; 
32'd167467: dataIn1 = 32'd5112
; 
32'd167468: dataIn1 = 32'd6077
; 
32'd167469: dataIn1 = 32'd6078
; 
32'd167470: dataIn1 = 32'd7074
; 
32'd167471: dataIn1 = 32'd7078
; 
32'd167472: dataIn1 = 32'd7081
; 
32'd167473: dataIn1 = 32'd5115
; 
32'd167474: dataIn1 = 32'd6076
; 
32'd167475: dataIn1 = 32'd6078
; 
32'd167476: dataIn1 = 32'd7079
; 
32'd167477: dataIn1 = 32'd7082
; 
32'd167478: dataIn1 = 32'd7083
; 
32'd167479: dataIn1 = 32'd5115
; 
32'd167480: dataIn1 = 32'd6082
; 
32'd167481: dataIn1 = 32'd7079
; 
32'd167482: dataIn1 = 32'd7082
; 
32'd167483: dataIn1 = 32'd7083
; 
32'd167484: dataIn1 = 32'd7191
; 
32'd167485: dataIn1 = 32'd7201
; 
32'd167486: dataIn1 = 32'd2694
; 
32'd167487: dataIn1 = 32'd6082
; 
32'd167488: dataIn1 = 32'd7076
; 
32'd167489: dataIn1 = 32'd7080
; 
32'd167490: dataIn1 = 32'd7084
; 
32'd167491: dataIn1 = 32'd7184
; 
32'd167492: dataIn1 = 32'd7202
; 
32'd167493: dataIn1 = 32'd6084
; 
32'd167494: dataIn1 = 32'd6085
; 
32'd167495: dataIn1 = 32'd7085
; 
32'd167496: dataIn1 = 32'd7086
; 
32'd167497: dataIn1 = 32'd7087
; 
32'd167498: dataIn1 = 32'd7088
; 
32'd167499: dataIn1 = 32'd7089
; 
32'd167500: dataIn1 = 32'd6083
; 
32'd167501: dataIn1 = 32'd6085
; 
32'd167502: dataIn1 = 32'd7085
; 
32'd167503: dataIn1 = 32'd7086
; 
32'd167504: dataIn1 = 32'd7087
; 
32'd167505: dataIn1 = 32'd7090
; 
32'd167506: dataIn1 = 32'd7091
; 
32'd167507: dataIn1 = 32'd6083
; 
32'd167508: dataIn1 = 32'd6084
; 
32'd167509: dataIn1 = 32'd7085
; 
32'd167510: dataIn1 = 32'd7086
; 
32'd167511: dataIn1 = 32'd7087
; 
32'd167512: dataIn1 = 32'd7092
; 
32'd167513: dataIn1 = 32'd7093
; 
32'd167514: dataIn1 = 32'd5117
; 
32'd167515: dataIn1 = 32'd6085
; 
32'd167516: dataIn1 = 32'd7085
; 
32'd167517: dataIn1 = 32'd7088
; 
32'd167518: dataIn1 = 32'd7089
; 
32'd167519: dataIn1 = 32'd7099
; 
32'd167520: dataIn1 = 32'd7102
; 
32'd167521: dataIn1 = 32'd5117
; 
32'd167522: dataIn1 = 32'd6084
; 
32'd167523: dataIn1 = 32'd7085
; 
32'd167524: dataIn1 = 32'd7088
; 
32'd167525: dataIn1 = 32'd7089
; 
32'd167526: dataIn1 = 32'd9791
; 
32'd167527: dataIn1 = 32'd9792
; 
32'd167528: dataIn1 = 32'd5113
; 
32'd167529: dataIn1 = 32'd6085
; 
32'd167530: dataIn1 = 32'd7075
; 
32'd167531: dataIn1 = 32'd7086
; 
32'd167532: dataIn1 = 32'd7090
; 
32'd167533: dataIn1 = 32'd7091
; 
32'd167534: dataIn1 = 32'd7100
; 
32'd167535: dataIn1 = 32'd5113
; 
32'd167536: dataIn1 = 32'd6083
; 
32'd167537: dataIn1 = 32'd7069
; 
32'd167538: dataIn1 = 32'd7086
; 
32'd167539: dataIn1 = 32'd7090
; 
32'd167540: dataIn1 = 32'd7091
; 
32'd167541: dataIn1 = 32'd7095
; 
32'd167542: dataIn1 = 32'd5118
; 
32'd167543: dataIn1 = 32'd6084
; 
32'd167544: dataIn1 = 32'd7087
; 
32'd167545: dataIn1 = 32'd7092
; 
32'd167546: dataIn1 = 32'd7093
; 
32'd167547: dataIn1 = 32'd9793
; 
32'd167548: dataIn1 = 32'd9794
; 
32'd167549: dataIn1 = 32'd5118
; 
32'd167550: dataIn1 = 32'd6083
; 
32'd167551: dataIn1 = 32'd7087
; 
32'd167552: dataIn1 = 32'd7092
; 
32'd167553: dataIn1 = 32'd7093
; 
32'd167554: dataIn1 = 32'd7096
; 
32'd167555: dataIn1 = 32'd7098
; 
32'd167556: dataIn1 = 32'd6071
; 
32'd167557: dataIn1 = 32'd6086
; 
32'd167558: dataIn1 = 32'd7067
; 
32'd167559: dataIn1 = 32'd7094
; 
32'd167560: dataIn1 = 32'd7095
; 
32'd167561: dataIn1 = 32'd7096
; 
32'd167562: dataIn1 = 32'd7097
; 
32'd167563: dataIn1 = 32'd6071
; 
32'd167564: dataIn1 = 32'd6083
; 
32'd167565: dataIn1 = 32'd7069
; 
32'd167566: dataIn1 = 32'd7091
; 
32'd167567: dataIn1 = 32'd7094
; 
32'd167568: dataIn1 = 32'd7095
; 
32'd167569: dataIn1 = 32'd7096
; 
32'd167570: dataIn1 = 32'd6083
; 
32'd167571: dataIn1 = 32'd6086
; 
32'd167572: dataIn1 = 32'd7093
; 
32'd167573: dataIn1 = 32'd7094
; 
32'd167574: dataIn1 = 32'd7095
; 
32'd167575: dataIn1 = 32'd7096
; 
32'd167576: dataIn1 = 32'd7098
; 
32'd167577: dataIn1 = 32'd2692
; 
32'd167578: dataIn1 = 32'd6086
; 
32'd167579: dataIn1 = 32'd7067
; 
32'd167580: dataIn1 = 32'd7094
; 
32'd167581: dataIn1 = 32'd7097
; 
32'd167582: dataIn1 = 32'd7123
; 
32'd167583: dataIn1 = 32'd7141
; 
32'd167584: dataIn1 = 32'd5118
; 
32'd167585: dataIn1 = 32'd6086
; 
32'd167586: dataIn1 = 32'd7093
; 
32'd167587: dataIn1 = 32'd7096
; 
32'd167588: dataIn1 = 32'd7098
; 
32'd167589: dataIn1 = 32'd7143
; 
32'd167590: dataIn1 = 32'd7145
; 
32'd167591: dataIn1 = 32'd6085
; 
32'd167592: dataIn1 = 32'd6089
; 
32'd167593: dataIn1 = 32'd7088
; 
32'd167594: dataIn1 = 32'd7099
; 
32'd167595: dataIn1 = 32'd7100
; 
32'd167596: dataIn1 = 32'd7101
; 
32'd167597: dataIn1 = 32'd7102
; 
32'd167598: dataIn1 = 32'd6074
; 
32'd167599: dataIn1 = 32'd6085
; 
32'd167600: dataIn1 = 32'd7075
; 
32'd167601: dataIn1 = 32'd7090
; 
32'd167602: dataIn1 = 32'd7099
; 
32'd167603: dataIn1 = 32'd7100
; 
32'd167604: dataIn1 = 32'd7101
; 
32'd167605: dataIn1 = 32'd6074
; 
32'd167606: dataIn1 = 32'd6089
; 
32'd167607: dataIn1 = 32'd7077
; 
32'd167608: dataIn1 = 32'd7099
; 
32'd167609: dataIn1 = 32'd7100
; 
32'd167610: dataIn1 = 32'd7101
; 
32'd167611: dataIn1 = 32'd7103
; 
32'd167612: dataIn1 = 32'd5117
; 
32'd167613: dataIn1 = 32'd6089
; 
32'd167614: dataIn1 = 32'd7088
; 
32'd167615: dataIn1 = 32'd7099
; 
32'd167616: dataIn1 = 32'd7102
; 
32'd167617: dataIn1 = 32'd7203
; 
32'd167618: dataIn1 = 32'd7206
; 
32'd167619: dataIn1 = 32'd2694
; 
32'd167620: dataIn1 = 32'd6089
; 
32'd167621: dataIn1 = 32'd7077
; 
32'd167622: dataIn1 = 32'd7101
; 
32'd167623: dataIn1 = 32'd7103
; 
32'd167624: dataIn1 = 32'd7185
; 
32'd167625: dataIn1 = 32'd7205
; 
32'd167626: dataIn1 = 32'd6070
; 
32'd167627: dataIn1 = 32'd6093
; 
32'd167628: dataIn1 = 32'd7068
; 
32'd167629: dataIn1 = 32'd7104
; 
32'd167630: dataIn1 = 32'd7105
; 
32'd167631: dataIn1 = 32'd7106
; 
32'd167632: dataIn1 = 32'd7107
; 
32'd167633: dataIn1 = 32'd6090
; 
32'd167634: dataIn1 = 32'd6093
; 
32'd167635: dataIn1 = 32'd7104
; 
32'd167636: dataIn1 = 32'd7105
; 
32'd167637: dataIn1 = 32'd7106
; 
32'd167638: dataIn1 = 32'd7108
; 
32'd167639: dataIn1 = 32'd7109
; 
32'd167640: dataIn1 = 32'd6070
; 
32'd167641: dataIn1 = 32'd6090
; 
32'd167642: dataIn1 = 32'd7070
; 
32'd167643: dataIn1 = 32'd7104
; 
32'd167644: dataIn1 = 32'd7105
; 
32'd167645: dataIn1 = 32'd7106
; 
32'd167646: dataIn1 = 32'd7110
; 
32'd167647: dataIn1 = 32'd2692
; 
32'd167648: dataIn1 = 32'd6093
; 
32'd167649: dataIn1 = 32'd7068
; 
32'd167650: dataIn1 = 32'd7104
; 
32'd167651: dataIn1 = 32'd7107
; 
32'd167652: dataIn1 = 32'd7124
; 
32'd167653: dataIn1 = 32'd7155
; 
32'd167654: dataIn1 = 32'd5120
; 
32'd167655: dataIn1 = 32'd6093
; 
32'd167656: dataIn1 = 32'd7105
; 
32'd167657: dataIn1 = 32'd7108
; 
32'd167658: dataIn1 = 32'd7109
; 
32'd167659: dataIn1 = 32'd7152
; 
32'd167660: dataIn1 = 32'd7156
; 
32'd167661: dataIn1 = 32'd5120
; 
32'd167662: dataIn1 = 32'd6090
; 
32'd167663: dataIn1 = 32'd6092
; 
32'd167664: dataIn1 = 32'd7105
; 
32'd167665: dataIn1 = 32'd7108
; 
32'd167666: dataIn1 = 32'd7109
; 
32'd167667: dataIn1 = 32'd5114
; 
32'd167668: dataIn1 = 32'd6090
; 
32'd167669: dataIn1 = 32'd6091
; 
32'd167670: dataIn1 = 32'd7070
; 
32'd167671: dataIn1 = 32'd7106
; 
32'd167672: dataIn1 = 32'd7110
; 
32'd167673: dataIn1 = 32'd6098
; 
32'd167674: dataIn1 = 32'd6099
; 
32'd167675: dataIn1 = 32'd7111
; 
32'd167676: dataIn1 = 32'd7112
; 
32'd167677: dataIn1 = 32'd7113
; 
32'd167678: dataIn1 = 32'd7114
; 
32'd167679: dataIn1 = 32'd7115
; 
32'd167680: dataIn1 = 32'd6097
; 
32'd167681: dataIn1 = 32'd6099
; 
32'd167682: dataIn1 = 32'd7111
; 
32'd167683: dataIn1 = 32'd7112
; 
32'd167684: dataIn1 = 32'd7113
; 
32'd167685: dataIn1 = 32'd7116
; 
32'd167686: dataIn1 = 32'd7117
; 
32'd167687: dataIn1 = 32'd6097
; 
32'd167688: dataIn1 = 32'd6098
; 
32'd167689: dataIn1 = 32'd7111
; 
32'd167690: dataIn1 = 32'd7112
; 
32'd167691: dataIn1 = 32'd7113
; 
32'd167692: dataIn1 = 32'd7118
; 
32'd167693: dataIn1 = 32'd7119
; 
32'd167694: dataIn1 = 32'd5121
; 
32'd167695: dataIn1 = 32'd6099
; 
32'd167696: dataIn1 = 32'd7111
; 
32'd167697: dataIn1 = 32'd7114
; 
32'd167698: dataIn1 = 32'd7115
; 
32'd167699: dataIn1 = 32'd9801
; 
32'd167700: dataIn1 = 32'd9802
; 
32'd167701: dataIn1 = 32'd5121
; 
32'd167702: dataIn1 = 32'd6098
; 
32'd167703: dataIn1 = 32'd7111
; 
32'd167704: dataIn1 = 32'd7114
; 
32'd167705: dataIn1 = 32'd7115
; 
32'd167706: dataIn1 = 32'd7127
; 
32'd167707: dataIn1 = 32'd7130
; 
32'd167708: dataIn1 = 32'd5122
; 
32'd167709: dataIn1 = 32'd6099
; 
32'd167710: dataIn1 = 32'd7112
; 
32'd167711: dataIn1 = 32'd7116
; 
32'd167712: dataIn1 = 32'd7117
; 
32'd167713: dataIn1 = 32'd9799
; 
32'd167714: dataIn1 = 32'd9800
; 
32'd167715: dataIn1 = 32'd5122
; 
32'd167716: dataIn1 = 32'd6097
; 
32'd167717: dataIn1 = 32'd7112
; 
32'd167718: dataIn1 = 32'd7116
; 
32'd167719: dataIn1 = 32'd7117
; 
32'd167720: dataIn1 = 32'd7121
; 
32'd167721: dataIn1 = 32'd7125
; 
32'd167722: dataIn1 = 32'd5123
; 
32'd167723: dataIn1 = 32'd6098
; 
32'd167724: dataIn1 = 32'd7113
; 
32'd167725: dataIn1 = 32'd7118
; 
32'd167726: dataIn1 = 32'd7119
; 
32'd167727: dataIn1 = 32'd7129
; 
32'd167728: dataIn1 = 32'd7133
; 
32'd167729: dataIn1 = 32'd5123
; 
32'd167730: dataIn1 = 32'd6097
; 
32'd167731: dataIn1 = 32'd7113
; 
32'd167732: dataIn1 = 32'd7118
; 
32'd167733: dataIn1 = 32'd7119
; 
32'd167734: dataIn1 = 32'd7122
; 
32'd167735: dataIn1 = 32'd7126
; 
32'd167736: dataIn1 = 32'd6100
; 
32'd167737: dataIn1 = 32'd6101
; 
32'd167738: dataIn1 = 32'd7120
; 
32'd167739: dataIn1 = 32'd7121
; 
32'd167740: dataIn1 = 32'd7122
; 
32'd167741: dataIn1 = 32'd7123
; 
32'd167742: dataIn1 = 32'd7124
; 
32'd167743: dataIn1 = 32'd6097
; 
32'd167744: dataIn1 = 32'd6101
; 
32'd167745: dataIn1 = 32'd7117
; 
32'd167746: dataIn1 = 32'd7120
; 
32'd167747: dataIn1 = 32'd7121
; 
32'd167748: dataIn1 = 32'd7122
; 
32'd167749: dataIn1 = 32'd7125
; 
32'd167750: dataIn1 = 32'd6097
; 
32'd167751: dataIn1 = 32'd6100
; 
32'd167752: dataIn1 = 32'd7119
; 
32'd167753: dataIn1 = 32'd7120
; 
32'd167754: dataIn1 = 32'd7121
; 
32'd167755: dataIn1 = 32'd7122
; 
32'd167756: dataIn1 = 32'd7126
; 
32'd167757: dataIn1 = 32'd2692
; 
32'd167758: dataIn1 = 32'd6101
; 
32'd167759: dataIn1 = 32'd7097
; 
32'd167760: dataIn1 = 32'd7120
; 
32'd167761: dataIn1 = 32'd7123
; 
32'd167762: dataIn1 = 32'd7124
; 
32'd167763: dataIn1 = 32'd7141
; 
32'd167764: dataIn1 = 32'd2692
; 
32'd167765: dataIn1 = 32'd6100
; 
32'd167766: dataIn1 = 32'd7107
; 
32'd167767: dataIn1 = 32'd7120
; 
32'd167768: dataIn1 = 32'd7123
; 
32'd167769: dataIn1 = 32'd7124
; 
32'd167770: dataIn1 = 32'd7155
; 
32'd167771: dataIn1 = 32'd5122
; 
32'd167772: dataIn1 = 32'd6101
; 
32'd167773: dataIn1 = 32'd7117
; 
32'd167774: dataIn1 = 32'd7121
; 
32'd167775: dataIn1 = 32'd7125
; 
32'd167776: dataIn1 = 32'd7142
; 
32'd167777: dataIn1 = 32'd7144
; 
32'd167778: dataIn1 = 32'd5123
; 
32'd167779: dataIn1 = 32'd6100
; 
32'd167780: dataIn1 = 32'd7119
; 
32'd167781: dataIn1 = 32'd7122
; 
32'd167782: dataIn1 = 32'd7126
; 
32'd167783: dataIn1 = 32'd7154
; 
32'd167784: dataIn1 = 32'd7157
; 
32'd167785: dataIn1 = 32'd6098
; 
32'd167786: dataIn1 = 32'd6103
; 
32'd167787: dataIn1 = 32'd7115
; 
32'd167788: dataIn1 = 32'd7127
; 
32'd167789: dataIn1 = 32'd7128
; 
32'd167790: dataIn1 = 32'd7129
; 
32'd167791: dataIn1 = 32'd7130
; 
32'd167792: dataIn1 = 32'd6102
; 
32'd167793: dataIn1 = 32'd6103
; 
32'd167794: dataIn1 = 32'd7127
; 
32'd167795: dataIn1 = 32'd7128
; 
32'd167796: dataIn1 = 32'd7129
; 
32'd167797: dataIn1 = 32'd7131
; 
32'd167798: dataIn1 = 32'd7132
; 
32'd167799: dataIn1 = 32'd6098
; 
32'd167800: dataIn1 = 32'd6102
; 
32'd167801: dataIn1 = 32'd7118
; 
32'd167802: dataIn1 = 32'd7127
; 
32'd167803: dataIn1 = 32'd7128
; 
32'd167804: dataIn1 = 32'd7129
; 
32'd167805: dataIn1 = 32'd7133
; 
32'd167806: dataIn1 = 32'd5121
; 
32'd167807: dataIn1 = 32'd6103
; 
32'd167808: dataIn1 = 32'd7115
; 
32'd167809: dataIn1 = 32'd7127
; 
32'd167810: dataIn1 = 32'd7130
; 
32'd167811: dataIn1 = 32'd7134
; 
32'd167812: dataIn1 = 32'd7137
; 
32'd167813: dataIn1 = 32'd2695
; 
32'd167814: dataIn1 = 32'd6103
; 
32'd167815: dataIn1 = 32'd7128
; 
32'd167816: dataIn1 = 32'd7131
; 
32'd167817: dataIn1 = 32'd7132
; 
32'd167818: dataIn1 = 32'd7135
; 
32'd167819: dataIn1 = 32'd7138
; 
32'd167820: dataIn1 = 32'd2695
; 
32'd167821: dataIn1 = 32'd6102
; 
32'd167822: dataIn1 = 32'd7128
; 
32'd167823: dataIn1 = 32'd7131
; 
32'd167824: dataIn1 = 32'd7132
; 
32'd167825: dataIn1 = 32'd7159
; 
32'd167826: dataIn1 = 32'd7162
; 
32'd167827: dataIn1 = 32'd5123
; 
32'd167828: dataIn1 = 32'd6102
; 
32'd167829: dataIn1 = 32'd7118
; 
32'd167830: dataIn1 = 32'd7129
; 
32'd167831: dataIn1 = 32'd7133
; 
32'd167832: dataIn1 = 32'd7153
; 
32'd167833: dataIn1 = 32'd7160
; 
32'd167834: dataIn1 = 32'd6103
; 
32'd167835: dataIn1 = 32'd6107
; 
32'd167836: dataIn1 = 32'd7130
; 
32'd167837: dataIn1 = 32'd7134
; 
32'd167838: dataIn1 = 32'd7135
; 
32'd167839: dataIn1 = 32'd7136
; 
32'd167840: dataIn1 = 32'd7137
; 
32'd167841: dataIn1 = 32'd6103
; 
32'd167842: dataIn1 = 32'd6110
; 
32'd167843: dataIn1 = 32'd7131
; 
32'd167844: dataIn1 = 32'd7134
; 
32'd167845: dataIn1 = 32'd7135
; 
32'd167846: dataIn1 = 32'd7136
; 
32'd167847: dataIn1 = 32'd7138
; 
32'd167848: dataIn1 = 32'd6107
; 
32'd167849: dataIn1 = 32'd6110
; 
32'd167850: dataIn1 = 32'd7134
; 
32'd167851: dataIn1 = 32'd7135
; 
32'd167852: dataIn1 = 32'd7136
; 
32'd167853: dataIn1 = 32'd7139
; 
32'd167854: dataIn1 = 32'd7140
; 
32'd167855: dataIn1 = 32'd5121
; 
32'd167856: dataIn1 = 32'd6107
; 
32'd167857: dataIn1 = 32'd7130
; 
32'd167858: dataIn1 = 32'd7134
; 
32'd167859: dataIn1 = 32'd7137
; 
32'd167860: dataIn1 = 32'd9803
; 
32'd167861: dataIn1 = 32'd9804
; 
32'd167862: dataIn1 = 32'd2695
; 
32'd167863: dataIn1 = 32'd6110
; 
32'd167864: dataIn1 = 32'd7131
; 
32'd167865: dataIn1 = 32'd7135
; 
32'd167866: dataIn1 = 32'd7138
; 
32'd167867: dataIn1 = 32'd9361
; 
32'd167868: dataIn1 = 32'd9379
; 
32'd167869: dataIn1 = 32'd5124
; 
32'd167870: dataIn1 = 32'd6107
; 
32'd167871: dataIn1 = 32'd7136
; 
32'd167872: dataIn1 = 32'd7139
; 
32'd167873: dataIn1 = 32'd7140
; 
32'd167874: dataIn1 = 32'd9805
; 
32'd167875: dataIn1 = 32'd9806
; 
32'd167876: dataIn1 = 32'd5124
; 
32'd167877: dataIn1 = 32'd6110
; 
32'd167878: dataIn1 = 32'd7136
; 
32'd167879: dataIn1 = 32'd7139
; 
32'd167880: dataIn1 = 32'd7140
; 
32'd167881: dataIn1 = 32'd9368
; 
32'd167882: dataIn1 = 32'd9378
; 
32'd167883: dataIn1 = 32'd6086
; 
32'd167884: dataIn1 = 32'd6101
; 
32'd167885: dataIn1 = 32'd7097
; 
32'd167886: dataIn1 = 32'd7123
; 
32'd167887: dataIn1 = 32'd7141
; 
32'd167888: dataIn1 = 32'd7142
; 
32'd167889: dataIn1 = 32'd7143
; 
32'd167890: dataIn1 = 32'd6101
; 
32'd167891: dataIn1 = 32'd6111
; 
32'd167892: dataIn1 = 32'd7125
; 
32'd167893: dataIn1 = 32'd7141
; 
32'd167894: dataIn1 = 32'd7142
; 
32'd167895: dataIn1 = 32'd7143
; 
32'd167896: dataIn1 = 32'd7144
; 
32'd167897: dataIn1 = 32'd6086
; 
32'd167898: dataIn1 = 32'd6111
; 
32'd167899: dataIn1 = 32'd7098
; 
32'd167900: dataIn1 = 32'd7141
; 
32'd167901: dataIn1 = 32'd7142
; 
32'd167902: dataIn1 = 32'd7143
; 
32'd167903: dataIn1 = 32'd7145
; 
32'd167904: dataIn1 = 32'd5122
; 
32'd167905: dataIn1 = 32'd6111
; 
32'd167906: dataIn1 = 32'd7125
; 
32'd167907: dataIn1 = 32'd7142
; 
32'd167908: dataIn1 = 32'd7144
; 
32'd167909: dataIn1 = 32'd9797
; 
32'd167910: dataIn1 = 32'd9798
; 
32'd167911: dataIn1 = 32'd5118
; 
32'd167912: dataIn1 = 32'd6111
; 
32'd167913: dataIn1 = 32'd7098
; 
32'd167914: dataIn1 = 32'd7143
; 
32'd167915: dataIn1 = 32'd7145
; 
32'd167916: dataIn1 = 32'd9795
; 
32'd167917: dataIn1 = 32'd9796
; 
32'd167918: dataIn1 = 32'd6115
; 
32'd167919: dataIn1 = 32'd6116
; 
32'd167920: dataIn1 = 32'd7146
; 
32'd167921: dataIn1 = 32'd7147
; 
32'd167922: dataIn1 = 32'd7148
; 
32'd167923: dataIn1 = 32'd7149
; 
32'd167924: dataIn1 = 32'd7150
; 
32'd167925: dataIn1 = 32'd6114
; 
32'd167926: dataIn1 = 32'd6116
; 
32'd167927: dataIn1 = 32'd7146
; 
32'd167928: dataIn1 = 32'd7147
; 
32'd167929: dataIn1 = 32'd7148
; 
32'd167930: dataIn1 = 32'd7151
; 
32'd167931: dataIn1 = 32'd7152
; 
32'd167932: dataIn1 = 32'd6114
; 
32'd167933: dataIn1 = 32'd6115
; 
32'd167934: dataIn1 = 32'd7146
; 
32'd167935: dataIn1 = 32'd7147
; 
32'd167936: dataIn1 = 32'd7148
; 
32'd167937: dataIn1 = 32'd7153
; 
32'd167938: dataIn1 = 32'd7154
; 
32'd167939: dataIn1 = 32'd5125
; 
32'd167940: dataIn1 = 32'd6116
; 
32'd167941: dataIn1 = 32'd6118
; 
32'd167942: dataIn1 = 32'd7146
; 
32'd167943: dataIn1 = 32'd7149
; 
32'd167944: dataIn1 = 32'd7150
; 
32'd167945: dataIn1 = 32'd5125
; 
32'd167946: dataIn1 = 32'd6115
; 
32'd167947: dataIn1 = 32'd7146
; 
32'd167948: dataIn1 = 32'd7149
; 
32'd167949: dataIn1 = 32'd7150
; 
32'd167950: dataIn1 = 32'd7158
; 
32'd167951: dataIn1 = 32'd7161
; 
32'd167952: dataIn1 = 32'd5120
; 
32'd167953: dataIn1 = 32'd6095
; 
32'd167954: dataIn1 = 32'd6116
; 
32'd167955: dataIn1 = 32'd7147
; 
32'd167956: dataIn1 = 32'd7151
; 
32'd167957: dataIn1 = 32'd7152
; 
32'd167958: dataIn1 = 32'd5120
; 
32'd167959: dataIn1 = 32'd6114
; 
32'd167960: dataIn1 = 32'd7108
; 
32'd167961: dataIn1 = 32'd7147
; 
32'd167962: dataIn1 = 32'd7151
; 
32'd167963: dataIn1 = 32'd7152
; 
32'd167964: dataIn1 = 32'd7156
; 
32'd167965: dataIn1 = 32'd5123
; 
32'd167966: dataIn1 = 32'd6115
; 
32'd167967: dataIn1 = 32'd7133
; 
32'd167968: dataIn1 = 32'd7148
; 
32'd167969: dataIn1 = 32'd7153
; 
32'd167970: dataIn1 = 32'd7154
; 
32'd167971: dataIn1 = 32'd7160
; 
32'd167972: dataIn1 = 32'd5123
; 
32'd167973: dataIn1 = 32'd6114
; 
32'd167974: dataIn1 = 32'd7126
; 
32'd167975: dataIn1 = 32'd7148
; 
32'd167976: dataIn1 = 32'd7153
; 
32'd167977: dataIn1 = 32'd7154
; 
32'd167978: dataIn1 = 32'd7157
; 
32'd167979: dataIn1 = 32'd6093
; 
32'd167980: dataIn1 = 32'd6100
; 
32'd167981: dataIn1 = 32'd7107
; 
32'd167982: dataIn1 = 32'd7124
; 
32'd167983: dataIn1 = 32'd7155
; 
32'd167984: dataIn1 = 32'd7156
; 
32'd167985: dataIn1 = 32'd7157
; 
32'd167986: dataIn1 = 32'd6093
; 
32'd167987: dataIn1 = 32'd6114
; 
32'd167988: dataIn1 = 32'd7108
; 
32'd167989: dataIn1 = 32'd7152
; 
32'd167990: dataIn1 = 32'd7155
; 
32'd167991: dataIn1 = 32'd7156
; 
32'd167992: dataIn1 = 32'd7157
; 
32'd167993: dataIn1 = 32'd6100
; 
32'd167994: dataIn1 = 32'd6114
; 
32'd167995: dataIn1 = 32'd7126
; 
32'd167996: dataIn1 = 32'd7154
; 
32'd167997: dataIn1 = 32'd7155
; 
32'd167998: dataIn1 = 32'd7156
; 
32'd167999: dataIn1 = 32'd7157
; 
32'd168000: dataIn1 = 32'd6115
; 
32'd168001: dataIn1 = 32'd6117
; 
32'd168002: dataIn1 = 32'd7150
; 
32'd168003: dataIn1 = 32'd7158
; 
32'd168004: dataIn1 = 32'd7159
; 
32'd168005: dataIn1 = 32'd7160
; 
32'd168006: dataIn1 = 32'd7161
; 
32'd168007: dataIn1 = 32'd6102
; 
32'd168008: dataIn1 = 32'd6117
; 
32'd168009: dataIn1 = 32'd7132
; 
32'd168010: dataIn1 = 32'd7158
; 
32'd168011: dataIn1 = 32'd7159
; 
32'd168012: dataIn1 = 32'd7160
; 
32'd168013: dataIn1 = 32'd7162
; 
32'd168014: dataIn1 = 32'd6102
; 
32'd168015: dataIn1 = 32'd6115
; 
32'd168016: dataIn1 = 32'd7133
; 
32'd168017: dataIn1 = 32'd7153
; 
32'd168018: dataIn1 = 32'd7158
; 
32'd168019: dataIn1 = 32'd7159
; 
32'd168020: dataIn1 = 32'd7160
; 
32'd168021: dataIn1 = 32'd5125
; 
32'd168022: dataIn1 = 32'd6117
; 
32'd168023: dataIn1 = 32'd7150
; 
32'd168024: dataIn1 = 32'd7158
; 
32'd168025: dataIn1 = 32'd7161
; 
32'd168026: dataIn1 = 32'd9380
; 
32'd168027: dataIn1 = 32'd9446
; 
32'd168028: dataIn1 = 32'd2695
; 
32'd168029: dataIn1 = 32'd6117
; 
32'd168030: dataIn1 = 32'd7132
; 
32'd168031: dataIn1 = 32'd7159
; 
32'd168032: dataIn1 = 32'd7162
; 
32'd168033: dataIn1 = 32'd9362
; 
32'd168034: dataIn1 = 32'd9382
; 
32'd168035: dataIn1 = 32'd6120
; 
32'd168036: dataIn1 = 32'd6121
; 
32'd168037: dataIn1 = 32'd7163
; 
32'd168038: dataIn1 = 32'd7164
; 
32'd168039: dataIn1 = 32'd7165
; 
32'd168040: dataIn1 = 32'd7166
; 
32'd168041: dataIn1 = 32'd7167
; 
32'd168042: dataIn1 = 32'd6119
; 
32'd168043: dataIn1 = 32'd6121
; 
32'd168044: dataIn1 = 32'd7163
; 
32'd168045: dataIn1 = 32'd7164
; 
32'd168046: dataIn1 = 32'd7165
; 
32'd168047: dataIn1 = 32'd7168
; 
32'd168048: dataIn1 = 32'd7169
; 
32'd168049: dataIn1 = 32'd6119
; 
32'd168050: dataIn1 = 32'd6120
; 
32'd168051: dataIn1 = 32'd7163
; 
32'd168052: dataIn1 = 32'd7164
; 
32'd168053: dataIn1 = 32'd7165
; 
32'd168054: dataIn1 = 32'd7170
; 
32'd168055: dataIn1 = 32'd7171
; 
32'd168056: dataIn1 = 32'd5126
; 
32'd168057: dataIn1 = 32'd6121
; 
32'd168058: dataIn1 = 32'd7163
; 
32'd168059: dataIn1 = 32'd7166
; 
32'd168060: dataIn1 = 32'd7167
; 
32'd168061: dataIn1 = 32'd7179
; 
32'd168062: dataIn1 = 32'd7182
; 
32'd168063: dataIn1 = 32'd5126
; 
32'd168064: dataIn1 = 32'd6120
; 
32'd168065: dataIn1 = 32'd7163
; 
32'd168066: dataIn1 = 32'd7166
; 
32'd168067: dataIn1 = 32'd7167
; 
32'd168068: dataIn1 = 32'd7172
; 
32'd168069: dataIn1 = 32'd7175
; 
32'd168070: dataIn1 = 32'd5127
; 
32'd168071: dataIn1 = 32'd6121
; 
32'd168072: dataIn1 = 32'd7164
; 
32'd168073: dataIn1 = 32'd7168
; 
32'd168074: dataIn1 = 32'd7169
; 
32'd168075: dataIn1 = 32'd7180
; 
32'd168076: dataIn1 = 32'd7183
; 
32'd168077: dataIn1 = 32'd5127
; 
32'd168078: dataIn1 = 32'd6119
; 
32'd168079: dataIn1 = 32'd7164
; 
32'd168080: dataIn1 = 32'd7168
; 
32'd168081: dataIn1 = 32'd7169
; 
32'd168082: dataIn1 = 32'd9785
; 
32'd168083: dataIn1 = 32'd9786
; 
32'd168084: dataIn1 = 32'd5128
; 
32'd168085: dataIn1 = 32'd6120
; 
32'd168086: dataIn1 = 32'd7165
; 
32'd168087: dataIn1 = 32'd7170
; 
32'd168088: dataIn1 = 32'd7171
; 
32'd168089: dataIn1 = 32'd7174
; 
32'd168090: dataIn1 = 32'd7178
; 
32'd168091: dataIn1 = 32'd5128
; 
32'd168092: dataIn1 = 32'd6119
; 
32'd168093: dataIn1 = 32'd7165
; 
32'd168094: dataIn1 = 32'd7170
; 
32'd168095: dataIn1 = 32'd7171
; 
32'd168096: dataIn1 = 32'd9759
; 
32'd168097: dataIn1 = 32'd9777
; 
32'd168098: dataIn1 = 32'd6120
; 
32'd168099: dataIn1 = 32'd6125
; 
32'd168100: dataIn1 = 32'd7167
; 
32'd168101: dataIn1 = 32'd7172
; 
32'd168102: dataIn1 = 32'd7173
; 
32'd168103: dataIn1 = 32'd7174
; 
32'd168104: dataIn1 = 32'd7175
; 
32'd168105: dataIn1 = 32'd6124
; 
32'd168106: dataIn1 = 32'd6125
; 
32'd168107: dataIn1 = 32'd7172
; 
32'd168108: dataIn1 = 32'd7173
; 
32'd168109: dataIn1 = 32'd7174
; 
32'd168110: dataIn1 = 32'd7176
; 
32'd168111: dataIn1 = 32'd7177
; 
32'd168112: dataIn1 = 32'd6120
; 
32'd168113: dataIn1 = 32'd6124
; 
32'd168114: dataIn1 = 32'd7170
; 
32'd168115: dataIn1 = 32'd7172
; 
32'd168116: dataIn1 = 32'd7173
; 
32'd168117: dataIn1 = 32'd7174
; 
32'd168118: dataIn1 = 32'd7178
; 
32'd168119: dataIn1 = 32'd5126
; 
32'd168120: dataIn1 = 32'd6125
; 
32'd168121: dataIn1 = 32'd7167
; 
32'd168122: dataIn1 = 32'd7172
; 
32'd168123: dataIn1 = 32'd7175
; 
32'd168124: dataIn1 = 32'd7190
; 
32'd168125: dataIn1 = 32'd7195
; 
32'd168126: dataIn1 = 32'd2696
; 
32'd168127: dataIn1 = 32'd6125
; 
32'd168128: dataIn1 = 32'd7173
; 
32'd168129: dataIn1 = 32'd7176
; 
32'd168130: dataIn1 = 32'd7177
; 
32'd168131: dataIn1 = 32'd7196
; 
32'd168132: dataIn1 = 32'd7198
; 
32'd168133: dataIn1 = 32'd2696
; 
32'd168134: dataIn1 = 32'd6124
; 
32'd168135: dataIn1 = 32'd7173
; 
32'd168136: dataIn1 = 32'd7176
; 
32'd168137: dataIn1 = 32'd7177
; 
32'd168138: dataIn1 = 32'd7216
; 
32'd168139: dataIn1 = 32'd7219
; 
32'd168140: dataIn1 = 32'd5128
; 
32'd168141: dataIn1 = 32'd6124
; 
32'd168142: dataIn1 = 32'd7170
; 
32'd168143: dataIn1 = 32'd7174
; 
32'd168144: dataIn1 = 32'd7178
; 
32'd168145: dataIn1 = 32'd7213
; 
32'd168146: dataIn1 = 32'd7217
; 
32'd168147: dataIn1 = 32'd6121
; 
32'd168148: dataIn1 = 32'd6127
; 
32'd168149: dataIn1 = 32'd7166
; 
32'd168150: dataIn1 = 32'd7179
; 
32'd168151: dataIn1 = 32'd7180
; 
32'd168152: dataIn1 = 32'd7181
; 
32'd168153: dataIn1 = 32'd7182
; 
32'd168154: dataIn1 = 32'd6121
; 
32'd168155: dataIn1 = 32'd6126
; 
32'd168156: dataIn1 = 32'd7168
; 
32'd168157: dataIn1 = 32'd7179
; 
32'd168158: dataIn1 = 32'd7180
; 
32'd168159: dataIn1 = 32'd7181
; 
32'd168160: dataIn1 = 32'd7183
; 
32'd168161: dataIn1 = 32'd6126
; 
32'd168162: dataIn1 = 32'd6127
; 
32'd168163: dataIn1 = 32'd7179
; 
32'd168164: dataIn1 = 32'd7180
; 
32'd168165: dataIn1 = 32'd7181
; 
32'd168166: dataIn1 = 32'd7184
; 
32'd168167: dataIn1 = 32'd7185
; 
32'd168168: dataIn1 = 32'd5126
; 
32'd168169: dataIn1 = 32'd6127
; 
32'd168170: dataIn1 = 32'd7166
; 
32'd168171: dataIn1 = 32'd7179
; 
32'd168172: dataIn1 = 32'd7182
; 
32'd168173: dataIn1 = 32'd7189
; 
32'd168174: dataIn1 = 32'd7200
; 
32'd168175: dataIn1 = 32'd5127
; 
32'd168176: dataIn1 = 32'd6126
; 
32'd168177: dataIn1 = 32'd7168
; 
32'd168178: dataIn1 = 32'd7180
; 
32'd168179: dataIn1 = 32'd7183
; 
32'd168180: dataIn1 = 32'd7204
; 
32'd168181: dataIn1 = 32'd7207
; 
32'd168182: dataIn1 = 32'd2694
; 
32'd168183: dataIn1 = 32'd6127
; 
32'd168184: dataIn1 = 32'd7084
; 
32'd168185: dataIn1 = 32'd7181
; 
32'd168186: dataIn1 = 32'd7184
; 
32'd168187: dataIn1 = 32'd7185
; 
32'd168188: dataIn1 = 32'd7202
; 
32'd168189: dataIn1 = 32'd2694
; 
32'd168190: dataIn1 = 32'd6126
; 
32'd168191: dataIn1 = 32'd7103
; 
32'd168192: dataIn1 = 32'd7181
; 
32'd168193: dataIn1 = 32'd7184
; 
32'd168194: dataIn1 = 32'd7185
; 
32'd168195: dataIn1 = 32'd7205
; 
32'd168196: dataIn1 = 32'd6129
; 
32'd168197: dataIn1 = 32'd6130
; 
32'd168198: dataIn1 = 32'd7186
; 
32'd168199: dataIn1 = 32'd7187
; 
32'd168200: dataIn1 = 32'd7188
; 
32'd168201: dataIn1 = 32'd7189
; 
32'd168202: dataIn1 = 32'd7190
; 
32'd168203: dataIn1 = 32'd6128
; 
32'd168204: dataIn1 = 32'd6130
; 
32'd168205: dataIn1 = 32'd7186
; 
32'd168206: dataIn1 = 32'd7187
; 
32'd168207: dataIn1 = 32'd7188
; 
32'd168208: dataIn1 = 32'd7191
; 
32'd168209: dataIn1 = 32'd7192
; 
32'd168210: dataIn1 = 32'd6128
; 
32'd168211: dataIn1 = 32'd6129
; 
32'd168212: dataIn1 = 32'd7186
; 
32'd168213: dataIn1 = 32'd7187
; 
32'd168214: dataIn1 = 32'd7188
; 
32'd168215: dataIn1 = 32'd7193
; 
32'd168216: dataIn1 = 32'd7194
; 
32'd168217: dataIn1 = 32'd5126
; 
32'd168218: dataIn1 = 32'd6130
; 
32'd168219: dataIn1 = 32'd7182
; 
32'd168220: dataIn1 = 32'd7186
; 
32'd168221: dataIn1 = 32'd7189
; 
32'd168222: dataIn1 = 32'd7190
; 
32'd168223: dataIn1 = 32'd7200
; 
32'd168224: dataIn1 = 32'd5126
; 
32'd168225: dataIn1 = 32'd6129
; 
32'd168226: dataIn1 = 32'd7175
; 
32'd168227: dataIn1 = 32'd7186
; 
32'd168228: dataIn1 = 32'd7189
; 
32'd168229: dataIn1 = 32'd7190
; 
32'd168230: dataIn1 = 32'd7195
; 
32'd168231: dataIn1 = 32'd5115
; 
32'd168232: dataIn1 = 32'd6130
; 
32'd168233: dataIn1 = 32'd7083
; 
32'd168234: dataIn1 = 32'd7187
; 
32'd168235: dataIn1 = 32'd7191
; 
32'd168236: dataIn1 = 32'd7192
; 
32'd168237: dataIn1 = 32'd7201
; 
32'd168238: dataIn1 = 32'd5115
; 
32'd168239: dataIn1 = 32'd6080
; 
32'd168240: dataIn1 = 32'd6128
; 
32'd168241: dataIn1 = 32'd7187
; 
32'd168242: dataIn1 = 32'd7191
; 
32'd168243: dataIn1 = 32'd7192
; 
32'd168244: dataIn1 = 32'd5129
; 
32'd168245: dataIn1 = 32'd6129
; 
32'd168246: dataIn1 = 32'd7188
; 
32'd168247: dataIn1 = 32'd7193
; 
32'd168248: dataIn1 = 32'd7194
; 
32'd168249: dataIn1 = 32'd7197
; 
32'd168250: dataIn1 = 32'd7199
; 
32'd168251: dataIn1 = 32'd5129
; 
32'd168252: dataIn1 = 32'd6128
; 
32'd168253: dataIn1 = 32'd6131
; 
32'd168254: dataIn1 = 32'd7188
; 
32'd168255: dataIn1 = 32'd7193
; 
32'd168256: dataIn1 = 32'd7194
; 
32'd168257: dataIn1 = 32'd6125
; 
32'd168258: dataIn1 = 32'd6129
; 
32'd168259: dataIn1 = 32'd7175
; 
32'd168260: dataIn1 = 32'd7190
; 
32'd168261: dataIn1 = 32'd7195
; 
32'd168262: dataIn1 = 32'd7196
; 
32'd168263: dataIn1 = 32'd7197
; 
32'd168264: dataIn1 = 32'd6125
; 
32'd168265: dataIn1 = 32'd6132
; 
32'd168266: dataIn1 = 32'd7176
; 
32'd168267: dataIn1 = 32'd7195
; 
32'd168268: dataIn1 = 32'd7196
; 
32'd168269: dataIn1 = 32'd7197
; 
32'd168270: dataIn1 = 32'd7198
; 
32'd168271: dataIn1 = 32'd6129
; 
32'd168272: dataIn1 = 32'd6132
; 
32'd168273: dataIn1 = 32'd7193
; 
32'd168274: dataIn1 = 32'd7195
; 
32'd168275: dataIn1 = 32'd7196
; 
32'd168276: dataIn1 = 32'd7197
; 
32'd168277: dataIn1 = 32'd7199
; 
32'd168278: dataIn1 = 32'd2696
; 
32'd168279: dataIn1 = 32'd6132
; 
32'd168280: dataIn1 = 32'd7176
; 
32'd168281: dataIn1 = 32'd7196
; 
32'd168282: dataIn1 = 32'd7198
; 
32'd168283: dataIn1 = 32'd8884
; 
32'd168284: dataIn1 = 32'd8917
; 
32'd168285: dataIn1 = 32'd5129
; 
32'd168286: dataIn1 = 32'd6132
; 
32'd168287: dataIn1 = 32'd7193
; 
32'd168288: dataIn1 = 32'd7197
; 
32'd168289: dataIn1 = 32'd7199
; 
32'd168290: dataIn1 = 32'd8916
; 
32'd168291: dataIn1 = 32'd8919
; 
32'd168292: dataIn1 = 32'd6127
; 
32'd168293: dataIn1 = 32'd6130
; 
32'd168294: dataIn1 = 32'd7182
; 
32'd168295: dataIn1 = 32'd7189
; 
32'd168296: dataIn1 = 32'd7200
; 
32'd168297: dataIn1 = 32'd7201
; 
32'd168298: dataIn1 = 32'd7202
; 
32'd168299: dataIn1 = 32'd6082
; 
32'd168300: dataIn1 = 32'd6130
; 
32'd168301: dataIn1 = 32'd7083
; 
32'd168302: dataIn1 = 32'd7191
; 
32'd168303: dataIn1 = 32'd7200
; 
32'd168304: dataIn1 = 32'd7201
; 
32'd168305: dataIn1 = 32'd7202
; 
32'd168306: dataIn1 = 32'd6082
; 
32'd168307: dataIn1 = 32'd6127
; 
32'd168308: dataIn1 = 32'd7084
; 
32'd168309: dataIn1 = 32'd7184
; 
32'd168310: dataIn1 = 32'd7200
; 
32'd168311: dataIn1 = 32'd7201
; 
32'd168312: dataIn1 = 32'd7202
; 
32'd168313: dataIn1 = 32'd6089
; 
32'd168314: dataIn1 = 32'd6135
; 
32'd168315: dataIn1 = 32'd7102
; 
32'd168316: dataIn1 = 32'd7203
; 
32'd168317: dataIn1 = 32'd7204
; 
32'd168318: dataIn1 = 32'd7205
; 
32'd168319: dataIn1 = 32'd7206
; 
32'd168320: dataIn1 = 32'd6126
; 
32'd168321: dataIn1 = 32'd6135
; 
32'd168322: dataIn1 = 32'd7183
; 
32'd168323: dataIn1 = 32'd7203
; 
32'd168324: dataIn1 = 32'd7204
; 
32'd168325: dataIn1 = 32'd7205
; 
32'd168326: dataIn1 = 32'd7207
; 
32'd168327: dataIn1 = 32'd6089
; 
32'd168328: dataIn1 = 32'd6126
; 
32'd168329: dataIn1 = 32'd7103
; 
32'd168330: dataIn1 = 32'd7185
; 
32'd168331: dataIn1 = 32'd7203
; 
32'd168332: dataIn1 = 32'd7204
; 
32'd168333: dataIn1 = 32'd7205
; 
32'd168334: dataIn1 = 32'd5117
; 
32'd168335: dataIn1 = 32'd6135
; 
32'd168336: dataIn1 = 32'd7102
; 
32'd168337: dataIn1 = 32'd7203
; 
32'd168338: dataIn1 = 32'd7206
; 
32'd168339: dataIn1 = 32'd9789
; 
32'd168340: dataIn1 = 32'd9790
; 
32'd168341: dataIn1 = 32'd5127
; 
32'd168342: dataIn1 = 32'd6135
; 
32'd168343: dataIn1 = 32'd7183
; 
32'd168344: dataIn1 = 32'd7204
; 
32'd168345: dataIn1 = 32'd7207
; 
32'd168346: dataIn1 = 32'd9787
; 
32'd168347: dataIn1 = 32'd9788
; 
32'd168348: dataIn1 = 32'd6137
; 
32'd168349: dataIn1 = 32'd6138
; 
32'd168350: dataIn1 = 32'd7208
; 
32'd168351: dataIn1 = 32'd7209
; 
32'd168352: dataIn1 = 32'd7210
; 
32'd168353: dataIn1 = 32'd7211
; 
32'd168354: dataIn1 = 32'd7212
; 
32'd168355: dataIn1 = 32'd6136
; 
32'd168356: dataIn1 = 32'd6138
; 
32'd168357: dataIn1 = 32'd7208
; 
32'd168358: dataIn1 = 32'd7209
; 
32'd168359: dataIn1 = 32'd7210
; 
32'd168360: dataIn1 = 32'd9731
; 
32'd168361: dataIn1 = 32'd9758
; 
32'd168362: dataIn1 = 32'd6136
; 
32'd168363: dataIn1 = 32'd6137
; 
32'd168364: dataIn1 = 32'd7208
; 
32'd168365: dataIn1 = 32'd7209
; 
32'd168366: dataIn1 = 32'd7210
; 
32'd168367: dataIn1 = 32'd7213
; 
32'd168368: dataIn1 = 32'd7214
; 
32'd168369: dataIn1 = 32'd5130
; 
32'd168370: dataIn1 = 32'd6138
; 
32'd168371: dataIn1 = 32'd7208
; 
32'd168372: dataIn1 = 32'd7211
; 
32'd168373: dataIn1 = 32'd7212
; 
32'd168374: dataIn1 = 32'd7220
; 
32'd168375: dataIn1 = 32'd7221
; 
32'd168376: dataIn1 = 32'd5130
; 
32'd168377: dataIn1 = 32'd6137
; 
32'd168378: dataIn1 = 32'd7208
; 
32'd168379: dataIn1 = 32'd7211
; 
32'd168380: dataIn1 = 32'd7212
; 
32'd168381: dataIn1 = 32'd7215
; 
32'd168382: dataIn1 = 32'd7218
; 
32'd168383: dataIn1 = 32'd5128
; 
32'd168384: dataIn1 = 32'd6137
; 
32'd168385: dataIn1 = 32'd7178
; 
32'd168386: dataIn1 = 32'd7210
; 
32'd168387: dataIn1 = 32'd7213
; 
32'd168388: dataIn1 = 32'd7214
; 
32'd168389: dataIn1 = 32'd7217
; 
32'd168390: dataIn1 = 32'd5128
; 
32'd168391: dataIn1 = 32'd6136
; 
32'd168392: dataIn1 = 32'd7210
; 
32'd168393: dataIn1 = 32'd7213
; 
32'd168394: dataIn1 = 32'd7214
; 
32'd168395: dataIn1 = 32'd9728
; 
32'd168396: dataIn1 = 32'd9759
; 
32'd168397: dataIn1 = 32'd6137
; 
32'd168398: dataIn1 = 32'd6139
; 
32'd168399: dataIn1 = 32'd7212
; 
32'd168400: dataIn1 = 32'd7215
; 
32'd168401: dataIn1 = 32'd7216
; 
32'd168402: dataIn1 = 32'd7217
; 
32'd168403: dataIn1 = 32'd7218
; 
32'd168404: dataIn1 = 32'd6124
; 
32'd168405: dataIn1 = 32'd6139
; 
32'd168406: dataIn1 = 32'd7177
; 
32'd168407: dataIn1 = 32'd7215
; 
32'd168408: dataIn1 = 32'd7216
; 
32'd168409: dataIn1 = 32'd7217
; 
32'd168410: dataIn1 = 32'd7219
; 
32'd168411: dataIn1 = 32'd6124
; 
32'd168412: dataIn1 = 32'd6137
; 
32'd168413: dataIn1 = 32'd7178
; 
32'd168414: dataIn1 = 32'd7213
; 
32'd168415: dataIn1 = 32'd7215
; 
32'd168416: dataIn1 = 32'd7216
; 
32'd168417: dataIn1 = 32'd7217
; 
32'd168418: dataIn1 = 32'd5130
; 
32'd168419: dataIn1 = 32'd6139
; 
32'd168420: dataIn1 = 32'd7212
; 
32'd168421: dataIn1 = 32'd7215
; 
32'd168422: dataIn1 = 32'd7218
; 
32'd168423: dataIn1 = 32'd8900
; 
32'd168424: dataIn1 = 32'd8907
; 
32'd168425: dataIn1 = 32'd2696
; 
32'd168426: dataIn1 = 32'd6139
; 
32'd168427: dataIn1 = 32'd7177
; 
32'd168428: dataIn1 = 32'd7216
; 
32'd168429: dataIn1 = 32'd7219
; 
32'd168430: dataIn1 = 32'd8883
; 
32'd168431: dataIn1 = 32'd8906
; 
32'd168432: dataIn1 = 32'd4817
; 
32'd168433: dataIn1 = 32'd6138
; 
32'd168434: dataIn1 = 32'd6140
; 
32'd168435: dataIn1 = 32'd7211
; 
32'd168436: dataIn1 = 32'd7220
; 
32'd168437: dataIn1 = 32'd7221
; 
32'd168438: dataIn1 = 32'd5130
; 
32'd168439: dataIn1 = 32'd6140
; 
32'd168440: dataIn1 = 32'd7211
; 
32'd168441: dataIn1 = 32'd7220
; 
32'd168442: dataIn1 = 32'd7221
; 
32'd168443: dataIn1 = 32'd8901
; 
32'd168444: dataIn1 = 32'd8904
; 
32'd168445: dataIn1 = 32'd6147
; 
32'd168446: dataIn1 = 32'd6148
; 
32'd168447: dataIn1 = 32'd7222
; 
32'd168448: dataIn1 = 32'd7223
; 
32'd168449: dataIn1 = 32'd7224
; 
32'd168450: dataIn1 = 32'd7225
; 
32'd168451: dataIn1 = 32'd7226
; 
32'd168452: dataIn1 = 32'd6146
; 
32'd168453: dataIn1 = 32'd6148
; 
32'd168454: dataIn1 = 32'd7222
; 
32'd168455: dataIn1 = 32'd7223
; 
32'd168456: dataIn1 = 32'd7224
; 
32'd168457: dataIn1 = 32'd7227
; 
32'd168458: dataIn1 = 32'd7228
; 
32'd168459: dataIn1 = 32'd6146
; 
32'd168460: dataIn1 = 32'd6147
; 
32'd168461: dataIn1 = 32'd7222
; 
32'd168462: dataIn1 = 32'd7223
; 
32'd168463: dataIn1 = 32'd7224
; 
32'd168464: dataIn1 = 32'd7229
; 
32'd168465: dataIn1 = 32'd7230
; 
32'd168466: dataIn1 = 32'd5136
; 
32'd168467: dataIn1 = 32'd6148
; 
32'd168468: dataIn1 = 32'd7222
; 
32'd168469: dataIn1 = 32'd7225
; 
32'd168470: dataIn1 = 32'd7226
; 
32'd168471: dataIn1 = 32'd7240
; 
32'd168472: dataIn1 = 32'd7243
; 
32'd168473: dataIn1 = 32'd5136
; 
32'd168474: dataIn1 = 32'd6147
; 
32'd168475: dataIn1 = 32'd7222
; 
32'd168476: dataIn1 = 32'd7225
; 
32'd168477: dataIn1 = 32'd7226
; 
32'd168478: dataIn1 = 32'd7233
; 
32'd168479: dataIn1 = 32'd7236
; 
32'd168480: dataIn1 = 32'd5132
; 
32'd168481: dataIn1 = 32'd6148
; 
32'd168482: dataIn1 = 32'd7223
; 
32'd168483: dataIn1 = 32'd7227
; 
32'd168484: dataIn1 = 32'd7228
; 
32'd168485: dataIn1 = 32'd7241
; 
32'd168486: dataIn1 = 32'd7244
; 
32'd168487: dataIn1 = 32'd5132
; 
32'd168488: dataIn1 = 32'd6146
; 
32'd168489: dataIn1 = 32'd6150
; 
32'd168490: dataIn1 = 32'd7223
; 
32'd168491: dataIn1 = 32'd7227
; 
32'd168492: dataIn1 = 32'd7228
; 
32'd168493: dataIn1 = 32'd5137
; 
32'd168494: dataIn1 = 32'd6147
; 
32'd168495: dataIn1 = 32'd7224
; 
32'd168496: dataIn1 = 32'd7229
; 
32'd168497: dataIn1 = 32'd7230
; 
32'd168498: dataIn1 = 32'd7235
; 
32'd168499: dataIn1 = 32'd7239
; 
32'd168500: dataIn1 = 32'd5137
; 
32'd168501: dataIn1 = 32'd6146
; 
32'd168502: dataIn1 = 32'd7224
; 
32'd168503: dataIn1 = 32'd7229
; 
32'd168504: dataIn1 = 32'd7230
; 
32'd168505: dataIn1 = 32'd7231
; 
32'd168506: dataIn1 = 32'd7232
; 
32'd168507: dataIn1 = 32'd5137
; 
32'd168508: dataIn1 = 32'd6149
; 
32'd168509: dataIn1 = 32'd7230
; 
32'd168510: dataIn1 = 32'd7231
; 
32'd168511: dataIn1 = 32'd7232
; 
32'd168512: dataIn1 = 32'd7271
; 
32'd168513: dataIn1 = 32'd7274
; 
32'd168514: dataIn1 = 32'd6146
; 
32'd168515: dataIn1 = 32'd6149
; 
32'd168516: dataIn1 = 32'd6150
; 
32'd168517: dataIn1 = 32'd7230
; 
32'd168518: dataIn1 = 32'd7231
; 
32'd168519: dataIn1 = 32'd7232
; 
32'd168520: dataIn1 = 32'd6147
; 
32'd168521: dataIn1 = 32'd6152
; 
32'd168522: dataIn1 = 32'd7226
; 
32'd168523: dataIn1 = 32'd7233
; 
32'd168524: dataIn1 = 32'd7234
; 
32'd168525: dataIn1 = 32'd7235
; 
32'd168526: dataIn1 = 32'd7236
; 
32'd168527: dataIn1 = 32'd6151
; 
32'd168528: dataIn1 = 32'd6152
; 
32'd168529: dataIn1 = 32'd7233
; 
32'd168530: dataIn1 = 32'd7234
; 
32'd168531: dataIn1 = 32'd7235
; 
32'd168532: dataIn1 = 32'd7237
; 
32'd168533: dataIn1 = 32'd7238
; 
32'd168534: dataIn1 = 32'd6147
; 
32'd168535: dataIn1 = 32'd6151
; 
32'd168536: dataIn1 = 32'd7229
; 
32'd168537: dataIn1 = 32'd7233
; 
32'd168538: dataIn1 = 32'd7234
; 
32'd168539: dataIn1 = 32'd7235
; 
32'd168540: dataIn1 = 32'd7239
; 
32'd168541: dataIn1 = 32'd5136
; 
32'd168542: dataIn1 = 32'd6152
; 
32'd168543: dataIn1 = 32'd7226
; 
32'd168544: dataIn1 = 32'd7233
; 
32'd168545: dataIn1 = 32'd7236
; 
32'd168546: dataIn1 = 32'd7321
; 
32'd168547: dataIn1 = 32'd7329
; 
32'd168548: dataIn1 = 32'd130
; 
32'd168549: dataIn1 = 32'd5972
; 
32'd168550: dataIn1 = 32'd6152
; 
32'd168551: dataIn1 = 32'd7234
; 
32'd168552: dataIn1 = 32'd7237
; 
32'd168553: dataIn1 = 32'd7238
; 
32'd168554: dataIn1 = 32'd7330
; 
32'd168555: dataIn1 = 32'd130
; 
32'd168556: dataIn1 = 32'd6033
; 
32'd168557: dataIn1 = 32'd6151
; 
32'd168558: dataIn1 = 32'd7234
; 
32'd168559: dataIn1 = 32'd7237
; 
32'd168560: dataIn1 = 32'd7238
; 
32'd168561: dataIn1 = 32'd7277
; 
32'd168562: dataIn1 = 32'd5137
; 
32'd168563: dataIn1 = 32'd6151
; 
32'd168564: dataIn1 = 32'd7229
; 
32'd168565: dataIn1 = 32'd7235
; 
32'd168566: dataIn1 = 32'd7239
; 
32'd168567: dataIn1 = 32'd7270
; 
32'd168568: dataIn1 = 32'd7278
; 
32'd168569: dataIn1 = 32'd6148
; 
32'd168570: dataIn1 = 32'd6153
; 
32'd168571: dataIn1 = 32'd7225
; 
32'd168572: dataIn1 = 32'd7240
; 
32'd168573: dataIn1 = 32'd7241
; 
32'd168574: dataIn1 = 32'd7242
; 
32'd168575: dataIn1 = 32'd7243
; 
32'd168576: dataIn1 = 32'd6141
; 
32'd168577: dataIn1 = 32'd6148
; 
32'd168578: dataIn1 = 32'd7227
; 
32'd168579: dataIn1 = 32'd7240
; 
32'd168580: dataIn1 = 32'd7241
; 
32'd168581: dataIn1 = 32'd7242
; 
32'd168582: dataIn1 = 32'd7244
; 
32'd168583: dataIn1 = 32'd6141
; 
32'd168584: dataIn1 = 32'd6153
; 
32'd168585: dataIn1 = 32'd7240
; 
32'd168586: dataIn1 = 32'd7241
; 
32'd168587: dataIn1 = 32'd7242
; 
32'd168588: dataIn1 = 32'd7245
; 
32'd168589: dataIn1 = 32'd7246
; 
32'd168590: dataIn1 = 32'd5136
; 
32'd168591: dataIn1 = 32'd6153
; 
32'd168592: dataIn1 = 32'd7225
; 
32'd168593: dataIn1 = 32'd7240
; 
32'd168594: dataIn1 = 32'd7243
; 
32'd168595: dataIn1 = 32'd7320
; 
32'd168596: dataIn1 = 32'd7332
; 
32'd168597: dataIn1 = 32'd5132
; 
32'd168598: dataIn1 = 32'd6141
; 
32'd168599: dataIn1 = 32'd6143
; 
32'd168600: dataIn1 = 32'd7227
; 
32'd168601: dataIn1 = 32'd7241
; 
32'd168602: dataIn1 = 32'd7244
; 
32'd168603: dataIn1 = 32'd2699
; 
32'd168604: dataIn1 = 32'd6153
; 
32'd168605: dataIn1 = 32'd7242
; 
32'd168606: dataIn1 = 32'd7245
; 
32'd168607: dataIn1 = 32'd7246
; 
32'd168608: dataIn1 = 32'd7311
; 
32'd168609: dataIn1 = 32'd7334
; 
32'd168610: dataIn1 = 32'd2699
; 
32'd168611: dataIn1 = 32'd6141
; 
32'd168612: dataIn1 = 32'd6142
; 
32'd168613: dataIn1 = 32'd7242
; 
32'd168614: dataIn1 = 32'd7245
; 
32'd168615: dataIn1 = 32'd7246
; 
32'd168616: dataIn1 = 32'd6156
; 
32'd168617: dataIn1 = 32'd6160
; 
32'd168618: dataIn1 = 32'd7247
; 
32'd168619: dataIn1 = 32'd7248
; 
32'd168620: dataIn1 = 32'd7249
; 
32'd168621: dataIn1 = 32'd7250
; 
32'd168622: dataIn1 = 32'd7251
; 
32'd168623: dataIn1 = 32'd6156
; 
32'd168624: dataIn1 = 32'd6159
; 
32'd168625: dataIn1 = 32'd7247
; 
32'd168626: dataIn1 = 32'd7248
; 
32'd168627: dataIn1 = 32'd7249
; 
32'd168628: dataIn1 = 32'd7252
; 
32'd168629: dataIn1 = 32'd7253
; 
32'd168630: dataIn1 = 32'd6159
; 
32'd168631: dataIn1 = 32'd6160
; 
32'd168632: dataIn1 = 32'd7247
; 
32'd168633: dataIn1 = 32'd7248
; 
32'd168634: dataIn1 = 32'd7249
; 
32'd168635: dataIn1 = 32'd7254
; 
32'd168636: dataIn1 = 32'd7255
; 
32'd168637: dataIn1 = 32'd5140
; 
32'd168638: dataIn1 = 32'd6156
; 
32'd168639: dataIn1 = 32'd7247
; 
32'd168640: dataIn1 = 32'd7250
; 
32'd168641: dataIn1 = 32'd7251
; 
32'd168642: dataIn1 = 32'd9732
; 
32'd168643: dataIn1 = 32'd9760
; 
32'd168644: dataIn1 = 32'd5140
; 
32'd168645: dataIn1 = 32'd6160
; 
32'd168646: dataIn1 = 32'd7247
; 
32'd168647: dataIn1 = 32'd7250
; 
32'd168648: dataIn1 = 32'd7251
; 
32'd168649: dataIn1 = 32'd7259
; 
32'd168650: dataIn1 = 32'd7262
; 
32'd168651: dataIn1 = 32'd5141
; 
32'd168652: dataIn1 = 32'd6156
; 
32'd168653: dataIn1 = 32'd7248
; 
32'd168654: dataIn1 = 32'd7252
; 
32'd168655: dataIn1 = 32'd7253
; 
32'd168656: dataIn1 = 32'd9733
; 
32'd168657: dataIn1 = 32'd9761
; 
32'd168658: dataIn1 = 32'd5141
; 
32'd168659: dataIn1 = 32'd6159
; 
32'd168660: dataIn1 = 32'd7248
; 
32'd168661: dataIn1 = 32'd7252
; 
32'd168662: dataIn1 = 32'd7253
; 
32'd168663: dataIn1 = 32'd7268
; 
32'd168664: dataIn1 = 32'd7280
; 
32'd168665: dataIn1 = 32'd1106
; 
32'd168666: dataIn1 = 32'd6060
; 
32'd168667: dataIn1 = 32'd6160
; 
32'd168668: dataIn1 = 32'd7249
; 
32'd168669: dataIn1 = 32'd7254
; 
32'd168670: dataIn1 = 32'd7255
; 
32'd168671: dataIn1 = 32'd7261
; 
32'd168672: dataIn1 = 32'd1106
; 
32'd168673: dataIn1 = 32'd6042
; 
32'd168674: dataIn1 = 32'd6159
; 
32'd168675: dataIn1 = 32'd7249
; 
32'd168676: dataIn1 = 32'd7254
; 
32'd168677: dataIn1 = 32'd7255
; 
32'd168678: dataIn1 = 32'd7281
; 
32'd168679: dataIn1 = 32'd4879
; 
32'd168680: dataIn1 = 32'd6055
; 
32'd168681: dataIn1 = 32'd6164
; 
32'd168682: dataIn1 = 32'd7256
; 
32'd168683: dataIn1 = 32'd7257
; 
32'd168684: dataIn1 = 32'd7258
; 
32'd168685: dataIn1 = 32'd8924
; 
32'd168686: dataIn1 = 32'd4879
; 
32'd168687: dataIn1 = 32'd6161
; 
32'd168688: dataIn1 = 32'd6703
; 
32'd168689: dataIn1 = 32'd7256
; 
32'd168690: dataIn1 = 32'd7257
; 
32'd168691: dataIn1 = 32'd7258
; 
32'd168692: dataIn1 = 32'd9232
; 
32'd168693: dataIn1 = 32'd6161
; 
32'd168694: dataIn1 = 32'd6164
; 
32'd168695: dataIn1 = 32'd7256
; 
32'd168696: dataIn1 = 32'd7257
; 
32'd168697: dataIn1 = 32'd7258
; 
32'd168698: dataIn1 = 32'd9767
; 
32'd168699: dataIn1 = 32'd9778
; 
32'd168700: dataIn1 = 32'd6160
; 
32'd168701: dataIn1 = 32'd6163
; 
32'd168702: dataIn1 = 32'd7251
; 
32'd168703: dataIn1 = 32'd7259
; 
32'd168704: dataIn1 = 32'd7260
; 
32'd168705: dataIn1 = 32'd7261
; 
32'd168706: dataIn1 = 32'd7262
; 
32'd168707: dataIn1 = 32'd4880
; 
32'd168708: dataIn1 = 32'd6059
; 
32'd168709: dataIn1 = 32'd6163
; 
32'd168710: dataIn1 = 32'd7259
; 
32'd168711: dataIn1 = 32'd7260
; 
32'd168712: dataIn1 = 32'd7261
; 
32'd168713: dataIn1 = 32'd9274
; 
32'd168714: dataIn1 = 32'd4880
; 
32'd168715: dataIn1 = 32'd6060
; 
32'd168716: dataIn1 = 32'd6160
; 
32'd168717: dataIn1 = 32'd7254
; 
32'd168718: dataIn1 = 32'd7259
; 
32'd168719: dataIn1 = 32'd7260
; 
32'd168720: dataIn1 = 32'd7261
; 
32'd168721: dataIn1 = 32'd5140
; 
32'd168722: dataIn1 = 32'd6163
; 
32'd168723: dataIn1 = 32'd7251
; 
32'd168724: dataIn1 = 32'd7259
; 
32'd168725: dataIn1 = 32'd7262
; 
32'd168726: dataIn1 = 32'd10123
; 
32'd168727: dataIn1 = 32'd10220
; 
32'd168728: dataIn1 = 32'd6166
; 
32'd168729: dataIn1 = 32'd6167
; 
32'd168730: dataIn1 = 32'd7263
; 
32'd168731: dataIn1 = 32'd7264
; 
32'd168732: dataIn1 = 32'd7265
; 
32'd168733: dataIn1 = 32'd7266
; 
32'd168734: dataIn1 = 32'd7267
; 
32'd168735: dataIn1 = 32'd6165
; 
32'd168736: dataIn1 = 32'd6167
; 
32'd168737: dataIn1 = 32'd7263
; 
32'd168738: dataIn1 = 32'd7264
; 
32'd168739: dataIn1 = 32'd7265
; 
32'd168740: dataIn1 = 32'd7268
; 
32'd168741: dataIn1 = 32'd7269
; 
32'd168742: dataIn1 = 32'd6165
; 
32'd168743: dataIn1 = 32'd6166
; 
32'd168744: dataIn1 = 32'd7263
; 
32'd168745: dataIn1 = 32'd7264
; 
32'd168746: dataIn1 = 32'd7265
; 
32'd168747: dataIn1 = 32'd7270
; 
32'd168748: dataIn1 = 32'd7271
; 
32'd168749: dataIn1 = 32'd2630
; 
32'd168750: dataIn1 = 32'd6041
; 
32'd168751: dataIn1 = 32'd6167
; 
32'd168752: dataIn1 = 32'd7263
; 
32'd168753: dataIn1 = 32'd7266
; 
32'd168754: dataIn1 = 32'd7267
; 
32'd168755: dataIn1 = 32'd7279
; 
32'd168756: dataIn1 = 32'd2630
; 
32'd168757: dataIn1 = 32'd6034
; 
32'd168758: dataIn1 = 32'd6166
; 
32'd168759: dataIn1 = 32'd7263
; 
32'd168760: dataIn1 = 32'd7266
; 
32'd168761: dataIn1 = 32'd7267
; 
32'd168762: dataIn1 = 32'd7276
; 
32'd168763: dataIn1 = 32'd5141
; 
32'd168764: dataIn1 = 32'd6167
; 
32'd168765: dataIn1 = 32'd7253
; 
32'd168766: dataIn1 = 32'd7264
; 
32'd168767: dataIn1 = 32'd7268
; 
32'd168768: dataIn1 = 32'd7269
; 
32'd168769: dataIn1 = 32'd7280
; 
32'd168770: dataIn1 = 32'd5141
; 
32'd168771: dataIn1 = 32'd6165
; 
32'd168772: dataIn1 = 32'd7264
; 
32'd168773: dataIn1 = 32'd7268
; 
32'd168774: dataIn1 = 32'd7269
; 
32'd168775: dataIn1 = 32'd7273
; 
32'd168776: dataIn1 = 32'd7275
; 
32'd168777: dataIn1 = 32'd5137
; 
32'd168778: dataIn1 = 32'd6166
; 
32'd168779: dataIn1 = 32'd7239
; 
32'd168780: dataIn1 = 32'd7265
; 
32'd168781: dataIn1 = 32'd7270
; 
32'd168782: dataIn1 = 32'd7271
; 
32'd168783: dataIn1 = 32'd7278
; 
32'd168784: dataIn1 = 32'd5137
; 
32'd168785: dataIn1 = 32'd6165
; 
32'd168786: dataIn1 = 32'd7231
; 
32'd168787: dataIn1 = 32'd7265
; 
32'd168788: dataIn1 = 32'd7270
; 
32'd168789: dataIn1 = 32'd7271
; 
32'd168790: dataIn1 = 32'd7274
; 
32'd168791: dataIn1 = 32'd2697
; 
32'd168792: dataIn1 = 32'd6149
; 
32'd168793: dataIn1 = 32'd6158
; 
32'd168794: dataIn1 = 32'd7272
; 
32'd168795: dataIn1 = 32'd7273
; 
32'd168796: dataIn1 = 32'd7274
; 
32'd168797: dataIn1 = 32'd6158
; 
32'd168798: dataIn1 = 32'd6165
; 
32'd168799: dataIn1 = 32'd7269
; 
32'd168800: dataIn1 = 32'd7272
; 
32'd168801: dataIn1 = 32'd7273
; 
32'd168802: dataIn1 = 32'd7274
; 
32'd168803: dataIn1 = 32'd7275
; 
32'd168804: dataIn1 = 32'd6149
; 
32'd168805: dataIn1 = 32'd6165
; 
32'd168806: dataIn1 = 32'd7231
; 
32'd168807: dataIn1 = 32'd7271
; 
32'd168808: dataIn1 = 32'd7272
; 
32'd168809: dataIn1 = 32'd7273
; 
32'd168810: dataIn1 = 32'd7274
; 
32'd168811: dataIn1 = 32'd5141
; 
32'd168812: dataIn1 = 32'd6158
; 
32'd168813: dataIn1 = 32'd7269
; 
32'd168814: dataIn1 = 32'd7273
; 
32'd168815: dataIn1 = 32'd7275
; 
32'd168816: dataIn1 = 32'd9761
; 
32'd168817: dataIn1 = 32'd9762
; 
32'd168818: dataIn1 = 32'd4874
; 
32'd168819: dataIn1 = 32'd6034
; 
32'd168820: dataIn1 = 32'd6166
; 
32'd168821: dataIn1 = 32'd7267
; 
32'd168822: dataIn1 = 32'd7276
; 
32'd168823: dataIn1 = 32'd7277
; 
32'd168824: dataIn1 = 32'd7278
; 
32'd168825: dataIn1 = 32'd4874
; 
32'd168826: dataIn1 = 32'd6033
; 
32'd168827: dataIn1 = 32'd6151
; 
32'd168828: dataIn1 = 32'd7238
; 
32'd168829: dataIn1 = 32'd7276
; 
32'd168830: dataIn1 = 32'd7277
; 
32'd168831: dataIn1 = 32'd7278
; 
32'd168832: dataIn1 = 32'd6151
; 
32'd168833: dataIn1 = 32'd6166
; 
32'd168834: dataIn1 = 32'd7239
; 
32'd168835: dataIn1 = 32'd7270
; 
32'd168836: dataIn1 = 32'd7276
; 
32'd168837: dataIn1 = 32'd7277
; 
32'd168838: dataIn1 = 32'd7278
; 
32'd168839: dataIn1 = 32'd4875
; 
32'd168840: dataIn1 = 32'd6041
; 
32'd168841: dataIn1 = 32'd6167
; 
32'd168842: dataIn1 = 32'd7266
; 
32'd168843: dataIn1 = 32'd7279
; 
32'd168844: dataIn1 = 32'd7280
; 
32'd168845: dataIn1 = 32'd7281
; 
32'd168846: dataIn1 = 32'd6159
; 
32'd168847: dataIn1 = 32'd6167
; 
32'd168848: dataIn1 = 32'd7253
; 
32'd168849: dataIn1 = 32'd7268
; 
32'd168850: dataIn1 = 32'd7279
; 
32'd168851: dataIn1 = 32'd7280
; 
32'd168852: dataIn1 = 32'd7281
; 
32'd168853: dataIn1 = 32'd4875
; 
32'd168854: dataIn1 = 32'd6042
; 
32'd168855: dataIn1 = 32'd6159
; 
32'd168856: dataIn1 = 32'd7255
; 
32'd168857: dataIn1 = 32'd7279
; 
32'd168858: dataIn1 = 32'd7280
; 
32'd168859: dataIn1 = 32'd7281
; 
32'd168860: dataIn1 = 32'd6169
; 
32'd168861: dataIn1 = 32'd6170
; 
32'd168862: dataIn1 = 32'd7282
; 
32'd168863: dataIn1 = 32'd7283
; 
32'd168864: dataIn1 = 32'd7284
; 
32'd168865: dataIn1 = 32'd7285
; 
32'd168866: dataIn1 = 32'd7286
; 
32'd168867: dataIn1 = 32'd6168
; 
32'd168868: dataIn1 = 32'd6170
; 
32'd168869: dataIn1 = 32'd7282
; 
32'd168870: dataIn1 = 32'd7283
; 
32'd168871: dataIn1 = 32'd7284
; 
32'd168872: dataIn1 = 32'd7287
; 
32'd168873: dataIn1 = 32'd7288
; 
32'd168874: dataIn1 = 32'd6168
; 
32'd168875: dataIn1 = 32'd6169
; 
32'd168876: dataIn1 = 32'd7282
; 
32'd168877: dataIn1 = 32'd7283
; 
32'd168878: dataIn1 = 32'd7284
; 
32'd168879: dataIn1 = 32'd7289
; 
32'd168880: dataIn1 = 32'd7290
; 
32'd168881: dataIn1 = 32'd5145
; 
32'd168882: dataIn1 = 32'd6170
; 
32'd168883: dataIn1 = 32'd7282
; 
32'd168884: dataIn1 = 32'd7285
; 
32'd168885: dataIn1 = 32'd7286
; 
32'd168886: dataIn1 = 32'd7305
; 
32'd168887: dataIn1 = 32'd7308
; 
32'd168888: dataIn1 = 32'd5145
; 
32'd168889: dataIn1 = 32'd6169
; 
32'd168890: dataIn1 = 32'd7282
; 
32'd168891: dataIn1 = 32'd7285
; 
32'd168892: dataIn1 = 32'd7286
; 
32'd168893: dataIn1 = 32'd7298
; 
32'd168894: dataIn1 = 32'd7301
; 
32'd168895: dataIn1 = 32'd5146
; 
32'd168896: dataIn1 = 32'd6170
; 
32'd168897: dataIn1 = 32'd7283
; 
32'd168898: dataIn1 = 32'd7287
; 
32'd168899: dataIn1 = 32'd7288
; 
32'd168900: dataIn1 = 32'd7306
; 
32'd168901: dataIn1 = 32'd7309
; 
32'd168902: dataIn1 = 32'd5146
; 
32'd168903: dataIn1 = 32'd6168
; 
32'd168904: dataIn1 = 32'd7283
; 
32'd168905: dataIn1 = 32'd7287
; 
32'd168906: dataIn1 = 32'd7288
; 
32'd168907: dataIn1 = 32'd7292
; 
32'd168908: dataIn1 = 32'd7296
; 
32'd168909: dataIn1 = 32'd5147
; 
32'd168910: dataIn1 = 32'd6169
; 
32'd168911: dataIn1 = 32'd7284
; 
32'd168912: dataIn1 = 32'd7289
; 
32'd168913: dataIn1 = 32'd7290
; 
32'd168914: dataIn1 = 32'd7300
; 
32'd168915: dataIn1 = 32'd7304
; 
32'd168916: dataIn1 = 32'd5147
; 
32'd168917: dataIn1 = 32'd6168
; 
32'd168918: dataIn1 = 32'd7284
; 
32'd168919: dataIn1 = 32'd7289
; 
32'd168920: dataIn1 = 32'd7290
; 
32'd168921: dataIn1 = 32'd7293
; 
32'd168922: dataIn1 = 32'd7297
; 
32'd168923: dataIn1 = 32'd6171
; 
32'd168924: dataIn1 = 32'd6172
; 
32'd168925: dataIn1 = 32'd7291
; 
32'd168926: dataIn1 = 32'd7292
; 
32'd168927: dataIn1 = 32'd7293
; 
32'd168928: dataIn1 = 32'd7294
; 
32'd168929: dataIn1 = 32'd7295
; 
32'd168930: dataIn1 = 32'd6168
; 
32'd168931: dataIn1 = 32'd6172
; 
32'd168932: dataIn1 = 32'd7288
; 
32'd168933: dataIn1 = 32'd7291
; 
32'd168934: dataIn1 = 32'd7292
; 
32'd168935: dataIn1 = 32'd7293
; 
32'd168936: dataIn1 = 32'd7296
; 
32'd168937: dataIn1 = 32'd6168
; 
32'd168938: dataIn1 = 32'd6171
; 
32'd168939: dataIn1 = 32'd7290
; 
32'd168940: dataIn1 = 32'd7291
; 
32'd168941: dataIn1 = 32'd7292
; 
32'd168942: dataIn1 = 32'd7293
; 
32'd168943: dataIn1 = 32'd7297
; 
32'd168944: dataIn1 = 32'd1105
; 
32'd168945: dataIn1 = 32'd5977
; 
32'd168946: dataIn1 = 32'd6172
; 
32'd168947: dataIn1 = 32'd7291
; 
32'd168948: dataIn1 = 32'd7294
; 
32'd168949: dataIn1 = 32'd7295
; 
32'd168950: dataIn1 = 32'd7326
; 
32'd168951: dataIn1 = 32'd1105
; 
32'd168952: dataIn1 = 32'd5990
; 
32'd168953: dataIn1 = 32'd6171
; 
32'd168954: dataIn1 = 32'd7291
; 
32'd168955: dataIn1 = 32'd7294
; 
32'd168956: dataIn1 = 32'd7295
; 
32'd168957: dataIn1 = 32'd7344
; 
32'd168958: dataIn1 = 32'd5146
; 
32'd168959: dataIn1 = 32'd6172
; 
32'd168960: dataIn1 = 32'd7288
; 
32'd168961: dataIn1 = 32'd7292
; 
32'd168962: dataIn1 = 32'd7296
; 
32'd168963: dataIn1 = 32'd7323
; 
32'd168964: dataIn1 = 32'd7327
; 
32'd168965: dataIn1 = 32'd5147
; 
32'd168966: dataIn1 = 32'd6171
; 
32'd168967: dataIn1 = 32'd7290
; 
32'd168968: dataIn1 = 32'd7293
; 
32'd168969: dataIn1 = 32'd7297
; 
32'd168970: dataIn1 = 32'd7343
; 
32'd168971: dataIn1 = 32'd7346
; 
32'd168972: dataIn1 = 32'd6169
; 
32'd168973: dataIn1 = 32'd6174
; 
32'd168974: dataIn1 = 32'd7286
; 
32'd168975: dataIn1 = 32'd7298
; 
32'd168976: dataIn1 = 32'd7299
; 
32'd168977: dataIn1 = 32'd7300
; 
32'd168978: dataIn1 = 32'd7301
; 
32'd168979: dataIn1 = 32'd6173
; 
32'd168980: dataIn1 = 32'd6174
; 
32'd168981: dataIn1 = 32'd7298
; 
32'd168982: dataIn1 = 32'd7299
; 
32'd168983: dataIn1 = 32'd7300
; 
32'd168984: dataIn1 = 32'd7302
; 
32'd168985: dataIn1 = 32'd7303
; 
32'd168986: dataIn1 = 32'd6169
; 
32'd168987: dataIn1 = 32'd6173
; 
32'd168988: dataIn1 = 32'd7289
; 
32'd168989: dataIn1 = 32'd7298
; 
32'd168990: dataIn1 = 32'd7299
; 
32'd168991: dataIn1 = 32'd7300
; 
32'd168992: dataIn1 = 32'd7304
; 
32'd168993: dataIn1 = 32'd5145
; 
32'd168994: dataIn1 = 32'd6174
; 
32'd168995: dataIn1 = 32'd7286
; 
32'd168996: dataIn1 = 32'd7298
; 
32'd168997: dataIn1 = 32'd7301
; 
32'd168998: dataIn1 = 32'd7312
; 
32'd168999: dataIn1 = 32'd7315
; 
32'd169000: dataIn1 = 32'd2703
; 
32'd169001: dataIn1 = 32'd6174
; 
32'd169002: dataIn1 = 32'd7299
; 
32'd169003: dataIn1 = 32'd7302
; 
32'd169004: dataIn1 = 32'd7303
; 
32'd169005: dataIn1 = 32'd7313
; 
32'd169006: dataIn1 = 32'd7316
; 
32'd169007: dataIn1 = 32'd2703
; 
32'd169008: dataIn1 = 32'd6173
; 
32'd169009: dataIn1 = 32'd7299
; 
32'd169010: dataIn1 = 32'd7302
; 
32'd169011: dataIn1 = 32'd7303
; 
32'd169012: dataIn1 = 32'd7348
; 
32'd169013: dataIn1 = 32'd7351
; 
32'd169014: dataIn1 = 32'd5147
; 
32'd169015: dataIn1 = 32'd6173
; 
32'd169016: dataIn1 = 32'd7289
; 
32'd169017: dataIn1 = 32'd7300
; 
32'd169018: dataIn1 = 32'd7304
; 
32'd169019: dataIn1 = 32'd7342
; 
32'd169020: dataIn1 = 32'd7349
; 
32'd169021: dataIn1 = 32'd6170
; 
32'd169022: dataIn1 = 32'd6176
; 
32'd169023: dataIn1 = 32'd7285
; 
32'd169024: dataIn1 = 32'd7305
; 
32'd169025: dataIn1 = 32'd7306
; 
32'd169026: dataIn1 = 32'd7307
; 
32'd169027: dataIn1 = 32'd7308
; 
32'd169028: dataIn1 = 32'd6170
; 
32'd169029: dataIn1 = 32'd6175
; 
32'd169030: dataIn1 = 32'd7287
; 
32'd169031: dataIn1 = 32'd7305
; 
32'd169032: dataIn1 = 32'd7306
; 
32'd169033: dataIn1 = 32'd7307
; 
32'd169034: dataIn1 = 32'd7309
; 
32'd169035: dataIn1 = 32'd6175
; 
32'd169036: dataIn1 = 32'd6176
; 
32'd169037: dataIn1 = 32'd7305
; 
32'd169038: dataIn1 = 32'd7306
; 
32'd169039: dataIn1 = 32'd7307
; 
32'd169040: dataIn1 = 32'd7310
; 
32'd169041: dataIn1 = 32'd7311
; 
32'd169042: dataIn1 = 32'd5145
; 
32'd169043: dataIn1 = 32'd6176
; 
32'd169044: dataIn1 = 32'd6179
; 
32'd169045: dataIn1 = 32'd7285
; 
32'd169046: dataIn1 = 32'd7305
; 
32'd169047: dataIn1 = 32'd7308
; 
32'd169048: dataIn1 = 32'd5146
; 
32'd169049: dataIn1 = 32'd6175
; 
32'd169050: dataIn1 = 32'd7287
; 
32'd169051: dataIn1 = 32'd7306
; 
32'd169052: dataIn1 = 32'd7309
; 
32'd169053: dataIn1 = 32'd7322
; 
32'd169054: dataIn1 = 32'd7333
; 
32'd169055: dataIn1 = 32'd2699
; 
32'd169056: dataIn1 = 32'd6144
; 
32'd169057: dataIn1 = 32'd6176
; 
32'd169058: dataIn1 = 32'd7307
; 
32'd169059: dataIn1 = 32'd7310
; 
32'd169060: dataIn1 = 32'd7311
; 
32'd169061: dataIn1 = 32'd2699
; 
32'd169062: dataIn1 = 32'd6175
; 
32'd169063: dataIn1 = 32'd7245
; 
32'd169064: dataIn1 = 32'd7307
; 
32'd169065: dataIn1 = 32'd7310
; 
32'd169066: dataIn1 = 32'd7311
; 
32'd169067: dataIn1 = 32'd7334
; 
32'd169068: dataIn1 = 32'd6174
; 
32'd169069: dataIn1 = 32'd6178
; 
32'd169070: dataIn1 = 32'd7301
; 
32'd169071: dataIn1 = 32'd7312
; 
32'd169072: dataIn1 = 32'd7313
; 
32'd169073: dataIn1 = 32'd7314
; 
32'd169074: dataIn1 = 32'd7315
; 
32'd169075: dataIn1 = 32'd6174
; 
32'd169076: dataIn1 = 32'd6180
; 
32'd169077: dataIn1 = 32'd7302
; 
32'd169078: dataIn1 = 32'd7312
; 
32'd169079: dataIn1 = 32'd7313
; 
32'd169080: dataIn1 = 32'd7314
; 
32'd169081: dataIn1 = 32'd7316
; 
32'd169082: dataIn1 = 32'd5148
; 
32'd169083: dataIn1 = 32'd6178
; 
32'd169084: dataIn1 = 32'd6180
; 
32'd169085: dataIn1 = 32'd7312
; 
32'd169086: dataIn1 = 32'd7313
; 
32'd169087: dataIn1 = 32'd7314
; 
32'd169088: dataIn1 = 32'd5145
; 
32'd169089: dataIn1 = 32'd6178
; 
32'd169090: dataIn1 = 32'd6179
; 
32'd169091: dataIn1 = 32'd7301
; 
32'd169092: dataIn1 = 32'd7312
; 
32'd169093: dataIn1 = 32'd7315
; 
32'd169094: dataIn1 = 32'd2703
; 
32'd169095: dataIn1 = 32'd6180
; 
32'd169096: dataIn1 = 32'd7302
; 
32'd169097: dataIn1 = 32'd7313
; 
32'd169098: dataIn1 = 32'd7316
; 
32'd169099: dataIn1 = 32'd8941
; 
32'd169100: dataIn1 = 32'd8975
; 
32'd169101: dataIn1 = 32'd6182
; 
32'd169102: dataIn1 = 32'd6183
; 
32'd169103: dataIn1 = 32'd7317
; 
32'd169104: dataIn1 = 32'd7318
; 
32'd169105: dataIn1 = 32'd7319
; 
32'd169106: dataIn1 = 32'd7320
; 
32'd169107: dataIn1 = 32'd7321
; 
32'd169108: dataIn1 = 32'd6181
; 
32'd169109: dataIn1 = 32'd6183
; 
32'd169110: dataIn1 = 32'd7317
; 
32'd169111: dataIn1 = 32'd7318
; 
32'd169112: dataIn1 = 32'd7319
; 
32'd169113: dataIn1 = 32'd7322
; 
32'd169114: dataIn1 = 32'd7323
; 
32'd169115: dataIn1 = 32'd6181
; 
32'd169116: dataIn1 = 32'd6182
; 
32'd169117: dataIn1 = 32'd7317
; 
32'd169118: dataIn1 = 32'd7318
; 
32'd169119: dataIn1 = 32'd7319
; 
32'd169120: dataIn1 = 32'd7324
; 
32'd169121: dataIn1 = 32'd7325
; 
32'd169122: dataIn1 = 32'd5136
; 
32'd169123: dataIn1 = 32'd6183
; 
32'd169124: dataIn1 = 32'd7243
; 
32'd169125: dataIn1 = 32'd7317
; 
32'd169126: dataIn1 = 32'd7320
; 
32'd169127: dataIn1 = 32'd7321
; 
32'd169128: dataIn1 = 32'd7332
; 
32'd169129: dataIn1 = 32'd5136
; 
32'd169130: dataIn1 = 32'd6182
; 
32'd169131: dataIn1 = 32'd7236
; 
32'd169132: dataIn1 = 32'd7317
; 
32'd169133: dataIn1 = 32'd7320
; 
32'd169134: dataIn1 = 32'd7321
; 
32'd169135: dataIn1 = 32'd7329
; 
32'd169136: dataIn1 = 32'd5146
; 
32'd169137: dataIn1 = 32'd6183
; 
32'd169138: dataIn1 = 32'd7309
; 
32'd169139: dataIn1 = 32'd7318
; 
32'd169140: dataIn1 = 32'd7322
; 
32'd169141: dataIn1 = 32'd7323
; 
32'd169142: dataIn1 = 32'd7333
; 
32'd169143: dataIn1 = 32'd5146
; 
32'd169144: dataIn1 = 32'd6181
; 
32'd169145: dataIn1 = 32'd7296
; 
32'd169146: dataIn1 = 32'd7318
; 
32'd169147: dataIn1 = 32'd7322
; 
32'd169148: dataIn1 = 32'd7323
; 
32'd169149: dataIn1 = 32'd7327
; 
32'd169150: dataIn1 = 32'd2625
; 
32'd169151: dataIn1 = 32'd5973
; 
32'd169152: dataIn1 = 32'd6182
; 
32'd169153: dataIn1 = 32'd7319
; 
32'd169154: dataIn1 = 32'd7324
; 
32'd169155: dataIn1 = 32'd7325
; 
32'd169156: dataIn1 = 32'd7331
; 
32'd169157: dataIn1 = 32'd2625
; 
32'd169158: dataIn1 = 32'd5978
; 
32'd169159: dataIn1 = 32'd6181
; 
32'd169160: dataIn1 = 32'd7319
; 
32'd169161: dataIn1 = 32'd7324
; 
32'd169162: dataIn1 = 32'd7325
; 
32'd169163: dataIn1 = 32'd7328
; 
32'd169164: dataIn1 = 32'd4852
; 
32'd169165: dataIn1 = 32'd5977
; 
32'd169166: dataIn1 = 32'd6172
; 
32'd169167: dataIn1 = 32'd7294
; 
32'd169168: dataIn1 = 32'd7326
; 
32'd169169: dataIn1 = 32'd7327
; 
32'd169170: dataIn1 = 32'd7328
; 
32'd169171: dataIn1 = 32'd6172
; 
32'd169172: dataIn1 = 32'd6181
; 
32'd169173: dataIn1 = 32'd7296
; 
32'd169174: dataIn1 = 32'd7323
; 
32'd169175: dataIn1 = 32'd7326
; 
32'd169176: dataIn1 = 32'd7327
; 
32'd169177: dataIn1 = 32'd7328
; 
32'd169178: dataIn1 = 32'd4852
; 
32'd169179: dataIn1 = 32'd5978
; 
32'd169180: dataIn1 = 32'd6181
; 
32'd169181: dataIn1 = 32'd7325
; 
32'd169182: dataIn1 = 32'd7326
; 
32'd169183: dataIn1 = 32'd7327
; 
32'd169184: dataIn1 = 32'd7328
; 
32'd169185: dataIn1 = 32'd6152
; 
32'd169186: dataIn1 = 32'd6182
; 
32'd169187: dataIn1 = 32'd7236
; 
32'd169188: dataIn1 = 32'd7321
; 
32'd169189: dataIn1 = 32'd7329
; 
32'd169190: dataIn1 = 32'd7330
; 
32'd169191: dataIn1 = 32'd7331
; 
32'd169192: dataIn1 = 32'd4851
; 
32'd169193: dataIn1 = 32'd5972
; 
32'd169194: dataIn1 = 32'd6152
; 
32'd169195: dataIn1 = 32'd7237
; 
32'd169196: dataIn1 = 32'd7329
; 
32'd169197: dataIn1 = 32'd7330
; 
32'd169198: dataIn1 = 32'd7331
; 
32'd169199: dataIn1 = 32'd4851
; 
32'd169200: dataIn1 = 32'd5973
; 
32'd169201: dataIn1 = 32'd6182
; 
32'd169202: dataIn1 = 32'd7324
; 
32'd169203: dataIn1 = 32'd7329
; 
32'd169204: dataIn1 = 32'd7330
; 
32'd169205: dataIn1 = 32'd7331
; 
32'd169206: dataIn1 = 32'd6153
; 
32'd169207: dataIn1 = 32'd6183
; 
32'd169208: dataIn1 = 32'd7243
; 
32'd169209: dataIn1 = 32'd7320
; 
32'd169210: dataIn1 = 32'd7332
; 
32'd169211: dataIn1 = 32'd7333
; 
32'd169212: dataIn1 = 32'd7334
; 
32'd169213: dataIn1 = 32'd6175
; 
32'd169214: dataIn1 = 32'd6183
; 
32'd169215: dataIn1 = 32'd7309
; 
32'd169216: dataIn1 = 32'd7322
; 
32'd169217: dataIn1 = 32'd7332
; 
32'd169218: dataIn1 = 32'd7333
; 
32'd169219: dataIn1 = 32'd7334
; 
32'd169220: dataIn1 = 32'd6153
; 
32'd169221: dataIn1 = 32'd6175
; 
32'd169222: dataIn1 = 32'd7245
; 
32'd169223: dataIn1 = 32'd7311
; 
32'd169224: dataIn1 = 32'd7332
; 
32'd169225: dataIn1 = 32'd7333
; 
32'd169226: dataIn1 = 32'd7334
; 
32'd169227: dataIn1 = 32'd6185
; 
32'd169228: dataIn1 = 32'd6186
; 
32'd169229: dataIn1 = 32'd7335
; 
32'd169230: dataIn1 = 32'd7336
; 
32'd169231: dataIn1 = 32'd7337
; 
32'd169232: dataIn1 = 32'd7338
; 
32'd169233: dataIn1 = 32'd7339
; 
32'd169234: dataIn1 = 32'd6184
; 
32'd169235: dataIn1 = 32'd6186
; 
32'd169236: dataIn1 = 32'd7335
; 
32'd169237: dataIn1 = 32'd7336
; 
32'd169238: dataIn1 = 32'd7337
; 
32'd169239: dataIn1 = 32'd7340
; 
32'd169240: dataIn1 = 32'd7341
; 
32'd169241: dataIn1 = 32'd6184
; 
32'd169242: dataIn1 = 32'd6185
; 
32'd169243: dataIn1 = 32'd7335
; 
32'd169244: dataIn1 = 32'd7336
; 
32'd169245: dataIn1 = 32'd7337
; 
32'd169246: dataIn1 = 32'd7342
; 
32'd169247: dataIn1 = 32'd7343
; 
32'd169248: dataIn1 = 32'd5149
; 
32'd169249: dataIn1 = 32'd6186
; 
32'd169250: dataIn1 = 32'd7335
; 
32'd169251: dataIn1 = 32'd7338
; 
32'd169252: dataIn1 = 32'd7339
; 
32'd169253: dataIn1 = 32'd7352
; 
32'd169254: dataIn1 = 32'd7355
; 
32'd169255: dataIn1 = 32'd5149
; 
32'd169256: dataIn1 = 32'd6185
; 
32'd169257: dataIn1 = 32'd7335
; 
32'd169258: dataIn1 = 32'd7338
; 
32'd169259: dataIn1 = 32'd7339
; 
32'd169260: dataIn1 = 32'd7347
; 
32'd169261: dataIn1 = 32'd7350
; 
32'd169262: dataIn1 = 32'd2626
; 
32'd169263: dataIn1 = 32'd5994
; 
32'd169264: dataIn1 = 32'd6186
; 
32'd169265: dataIn1 = 32'd7336
; 
32'd169266: dataIn1 = 32'd7340
; 
32'd169267: dataIn1 = 32'd7341
; 
32'd169268: dataIn1 = 32'd7353
; 
32'd169269: dataIn1 = 32'd2626
; 
32'd169270: dataIn1 = 32'd5989
; 
32'd169271: dataIn1 = 32'd6184
; 
32'd169272: dataIn1 = 32'd7336
; 
32'd169273: dataIn1 = 32'd7340
; 
32'd169274: dataIn1 = 32'd7341
; 
32'd169275: dataIn1 = 32'd7345
; 
32'd169276: dataIn1 = 32'd5147
; 
32'd169277: dataIn1 = 32'd6185
; 
32'd169278: dataIn1 = 32'd7304
; 
32'd169279: dataIn1 = 32'd7337
; 
32'd169280: dataIn1 = 32'd7342
; 
32'd169281: dataIn1 = 32'd7343
; 
32'd169282: dataIn1 = 32'd7349
; 
32'd169283: dataIn1 = 32'd5147
; 
32'd169284: dataIn1 = 32'd6184
; 
32'd169285: dataIn1 = 32'd7297
; 
32'd169286: dataIn1 = 32'd7337
; 
32'd169287: dataIn1 = 32'd7342
; 
32'd169288: dataIn1 = 32'd7343
; 
32'd169289: dataIn1 = 32'd7346
; 
32'd169290: dataIn1 = 32'd4860
; 
32'd169291: dataIn1 = 32'd5990
; 
32'd169292: dataIn1 = 32'd6171
; 
32'd169293: dataIn1 = 32'd7295
; 
32'd169294: dataIn1 = 32'd7344
; 
32'd169295: dataIn1 = 32'd7345
; 
32'd169296: dataIn1 = 32'd7346
; 
32'd169297: dataIn1 = 32'd4860
; 
32'd169298: dataIn1 = 32'd5989
; 
32'd169299: dataIn1 = 32'd6184
; 
32'd169300: dataIn1 = 32'd7341
; 
32'd169301: dataIn1 = 32'd7344
; 
32'd169302: dataIn1 = 32'd7345
; 
32'd169303: dataIn1 = 32'd7346
; 
32'd169304: dataIn1 = 32'd6171
; 
32'd169305: dataIn1 = 32'd6184
; 
32'd169306: dataIn1 = 32'd7297
; 
32'd169307: dataIn1 = 32'd7343
; 
32'd169308: dataIn1 = 32'd7344
; 
32'd169309: dataIn1 = 32'd7345
; 
32'd169310: dataIn1 = 32'd7346
; 
32'd169311: dataIn1 = 32'd6185
; 
32'd169312: dataIn1 = 32'd6187
; 
32'd169313: dataIn1 = 32'd7339
; 
32'd169314: dataIn1 = 32'd7347
; 
32'd169315: dataIn1 = 32'd7348
; 
32'd169316: dataIn1 = 32'd7349
; 
32'd169317: dataIn1 = 32'd7350
; 
32'd169318: dataIn1 = 32'd6173
; 
32'd169319: dataIn1 = 32'd6187
; 
32'd169320: dataIn1 = 32'd7303
; 
32'd169321: dataIn1 = 32'd7347
; 
32'd169322: dataIn1 = 32'd7348
; 
32'd169323: dataIn1 = 32'd7349
; 
32'd169324: dataIn1 = 32'd7351
; 
32'd169325: dataIn1 = 32'd6173
; 
32'd169326: dataIn1 = 32'd6185
; 
32'd169327: dataIn1 = 32'd7304
; 
32'd169328: dataIn1 = 32'd7342
; 
32'd169329: dataIn1 = 32'd7347
; 
32'd169330: dataIn1 = 32'd7348
; 
32'd169331: dataIn1 = 32'd7349
; 
32'd169332: dataIn1 = 32'd5149
; 
32'd169333: dataIn1 = 32'd6187
; 
32'd169334: dataIn1 = 32'd7339
; 
32'd169335: dataIn1 = 32'd7347
; 
32'd169336: dataIn1 = 32'd7350
; 
32'd169337: dataIn1 = 32'd8957
; 
32'd169338: dataIn1 = 32'd8966
; 
32'd169339: dataIn1 = 32'd2703
; 
32'd169340: dataIn1 = 32'd6187
; 
32'd169341: dataIn1 = 32'd7303
; 
32'd169342: dataIn1 = 32'd7348
; 
32'd169343: dataIn1 = 32'd7351
; 
32'd169344: dataIn1 = 32'd8940
; 
32'd169345: dataIn1 = 32'd8965
; 
32'd169346: dataIn1 = 32'd6186
; 
32'd169347: dataIn1 = 32'd6188
; 
32'd169348: dataIn1 = 32'd7338
; 
32'd169349: dataIn1 = 32'd7352
; 
32'd169350: dataIn1 = 32'd7353
; 
32'd169351: dataIn1 = 32'd7354
; 
32'd169352: dataIn1 = 32'd7355
; 
32'd169353: dataIn1 = 32'd4861
; 
32'd169354: dataIn1 = 32'd5994
; 
32'd169355: dataIn1 = 32'd6186
; 
32'd169356: dataIn1 = 32'd7340
; 
32'd169357: dataIn1 = 32'd7352
; 
32'd169358: dataIn1 = 32'd7353
; 
32'd169359: dataIn1 = 32'd7354
; 
32'd169360: dataIn1 = 32'd4861
; 
32'd169361: dataIn1 = 32'd5995
; 
32'd169362: dataIn1 = 32'd6188
; 
32'd169363: dataIn1 = 32'd7352
; 
32'd169364: dataIn1 = 32'd7353
; 
32'd169365: dataIn1 = 32'd7354
; 
32'd169366: dataIn1 = 32'd8963
; 
32'd169367: dataIn1 = 32'd5149
; 
32'd169368: dataIn1 = 32'd6188
; 
32'd169369: dataIn1 = 32'd7338
; 
32'd169370: dataIn1 = 32'd7352
; 
32'd169371: dataIn1 = 32'd7355
; 
32'd169372: dataIn1 = 32'd8958
; 
32'd169373: dataIn1 = 32'd8961
; 
32'd169374: dataIn1 = 32'd6190
; 
32'd169375: dataIn1 = 32'd6191
; 
32'd169376: dataIn1 = 32'd7356
; 
32'd169377: dataIn1 = 32'd7357
; 
32'd169378: dataIn1 = 32'd7358
; 
32'd169379: dataIn1 = 32'd7359
; 
32'd169380: dataIn1 = 32'd7360
; 
32'd169381: dataIn1 = 32'd6189
; 
32'd169382: dataIn1 = 32'd6191
; 
32'd169383: dataIn1 = 32'd7356
; 
32'd169384: dataIn1 = 32'd7357
; 
32'd169385: dataIn1 = 32'd7358
; 
32'd169386: dataIn1 = 32'd7361
; 
32'd169387: dataIn1 = 32'd7362
; 
32'd169388: dataIn1 = 32'd6189
; 
32'd169389: dataIn1 = 32'd6190
; 
32'd169390: dataIn1 = 32'd7356
; 
32'd169391: dataIn1 = 32'd7357
; 
32'd169392: dataIn1 = 32'd7358
; 
32'd169393: dataIn1 = 32'd7363
; 
32'd169394: dataIn1 = 32'd7364
; 
32'd169395: dataIn1 = 32'd5150
; 
32'd169396: dataIn1 = 32'd6191
; 
32'd169397: dataIn1 = 32'd7356
; 
32'd169398: dataIn1 = 32'd7359
; 
32'd169399: dataIn1 = 32'd7360
; 
32'd169400: dataIn1 = 32'd7372
; 
32'd169401: dataIn1 = 32'd7375
; 
32'd169402: dataIn1 = 32'd5150
; 
32'd169403: dataIn1 = 32'd6190
; 
32'd169404: dataIn1 = 32'd6745
; 
32'd169405: dataIn1 = 32'd7356
; 
32'd169406: dataIn1 = 32'd7359
; 
32'd169407: dataIn1 = 32'd7360
; 
32'd169408: dataIn1 = 32'd5151
; 
32'd169409: dataIn1 = 32'd6191
; 
32'd169410: dataIn1 = 32'd7357
; 
32'd169411: dataIn1 = 32'd7361
; 
32'd169412: dataIn1 = 32'd7362
; 
32'd169413: dataIn1 = 32'd7373
; 
32'd169414: dataIn1 = 32'd7376
; 
32'd169415: dataIn1 = 32'd5151
; 
32'd169416: dataIn1 = 32'd6189
; 
32'd169417: dataIn1 = 32'd7357
; 
32'd169418: dataIn1 = 32'd7361
; 
32'd169419: dataIn1 = 32'd7362
; 
32'd169420: dataIn1 = 32'd7366
; 
32'd169421: dataIn1 = 32'd7370
; 
32'd169422: dataIn1 = 32'd5152
; 
32'd169423: dataIn1 = 32'd6190
; 
32'd169424: dataIn1 = 32'd6744
; 
32'd169425: dataIn1 = 32'd7358
; 
32'd169426: dataIn1 = 32'd7363
; 
32'd169427: dataIn1 = 32'd7364
; 
32'd169428: dataIn1 = 32'd5152
; 
32'd169429: dataIn1 = 32'd6189
; 
32'd169430: dataIn1 = 32'd7358
; 
32'd169431: dataIn1 = 32'd7363
; 
32'd169432: dataIn1 = 32'd7364
; 
32'd169433: dataIn1 = 32'd7367
; 
32'd169434: dataIn1 = 32'd7371
; 
32'd169435: dataIn1 = 32'd6192
; 
32'd169436: dataIn1 = 32'd6193
; 
32'd169437: dataIn1 = 32'd7365
; 
32'd169438: dataIn1 = 32'd7366
; 
32'd169439: dataIn1 = 32'd7367
; 
32'd169440: dataIn1 = 32'd7368
; 
32'd169441: dataIn1 = 32'd7369
; 
32'd169442: dataIn1 = 32'd6189
; 
32'd169443: dataIn1 = 32'd6193
; 
32'd169444: dataIn1 = 32'd7362
; 
32'd169445: dataIn1 = 32'd7365
; 
32'd169446: dataIn1 = 32'd7366
; 
32'd169447: dataIn1 = 32'd7367
; 
32'd169448: dataIn1 = 32'd7370
; 
32'd169449: dataIn1 = 32'd6189
; 
32'd169450: dataIn1 = 32'd6192
; 
32'd169451: dataIn1 = 32'd7364
; 
32'd169452: dataIn1 = 32'd7365
; 
32'd169453: dataIn1 = 32'd7366
; 
32'd169454: dataIn1 = 32'd7367
; 
32'd169455: dataIn1 = 32'd7371
; 
32'd169456: dataIn1 = 32'd2704
; 
32'd169457: dataIn1 = 32'd6193
; 
32'd169458: dataIn1 = 32'd7365
; 
32'd169459: dataIn1 = 32'd7368
; 
32'd169460: dataIn1 = 32'd7369
; 
32'd169461: dataIn1 = 32'd7395
; 
32'd169462: dataIn1 = 32'd7398
; 
32'd169463: dataIn1 = 32'd2704
; 
32'd169464: dataIn1 = 32'd6192
; 
32'd169465: dataIn1 = 32'd7365
; 
32'd169466: dataIn1 = 32'd7368
; 
32'd169467: dataIn1 = 32'd7369
; 
32'd169468: dataIn1 = 32'd7412
; 
32'd169469: dataIn1 = 32'd7415
; 
32'd169470: dataIn1 = 32'd5151
; 
32'd169471: dataIn1 = 32'd6193
; 
32'd169472: dataIn1 = 32'd7362
; 
32'd169473: dataIn1 = 32'd7366
; 
32'd169474: dataIn1 = 32'd7370
; 
32'd169475: dataIn1 = 32'd7392
; 
32'd169476: dataIn1 = 32'd7396
; 
32'd169477: dataIn1 = 32'd5152
; 
32'd169478: dataIn1 = 32'd6192
; 
32'd169479: dataIn1 = 32'd7364
; 
32'd169480: dataIn1 = 32'd7367
; 
32'd169481: dataIn1 = 32'd7371
; 
32'd169482: dataIn1 = 32'd7414
; 
32'd169483: dataIn1 = 32'd7418
; 
32'd169484: dataIn1 = 32'd6191
; 
32'd169485: dataIn1 = 32'd6195
; 
32'd169486: dataIn1 = 32'd7359
; 
32'd169487: dataIn1 = 32'd7372
; 
32'd169488: dataIn1 = 32'd7373
; 
32'd169489: dataIn1 = 32'd7374
; 
32'd169490: dataIn1 = 32'd7375
; 
32'd169491: dataIn1 = 32'd6191
; 
32'd169492: dataIn1 = 32'd6194
; 
32'd169493: dataIn1 = 32'd7361
; 
32'd169494: dataIn1 = 32'd7372
; 
32'd169495: dataIn1 = 32'd7373
; 
32'd169496: dataIn1 = 32'd7374
; 
32'd169497: dataIn1 = 32'd7376
; 
32'd169498: dataIn1 = 32'd6194
; 
32'd169499: dataIn1 = 32'd6195
; 
32'd169500: dataIn1 = 32'd7372
; 
32'd169501: dataIn1 = 32'd7373
; 
32'd169502: dataIn1 = 32'd7374
; 
32'd169503: dataIn1 = 32'd7377
; 
32'd169504: dataIn1 = 32'd7378
; 
32'd169505: dataIn1 = 32'd5150
; 
32'd169506: dataIn1 = 32'd6195
; 
32'd169507: dataIn1 = 32'd7359
; 
32'd169508: dataIn1 = 32'd7372
; 
32'd169509: dataIn1 = 32'd7375
; 
32'd169510: dataIn1 = 32'd7379
; 
32'd169511: dataIn1 = 32'd7382
; 
32'd169512: dataIn1 = 32'd5151
; 
32'd169513: dataIn1 = 32'd6194
; 
32'd169514: dataIn1 = 32'd7361
; 
32'd169515: dataIn1 = 32'd7373
; 
32'd169516: dataIn1 = 32'd7376
; 
32'd169517: dataIn1 = 32'd7391
; 
32'd169518: dataIn1 = 32'd7408
; 
32'd169519: dataIn1 = 32'd2706
; 
32'd169520: dataIn1 = 32'd6195
; 
32'd169521: dataIn1 = 32'd7374
; 
32'd169522: dataIn1 = 32'd7377
; 
32'd169523: dataIn1 = 32'd7378
; 
32'd169524: dataIn1 = 32'd7381
; 
32'd169525: dataIn1 = 32'd7385
; 
32'd169526: dataIn1 = 32'd2706
; 
32'd169527: dataIn1 = 32'd6194
; 
32'd169528: dataIn1 = 32'd7374
; 
32'd169529: dataIn1 = 32'd7377
; 
32'd169530: dataIn1 = 32'd7378
; 
32'd169531: dataIn1 = 32'd7409
; 
32'd169532: dataIn1 = 32'd7411
; 
32'd169533: dataIn1 = 32'd6195
; 
32'd169534: dataIn1 = 32'd6197
; 
32'd169535: dataIn1 = 32'd7375
; 
32'd169536: dataIn1 = 32'd7379
; 
32'd169537: dataIn1 = 32'd7380
; 
32'd169538: dataIn1 = 32'd7381
; 
32'd169539: dataIn1 = 32'd7382
; 
32'd169540: dataIn1 = 32'd6196
; 
32'd169541: dataIn1 = 32'd6197
; 
32'd169542: dataIn1 = 32'd7379
; 
32'd169543: dataIn1 = 32'd7380
; 
32'd169544: dataIn1 = 32'd7381
; 
32'd169545: dataIn1 = 32'd7383
; 
32'd169546: dataIn1 = 32'd7384
; 
32'd169547: dataIn1 = 32'd6195
; 
32'd169548: dataIn1 = 32'd6196
; 
32'd169549: dataIn1 = 32'd7377
; 
32'd169550: dataIn1 = 32'd7379
; 
32'd169551: dataIn1 = 32'd7380
; 
32'd169552: dataIn1 = 32'd7381
; 
32'd169553: dataIn1 = 32'd7385
; 
32'd169554: dataIn1 = 32'd5150
; 
32'd169555: dataIn1 = 32'd6197
; 
32'd169556: dataIn1 = 32'd6747
; 
32'd169557: dataIn1 = 32'd7375
; 
32'd169558: dataIn1 = 32'd7379
; 
32'd169559: dataIn1 = 32'd7382
; 
32'd169560: dataIn1 = 32'd5153
; 
32'd169561: dataIn1 = 32'd6197
; 
32'd169562: dataIn1 = 32'd6746
; 
32'd169563: dataIn1 = 32'd7380
; 
32'd169564: dataIn1 = 32'd7383
; 
32'd169565: dataIn1 = 32'd7384
; 
32'd169566: dataIn1 = 32'd5153
; 
32'd169567: dataIn1 = 32'd6196
; 
32'd169568: dataIn1 = 32'd7380
; 
32'd169569: dataIn1 = 32'd7383
; 
32'd169570: dataIn1 = 32'd7384
; 
32'd169571: dataIn1 = 32'd7547
; 
32'd169572: dataIn1 = 32'd7557
; 
32'd169573: dataIn1 = 32'd2706
; 
32'd169574: dataIn1 = 32'd6196
; 
32'd169575: dataIn1 = 32'd7377
; 
32'd169576: dataIn1 = 32'd7381
; 
32'd169577: dataIn1 = 32'd7385
; 
32'd169578: dataIn1 = 32'd7540
; 
32'd169579: dataIn1 = 32'd7558
; 
32'd169580: dataIn1 = 32'd6199
; 
32'd169581: dataIn1 = 32'd6200
; 
32'd169582: dataIn1 = 32'd7386
; 
32'd169583: dataIn1 = 32'd7387
; 
32'd169584: dataIn1 = 32'd7388
; 
32'd169585: dataIn1 = 32'd7389
; 
32'd169586: dataIn1 = 32'd7390
; 
32'd169587: dataIn1 = 32'd6198
; 
32'd169588: dataIn1 = 32'd6200
; 
32'd169589: dataIn1 = 32'd7386
; 
32'd169590: dataIn1 = 32'd7387
; 
32'd169591: dataIn1 = 32'd7388
; 
32'd169592: dataIn1 = 32'd7391
; 
32'd169593: dataIn1 = 32'd7392
; 
32'd169594: dataIn1 = 32'd6198
; 
32'd169595: dataIn1 = 32'd6199
; 
32'd169596: dataIn1 = 32'd7386
; 
32'd169597: dataIn1 = 32'd7387
; 
32'd169598: dataIn1 = 32'd7388
; 
32'd169599: dataIn1 = 32'd7393
; 
32'd169600: dataIn1 = 32'd7394
; 
32'd169601: dataIn1 = 32'd5155
; 
32'd169602: dataIn1 = 32'd6200
; 
32'd169603: dataIn1 = 32'd7386
; 
32'd169604: dataIn1 = 32'd7389
; 
32'd169605: dataIn1 = 32'd7390
; 
32'd169606: dataIn1 = 32'd7407
; 
32'd169607: dataIn1 = 32'd7410
; 
32'd169608: dataIn1 = 32'd5155
; 
32'd169609: dataIn1 = 32'd6199
; 
32'd169610: dataIn1 = 32'd7386
; 
32'd169611: dataIn1 = 32'd7389
; 
32'd169612: dataIn1 = 32'd7390
; 
32'd169613: dataIn1 = 32'd7400
; 
32'd169614: dataIn1 = 32'd7403
; 
32'd169615: dataIn1 = 32'd5151
; 
32'd169616: dataIn1 = 32'd6200
; 
32'd169617: dataIn1 = 32'd7376
; 
32'd169618: dataIn1 = 32'd7387
; 
32'd169619: dataIn1 = 32'd7391
; 
32'd169620: dataIn1 = 32'd7392
; 
32'd169621: dataIn1 = 32'd7408
; 
32'd169622: dataIn1 = 32'd5151
; 
32'd169623: dataIn1 = 32'd6198
; 
32'd169624: dataIn1 = 32'd7370
; 
32'd169625: dataIn1 = 32'd7387
; 
32'd169626: dataIn1 = 32'd7391
; 
32'd169627: dataIn1 = 32'd7392
; 
32'd169628: dataIn1 = 32'd7396
; 
32'd169629: dataIn1 = 32'd5156
; 
32'd169630: dataIn1 = 32'd6199
; 
32'd169631: dataIn1 = 32'd7388
; 
32'd169632: dataIn1 = 32'd7393
; 
32'd169633: dataIn1 = 32'd7394
; 
32'd169634: dataIn1 = 32'd7402
; 
32'd169635: dataIn1 = 32'd7406
; 
32'd169636: dataIn1 = 32'd5156
; 
32'd169637: dataIn1 = 32'd6198
; 
32'd169638: dataIn1 = 32'd7388
; 
32'd169639: dataIn1 = 32'd7393
; 
32'd169640: dataIn1 = 32'd7394
; 
32'd169641: dataIn1 = 32'd7397
; 
32'd169642: dataIn1 = 32'd7399
; 
32'd169643: dataIn1 = 32'd6193
; 
32'd169644: dataIn1 = 32'd6201
; 
32'd169645: dataIn1 = 32'd7368
; 
32'd169646: dataIn1 = 32'd7395
; 
32'd169647: dataIn1 = 32'd7396
; 
32'd169648: dataIn1 = 32'd7397
; 
32'd169649: dataIn1 = 32'd7398
; 
32'd169650: dataIn1 = 32'd6193
; 
32'd169651: dataIn1 = 32'd6198
; 
32'd169652: dataIn1 = 32'd7370
; 
32'd169653: dataIn1 = 32'd7392
; 
32'd169654: dataIn1 = 32'd7395
; 
32'd169655: dataIn1 = 32'd7396
; 
32'd169656: dataIn1 = 32'd7397
; 
32'd169657: dataIn1 = 32'd6198
; 
32'd169658: dataIn1 = 32'd6201
; 
32'd169659: dataIn1 = 32'd7394
; 
32'd169660: dataIn1 = 32'd7395
; 
32'd169661: dataIn1 = 32'd7396
; 
32'd169662: dataIn1 = 32'd7397
; 
32'd169663: dataIn1 = 32'd7399
; 
32'd169664: dataIn1 = 32'd2704
; 
32'd169665: dataIn1 = 32'd6201
; 
32'd169666: dataIn1 = 32'd7368
; 
32'd169667: dataIn1 = 32'd7395
; 
32'd169668: dataIn1 = 32'd7398
; 
32'd169669: dataIn1 = 32'd7431
; 
32'd169670: dataIn1 = 32'd7482
; 
32'd169671: dataIn1 = 32'd5156
; 
32'd169672: dataIn1 = 32'd6201
; 
32'd169673: dataIn1 = 32'd7394
; 
32'd169674: dataIn1 = 32'd7397
; 
32'd169675: dataIn1 = 32'd7399
; 
32'd169676: dataIn1 = 32'd7481
; 
32'd169677: dataIn1 = 32'd7484
; 
32'd169678: dataIn1 = 32'd6199
; 
32'd169679: dataIn1 = 32'd6203
; 
32'd169680: dataIn1 = 32'd7390
; 
32'd169681: dataIn1 = 32'd7400
; 
32'd169682: dataIn1 = 32'd7401
; 
32'd169683: dataIn1 = 32'd7402
; 
32'd169684: dataIn1 = 32'd7403
; 
32'd169685: dataIn1 = 32'd6202
; 
32'd169686: dataIn1 = 32'd6203
; 
32'd169687: dataIn1 = 32'd7400
; 
32'd169688: dataIn1 = 32'd7401
; 
32'd169689: dataIn1 = 32'd7402
; 
32'd169690: dataIn1 = 32'd7404
; 
32'd169691: dataIn1 = 32'd7405
; 
32'd169692: dataIn1 = 32'd6199
; 
32'd169693: dataIn1 = 32'd6202
; 
32'd169694: dataIn1 = 32'd7393
; 
32'd169695: dataIn1 = 32'd7400
; 
32'd169696: dataIn1 = 32'd7401
; 
32'd169697: dataIn1 = 32'd7402
; 
32'd169698: dataIn1 = 32'd7406
; 
32'd169699: dataIn1 = 32'd5155
; 
32'd169700: dataIn1 = 32'd6203
; 
32'd169701: dataIn1 = 32'd7390
; 
32'd169702: dataIn1 = 32'd7400
; 
32'd169703: dataIn1 = 32'd7403
; 
32'd169704: dataIn1 = 32'd7563
; 
32'd169705: dataIn1 = 32'd7573
; 
32'd169706: dataIn1 = 32'd133
; 
32'd169707: dataIn1 = 32'd6203
; 
32'd169708: dataIn1 = 32'd7401
; 
32'd169709: dataIn1 = 32'd7404
; 
32'd169710: dataIn1 = 32'd7405
; 
32'd169711: dataIn1 = 32'd7574
; 
32'd169712: dataIn1 = 32'd7576
; 
32'd169713: dataIn1 = 32'd133
; 
32'd169714: dataIn1 = 32'd6202
; 
32'd169715: dataIn1 = 32'd7401
; 
32'd169716: dataIn1 = 32'd7404
; 
32'd169717: dataIn1 = 32'd7405
; 
32'd169718: dataIn1 = 32'd7486
; 
32'd169719: dataIn1 = 32'd7489
; 
32'd169720: dataIn1 = 32'd5156
; 
32'd169721: dataIn1 = 32'd6202
; 
32'd169722: dataIn1 = 32'd7393
; 
32'd169723: dataIn1 = 32'd7402
; 
32'd169724: dataIn1 = 32'd7406
; 
32'd169725: dataIn1 = 32'd7480
; 
32'd169726: dataIn1 = 32'd7487
; 
32'd169727: dataIn1 = 32'd6200
; 
32'd169728: dataIn1 = 32'd6204
; 
32'd169729: dataIn1 = 32'd7389
; 
32'd169730: dataIn1 = 32'd7407
; 
32'd169731: dataIn1 = 32'd7408
; 
32'd169732: dataIn1 = 32'd7409
; 
32'd169733: dataIn1 = 32'd7410
; 
32'd169734: dataIn1 = 32'd6194
; 
32'd169735: dataIn1 = 32'd6200
; 
32'd169736: dataIn1 = 32'd7376
; 
32'd169737: dataIn1 = 32'd7391
; 
32'd169738: dataIn1 = 32'd7407
; 
32'd169739: dataIn1 = 32'd7408
; 
32'd169740: dataIn1 = 32'd7409
; 
32'd169741: dataIn1 = 32'd6194
; 
32'd169742: dataIn1 = 32'd6204
; 
32'd169743: dataIn1 = 32'd7378
; 
32'd169744: dataIn1 = 32'd7407
; 
32'd169745: dataIn1 = 32'd7408
; 
32'd169746: dataIn1 = 32'd7409
; 
32'd169747: dataIn1 = 32'd7411
; 
32'd169748: dataIn1 = 32'd5155
; 
32'd169749: dataIn1 = 32'd6204
; 
32'd169750: dataIn1 = 32'd7389
; 
32'd169751: dataIn1 = 32'd7407
; 
32'd169752: dataIn1 = 32'd7410
; 
32'd169753: dataIn1 = 32'd7562
; 
32'd169754: dataIn1 = 32'd7578
; 
32'd169755: dataIn1 = 32'd2706
; 
32'd169756: dataIn1 = 32'd6204
; 
32'd169757: dataIn1 = 32'd7378
; 
32'd169758: dataIn1 = 32'd7409
; 
32'd169759: dataIn1 = 32'd7411
; 
32'd169760: dataIn1 = 32'd7541
; 
32'd169761: dataIn1 = 32'd7580
; 
32'd169762: dataIn1 = 32'd6192
; 
32'd169763: dataIn1 = 32'd6206
; 
32'd169764: dataIn1 = 32'd7369
; 
32'd169765: dataIn1 = 32'd7412
; 
32'd169766: dataIn1 = 32'd7413
; 
32'd169767: dataIn1 = 32'd7414
; 
32'd169768: dataIn1 = 32'd7415
; 
32'd169769: dataIn1 = 32'd6205
; 
32'd169770: dataIn1 = 32'd6206
; 
32'd169771: dataIn1 = 32'd7412
; 
32'd169772: dataIn1 = 32'd7413
; 
32'd169773: dataIn1 = 32'd7414
; 
32'd169774: dataIn1 = 32'd7416
; 
32'd169775: dataIn1 = 32'd7417
; 
32'd169776: dataIn1 = 32'd6192
; 
32'd169777: dataIn1 = 32'd6205
; 
32'd169778: dataIn1 = 32'd7371
; 
32'd169779: dataIn1 = 32'd7412
; 
32'd169780: dataIn1 = 32'd7413
; 
32'd169781: dataIn1 = 32'd7414
; 
32'd169782: dataIn1 = 32'd7418
; 
32'd169783: dataIn1 = 32'd2704
; 
32'd169784: dataIn1 = 32'd6206
; 
32'd169785: dataIn1 = 32'd7369
; 
32'd169786: dataIn1 = 32'd7412
; 
32'd169787: dataIn1 = 32'd7415
; 
32'd169788: dataIn1 = 32'd7432
; 
32'd169789: dataIn1 = 32'd7504
; 
32'd169790: dataIn1 = 32'd5158
; 
32'd169791: dataIn1 = 32'd6206
; 
32'd169792: dataIn1 = 32'd7413
; 
32'd169793: dataIn1 = 32'd7416
; 
32'd169794: dataIn1 = 32'd7417
; 
32'd169795: dataIn1 = 32'd7501
; 
32'd169796: dataIn1 = 32'd7505
; 
32'd169797: dataIn1 = 32'd5158
; 
32'd169798: dataIn1 = 32'd6205
; 
32'd169799: dataIn1 = 32'd6749
; 
32'd169800: dataIn1 = 32'd7413
; 
32'd169801: dataIn1 = 32'd7416
; 
32'd169802: dataIn1 = 32'd7417
; 
32'd169803: dataIn1 = 32'd5152
; 
32'd169804: dataIn1 = 32'd6205
; 
32'd169805: dataIn1 = 32'd6748
; 
32'd169806: dataIn1 = 32'd7371
; 
32'd169807: dataIn1 = 32'd7414
; 
32'd169808: dataIn1 = 32'd7418
; 
32'd169809: dataIn1 = 32'd6208
; 
32'd169810: dataIn1 = 32'd6209
; 
32'd169811: dataIn1 = 32'd7419
; 
32'd169812: dataIn1 = 32'd7420
; 
32'd169813: dataIn1 = 32'd7421
; 
32'd169814: dataIn1 = 32'd7422
; 
32'd169815: dataIn1 = 32'd7423
; 
32'd169816: dataIn1 = 32'd6207
; 
32'd169817: dataIn1 = 32'd6209
; 
32'd169818: dataIn1 = 32'd7419
; 
32'd169819: dataIn1 = 32'd7420
; 
32'd169820: dataIn1 = 32'd7421
; 
32'd169821: dataIn1 = 32'd7424
; 
32'd169822: dataIn1 = 32'd7425
; 
32'd169823: dataIn1 = 32'd6207
; 
32'd169824: dataIn1 = 32'd6208
; 
32'd169825: dataIn1 = 32'd7419
; 
32'd169826: dataIn1 = 32'd7420
; 
32'd169827: dataIn1 = 32'd7421
; 
32'd169828: dataIn1 = 32'd7426
; 
32'd169829: dataIn1 = 32'd7427
; 
32'd169830: dataIn1 = 32'd5159
; 
32'd169831: dataIn1 = 32'd6209
; 
32'd169832: dataIn1 = 32'd7419
; 
32'd169833: dataIn1 = 32'd7422
; 
32'd169834: dataIn1 = 32'd7423
; 
32'd169835: dataIn1 = 32'd7442
; 
32'd169836: dataIn1 = 32'd7445
; 
32'd169837: dataIn1 = 32'd5159
; 
32'd169838: dataIn1 = 32'd6208
; 
32'd169839: dataIn1 = 32'd7419
; 
32'd169840: dataIn1 = 32'd7422
; 
32'd169841: dataIn1 = 32'd7423
; 
32'd169842: dataIn1 = 32'd7435
; 
32'd169843: dataIn1 = 32'd7438
; 
32'd169844: dataIn1 = 32'd5160
; 
32'd169845: dataIn1 = 32'd6209
; 
32'd169846: dataIn1 = 32'd7420
; 
32'd169847: dataIn1 = 32'd7424
; 
32'd169848: dataIn1 = 32'd7425
; 
32'd169849: dataIn1 = 32'd7443
; 
32'd169850: dataIn1 = 32'd7446
; 
32'd169851: dataIn1 = 32'd5160
; 
32'd169852: dataIn1 = 32'd6207
; 
32'd169853: dataIn1 = 32'd7420
; 
32'd169854: dataIn1 = 32'd7424
; 
32'd169855: dataIn1 = 32'd7425
; 
32'd169856: dataIn1 = 32'd7429
; 
32'd169857: dataIn1 = 32'd7433
; 
32'd169858: dataIn1 = 32'd5161
; 
32'd169859: dataIn1 = 32'd6208
; 
32'd169860: dataIn1 = 32'd7421
; 
32'd169861: dataIn1 = 32'd7426
; 
32'd169862: dataIn1 = 32'd7427
; 
32'd169863: dataIn1 = 32'd7437
; 
32'd169864: dataIn1 = 32'd7441
; 
32'd169865: dataIn1 = 32'd5161
; 
32'd169866: dataIn1 = 32'd6207
; 
32'd169867: dataIn1 = 32'd7421
; 
32'd169868: dataIn1 = 32'd7426
; 
32'd169869: dataIn1 = 32'd7427
; 
32'd169870: dataIn1 = 32'd7430
; 
32'd169871: dataIn1 = 32'd7434
; 
32'd169872: dataIn1 = 32'd6210
; 
32'd169873: dataIn1 = 32'd6211
; 
32'd169874: dataIn1 = 32'd7428
; 
32'd169875: dataIn1 = 32'd7429
; 
32'd169876: dataIn1 = 32'd7430
; 
32'd169877: dataIn1 = 32'd7431
; 
32'd169878: dataIn1 = 32'd7432
; 
32'd169879: dataIn1 = 32'd6207
; 
32'd169880: dataIn1 = 32'd6211
; 
32'd169881: dataIn1 = 32'd7425
; 
32'd169882: dataIn1 = 32'd7428
; 
32'd169883: dataIn1 = 32'd7429
; 
32'd169884: dataIn1 = 32'd7430
; 
32'd169885: dataIn1 = 32'd7433
; 
32'd169886: dataIn1 = 32'd6207
; 
32'd169887: dataIn1 = 32'd6210
; 
32'd169888: dataIn1 = 32'd7427
; 
32'd169889: dataIn1 = 32'd7428
; 
32'd169890: dataIn1 = 32'd7429
; 
32'd169891: dataIn1 = 32'd7430
; 
32'd169892: dataIn1 = 32'd7434
; 
32'd169893: dataIn1 = 32'd2704
; 
32'd169894: dataIn1 = 32'd6211
; 
32'd169895: dataIn1 = 32'd7398
; 
32'd169896: dataIn1 = 32'd7428
; 
32'd169897: dataIn1 = 32'd7431
; 
32'd169898: dataIn1 = 32'd7432
; 
32'd169899: dataIn1 = 32'd7482
; 
32'd169900: dataIn1 = 32'd2704
; 
32'd169901: dataIn1 = 32'd6210
; 
32'd169902: dataIn1 = 32'd7415
; 
32'd169903: dataIn1 = 32'd7428
; 
32'd169904: dataIn1 = 32'd7431
; 
32'd169905: dataIn1 = 32'd7432
; 
32'd169906: dataIn1 = 32'd7504
; 
32'd169907: dataIn1 = 32'd5160
; 
32'd169908: dataIn1 = 32'd6211
; 
32'd169909: dataIn1 = 32'd7425
; 
32'd169910: dataIn1 = 32'd7429
; 
32'd169911: dataIn1 = 32'd7433
; 
32'd169912: dataIn1 = 32'd7479
; 
32'd169913: dataIn1 = 32'd7483
; 
32'd169914: dataIn1 = 32'd5161
; 
32'd169915: dataIn1 = 32'd6210
; 
32'd169916: dataIn1 = 32'd7427
; 
32'd169917: dataIn1 = 32'd7430
; 
32'd169918: dataIn1 = 32'd7434
; 
32'd169919: dataIn1 = 32'd7503
; 
32'd169920: dataIn1 = 32'd7506
; 
32'd169921: dataIn1 = 32'd6208
; 
32'd169922: dataIn1 = 32'd6213
; 
32'd169923: dataIn1 = 32'd7423
; 
32'd169924: dataIn1 = 32'd7435
; 
32'd169925: dataIn1 = 32'd7436
; 
32'd169926: dataIn1 = 32'd7437
; 
32'd169927: dataIn1 = 32'd7438
; 
32'd169928: dataIn1 = 32'd6212
; 
32'd169929: dataIn1 = 32'd6213
; 
32'd169930: dataIn1 = 32'd7435
; 
32'd169931: dataIn1 = 32'd7436
; 
32'd169932: dataIn1 = 32'd7437
; 
32'd169933: dataIn1 = 32'd7439
; 
32'd169934: dataIn1 = 32'd7440
; 
32'd169935: dataIn1 = 32'd6208
; 
32'd169936: dataIn1 = 32'd6212
; 
32'd169937: dataIn1 = 32'd7426
; 
32'd169938: dataIn1 = 32'd7435
; 
32'd169939: dataIn1 = 32'd7436
; 
32'd169940: dataIn1 = 32'd7437
; 
32'd169941: dataIn1 = 32'd7441
; 
32'd169942: dataIn1 = 32'd5159
; 
32'd169943: dataIn1 = 32'd6213
; 
32'd169944: dataIn1 = 32'd7423
; 
32'd169945: dataIn1 = 32'd7435
; 
32'd169946: dataIn1 = 32'd7438
; 
32'd169947: dataIn1 = 32'd7453
; 
32'd169948: dataIn1 = 32'd7463
; 
32'd169949: dataIn1 = 32'd2707
; 
32'd169950: dataIn1 = 32'd6213
; 
32'd169951: dataIn1 = 32'd7436
; 
32'd169952: dataIn1 = 32'd7439
; 
32'd169953: dataIn1 = 32'd7440
; 
32'd169954: dataIn1 = 32'd7464
; 
32'd169955: dataIn1 = 32'd7466
; 
32'd169956: dataIn1 = 32'd2707
; 
32'd169957: dataIn1 = 32'd6212
; 
32'd169958: dataIn1 = 32'd7436
; 
32'd169959: dataIn1 = 32'd7439
; 
32'd169960: dataIn1 = 32'd7440
; 
32'd169961: dataIn1 = 32'd7508
; 
32'd169962: dataIn1 = 32'd7511
; 
32'd169963: dataIn1 = 32'd5161
; 
32'd169964: dataIn1 = 32'd6212
; 
32'd169965: dataIn1 = 32'd7426
; 
32'd169966: dataIn1 = 32'd7437
; 
32'd169967: dataIn1 = 32'd7441
; 
32'd169968: dataIn1 = 32'd7502
; 
32'd169969: dataIn1 = 32'd7509
; 
32'd169970: dataIn1 = 32'd6209
; 
32'd169971: dataIn1 = 32'd6215
; 
32'd169972: dataIn1 = 32'd7422
; 
32'd169973: dataIn1 = 32'd7442
; 
32'd169974: dataIn1 = 32'd7443
; 
32'd169975: dataIn1 = 32'd7444
; 
32'd169976: dataIn1 = 32'd7445
; 
32'd169977: dataIn1 = 32'd6209
; 
32'd169978: dataIn1 = 32'd6214
; 
32'd169979: dataIn1 = 32'd7424
; 
32'd169980: dataIn1 = 32'd7442
; 
32'd169981: dataIn1 = 32'd7443
; 
32'd169982: dataIn1 = 32'd7444
; 
32'd169983: dataIn1 = 32'd7446
; 
32'd169984: dataIn1 = 32'd6214
; 
32'd169985: dataIn1 = 32'd6215
; 
32'd169986: dataIn1 = 32'd7442
; 
32'd169987: dataIn1 = 32'd7443
; 
32'd169988: dataIn1 = 32'd7444
; 
32'd169989: dataIn1 = 32'd7447
; 
32'd169990: dataIn1 = 32'd7448
; 
32'd169991: dataIn1 = 32'd5159
; 
32'd169992: dataIn1 = 32'd6215
; 
32'd169993: dataIn1 = 32'd7422
; 
32'd169994: dataIn1 = 32'd7442
; 
32'd169995: dataIn1 = 32'd7445
; 
32'd169996: dataIn1 = 32'd7452
; 
32'd169997: dataIn1 = 32'd7468
; 
32'd169998: dataIn1 = 32'd5160
; 
32'd169999: dataIn1 = 32'd6214
; 
32'd170000: dataIn1 = 32'd7424
; 
32'd170001: dataIn1 = 32'd7443
; 
32'd170002: dataIn1 = 32'd7446
; 
32'd170003: dataIn1 = 32'd7478
; 
32'd170004: dataIn1 = 32'd7491
; 
32'd170005: dataIn1 = 32'd1107
; 
32'd170006: dataIn1 = 32'd6215
; 
32'd170007: dataIn1 = 32'd7444
; 
32'd170008: dataIn1 = 32'd7447
; 
32'd170009: dataIn1 = 32'd7448
; 
32'd170010: dataIn1 = 32'd7470
; 
32'd170011: dataIn1 = 32'd7472
; 
32'd170012: dataIn1 = 32'd1107
; 
32'd170013: dataIn1 = 32'd6214
; 
32'd170014: dataIn1 = 32'd7444
; 
32'd170015: dataIn1 = 32'd7447
; 
32'd170016: dataIn1 = 32'd7448
; 
32'd170017: dataIn1 = 32'd7492
; 
32'd170018: dataIn1 = 32'd7494
; 
32'd170019: dataIn1 = 32'd6217
; 
32'd170020: dataIn1 = 32'd6218
; 
32'd170021: dataIn1 = 32'd7449
; 
32'd170022: dataIn1 = 32'd7450
; 
32'd170023: dataIn1 = 32'd7451
; 
32'd170024: dataIn1 = 32'd7452
; 
32'd170025: dataIn1 = 32'd7453
; 
32'd170026: dataIn1 = 32'd6216
; 
32'd170027: dataIn1 = 32'd6218
; 
32'd170028: dataIn1 = 32'd7449
; 
32'd170029: dataIn1 = 32'd7450
; 
32'd170030: dataIn1 = 32'd7451
; 
32'd170031: dataIn1 = 32'd7454
; 
32'd170032: dataIn1 = 32'd7455
; 
32'd170033: dataIn1 = 32'd6216
; 
32'd170034: dataIn1 = 32'd6217
; 
32'd170035: dataIn1 = 32'd7449
; 
32'd170036: dataIn1 = 32'd7450
; 
32'd170037: dataIn1 = 32'd7451
; 
32'd170038: dataIn1 = 32'd7456
; 
32'd170039: dataIn1 = 32'd7457
; 
32'd170040: dataIn1 = 32'd5159
; 
32'd170041: dataIn1 = 32'd6218
; 
32'd170042: dataIn1 = 32'd7445
; 
32'd170043: dataIn1 = 32'd7449
; 
32'd170044: dataIn1 = 32'd7452
; 
32'd170045: dataIn1 = 32'd7453
; 
32'd170046: dataIn1 = 32'd7468
; 
32'd170047: dataIn1 = 32'd5159
; 
32'd170048: dataIn1 = 32'd6217
; 
32'd170049: dataIn1 = 32'd7438
; 
32'd170050: dataIn1 = 32'd7449
; 
32'd170051: dataIn1 = 32'd7452
; 
32'd170052: dataIn1 = 32'd7453
; 
32'd170053: dataIn1 = 32'd7463
; 
32'd170054: dataIn1 = 32'd2636
; 
32'd170055: dataIn1 = 32'd6218
; 
32'd170056: dataIn1 = 32'd7450
; 
32'd170057: dataIn1 = 32'd7454
; 
32'd170058: dataIn1 = 32'd7455
; 
32'd170059: dataIn1 = 32'd7469
; 
32'd170060: dataIn1 = 32'd7471
; 
32'd170061: dataIn1 = 32'd2636
; 
32'd170062: dataIn1 = 32'd6216
; 
32'd170063: dataIn1 = 32'd7450
; 
32'd170064: dataIn1 = 32'd7454
; 
32'd170065: dataIn1 = 32'd7455
; 
32'd170066: dataIn1 = 32'd7459
; 
32'd170067: dataIn1 = 32'd7461
; 
32'd170068: dataIn1 = 32'd5162
; 
32'd170069: dataIn1 = 32'd6217
; 
32'd170070: dataIn1 = 32'd7451
; 
32'd170071: dataIn1 = 32'd7456
; 
32'd170072: dataIn1 = 32'd7457
; 
32'd170073: dataIn1 = 32'd7465
; 
32'd170074: dataIn1 = 32'd7467
; 
32'd170075: dataIn1 = 32'd5162
; 
32'd170076: dataIn1 = 32'd6216
; 
32'd170077: dataIn1 = 32'd7451
; 
32'd170078: dataIn1 = 32'd7456
; 
32'd170079: dataIn1 = 32'd7457
; 
32'd170080: dataIn1 = 32'd7460
; 
32'd170081: dataIn1 = 32'd7462
; 
32'd170082: dataIn1 = 32'd4901
; 
32'd170083: dataIn1 = 32'd6065
; 
32'd170084: dataIn1 = 32'd6219
; 
32'd170085: dataIn1 = 32'd7458
; 
32'd170086: dataIn1 = 32'd7459
; 
32'd170087: dataIn1 = 32'd7460
; 
32'd170088: dataIn1 = 32'd8962
; 
32'd170089: dataIn1 = 32'd4901
; 
32'd170090: dataIn1 = 32'd6216
; 
32'd170091: dataIn1 = 32'd7455
; 
32'd170092: dataIn1 = 32'd7458
; 
32'd170093: dataIn1 = 32'd7459
; 
32'd170094: dataIn1 = 32'd7460
; 
32'd170095: dataIn1 = 32'd7461
; 
32'd170096: dataIn1 = 32'd6216
; 
32'd170097: dataIn1 = 32'd6219
; 
32'd170098: dataIn1 = 32'd7457
; 
32'd170099: dataIn1 = 32'd7458
; 
32'd170100: dataIn1 = 32'd7459
; 
32'd170101: dataIn1 = 32'd7460
; 
32'd170102: dataIn1 = 32'd7462
; 
32'd170103: dataIn1 = 32'd2636
; 
32'd170104: dataIn1 = 32'd4899
; 
32'd170105: dataIn1 = 32'd4901
; 
32'd170106: dataIn1 = 32'd7455
; 
32'd170107: dataIn1 = 32'd7459
; 
32'd170108: dataIn1 = 32'd7461
; 
32'd170109: dataIn1 = 32'd5162
; 
32'd170110: dataIn1 = 32'd6219
; 
32'd170111: dataIn1 = 32'd7457
; 
32'd170112: dataIn1 = 32'd7460
; 
32'd170113: dataIn1 = 32'd7462
; 
32'd170114: dataIn1 = 32'd8956
; 
32'd170115: dataIn1 = 32'd8960
; 
32'd170116: dataIn1 = 32'd6213
; 
32'd170117: dataIn1 = 32'd6217
; 
32'd170118: dataIn1 = 32'd7438
; 
32'd170119: dataIn1 = 32'd7453
; 
32'd170120: dataIn1 = 32'd7463
; 
32'd170121: dataIn1 = 32'd7464
; 
32'd170122: dataIn1 = 32'd7465
; 
32'd170123: dataIn1 = 32'd6213
; 
32'd170124: dataIn1 = 32'd6220
; 
32'd170125: dataIn1 = 32'd7439
; 
32'd170126: dataIn1 = 32'd7463
; 
32'd170127: dataIn1 = 32'd7464
; 
32'd170128: dataIn1 = 32'd7465
; 
32'd170129: dataIn1 = 32'd7466
; 
32'd170130: dataIn1 = 32'd6217
; 
32'd170131: dataIn1 = 32'd6220
; 
32'd170132: dataIn1 = 32'd7456
; 
32'd170133: dataIn1 = 32'd7463
; 
32'd170134: dataIn1 = 32'd7464
; 
32'd170135: dataIn1 = 32'd7465
; 
32'd170136: dataIn1 = 32'd7467
; 
32'd170137: dataIn1 = 32'd2707
; 
32'd170138: dataIn1 = 32'd6220
; 
32'd170139: dataIn1 = 32'd7439
; 
32'd170140: dataIn1 = 32'd7464
; 
32'd170141: dataIn1 = 32'd7466
; 
32'd170142: dataIn1 = 32'd8948
; 
32'd170143: dataIn1 = 32'd8969
; 
32'd170144: dataIn1 = 32'd5162
; 
32'd170145: dataIn1 = 32'd6220
; 
32'd170146: dataIn1 = 32'd7456
; 
32'd170147: dataIn1 = 32'd7465
; 
32'd170148: dataIn1 = 32'd7467
; 
32'd170149: dataIn1 = 32'd8955
; 
32'd170150: dataIn1 = 32'd8968
; 
32'd170151: dataIn1 = 32'd6215
; 
32'd170152: dataIn1 = 32'd6218
; 
32'd170153: dataIn1 = 32'd7445
; 
32'd170154: dataIn1 = 32'd7452
; 
32'd170155: dataIn1 = 32'd7468
; 
32'd170156: dataIn1 = 32'd7469
; 
32'd170157: dataIn1 = 32'd7470
; 
32'd170158: dataIn1 = 32'd4902
; 
32'd170159: dataIn1 = 32'd6218
; 
32'd170160: dataIn1 = 32'd7454
; 
32'd170161: dataIn1 = 32'd7468
; 
32'd170162: dataIn1 = 32'd7469
; 
32'd170163: dataIn1 = 32'd7470
; 
32'd170164: dataIn1 = 32'd7471
; 
32'd170165: dataIn1 = 32'd4902
; 
32'd170166: dataIn1 = 32'd6215
; 
32'd170167: dataIn1 = 32'd7447
; 
32'd170168: dataIn1 = 32'd7468
; 
32'd170169: dataIn1 = 32'd7469
; 
32'd170170: dataIn1 = 32'd7470
; 
32'd170171: dataIn1 = 32'd7472
; 
32'd170172: dataIn1 = 32'd2636
; 
32'd170173: dataIn1 = 32'd4900
; 
32'd170174: dataIn1 = 32'd4902
; 
32'd170175: dataIn1 = 32'd7454
; 
32'd170176: dataIn1 = 32'd7469
; 
32'd170177: dataIn1 = 32'd7471
; 
32'd170178: dataIn1 = 32'd1107
; 
32'd170179: dataIn1 = 32'd4902
; 
32'd170180: dataIn1 = 32'd7447
; 
32'd170181: dataIn1 = 32'd7470
; 
32'd170182: dataIn1 = 32'd7472
; 
32'd170183: dataIn1 = 32'd9612
; 
32'd170184: dataIn1 = 32'd9763
; 
32'd170185: dataIn1 = 32'd6222
; 
32'd170186: dataIn1 = 32'd6223
; 
32'd170187: dataIn1 = 32'd7473
; 
32'd170188: dataIn1 = 32'd7474
; 
32'd170189: dataIn1 = 32'd7475
; 
32'd170190: dataIn1 = 32'd7476
; 
32'd170191: dataIn1 = 32'd7477
; 
32'd170192: dataIn1 = 32'd6221
; 
32'd170193: dataIn1 = 32'd6223
; 
32'd170194: dataIn1 = 32'd7473
; 
32'd170195: dataIn1 = 32'd7474
; 
32'd170196: dataIn1 = 32'd7475
; 
32'd170197: dataIn1 = 32'd7478
; 
32'd170198: dataIn1 = 32'd7479
; 
32'd170199: dataIn1 = 32'd6221
; 
32'd170200: dataIn1 = 32'd6222
; 
32'd170201: dataIn1 = 32'd7473
; 
32'd170202: dataIn1 = 32'd7474
; 
32'd170203: dataIn1 = 32'd7475
; 
32'd170204: dataIn1 = 32'd7480
; 
32'd170205: dataIn1 = 32'd7481
; 
32'd170206: dataIn1 = 32'd2635
; 
32'd170207: dataIn1 = 32'd6223
; 
32'd170208: dataIn1 = 32'd7473
; 
32'd170209: dataIn1 = 32'd7476
; 
32'd170210: dataIn1 = 32'd7477
; 
32'd170211: dataIn1 = 32'd7490
; 
32'd170212: dataIn1 = 32'd7493
; 
32'd170213: dataIn1 = 32'd2635
; 
32'd170214: dataIn1 = 32'd6222
; 
32'd170215: dataIn1 = 32'd7473
; 
32'd170216: dataIn1 = 32'd7476
; 
32'd170217: dataIn1 = 32'd7477
; 
32'd170218: dataIn1 = 32'd7485
; 
32'd170219: dataIn1 = 32'd7488
; 
32'd170220: dataIn1 = 32'd5160
; 
32'd170221: dataIn1 = 32'd6223
; 
32'd170222: dataIn1 = 32'd7446
; 
32'd170223: dataIn1 = 32'd7474
; 
32'd170224: dataIn1 = 32'd7478
; 
32'd170225: dataIn1 = 32'd7479
; 
32'd170226: dataIn1 = 32'd7491
; 
32'd170227: dataIn1 = 32'd5160
; 
32'd170228: dataIn1 = 32'd6221
; 
32'd170229: dataIn1 = 32'd7433
; 
32'd170230: dataIn1 = 32'd7474
; 
32'd170231: dataIn1 = 32'd7478
; 
32'd170232: dataIn1 = 32'd7479
; 
32'd170233: dataIn1 = 32'd7483
; 
32'd170234: dataIn1 = 32'd5156
; 
32'd170235: dataIn1 = 32'd6222
; 
32'd170236: dataIn1 = 32'd7406
; 
32'd170237: dataIn1 = 32'd7475
; 
32'd170238: dataIn1 = 32'd7480
; 
32'd170239: dataIn1 = 32'd7481
; 
32'd170240: dataIn1 = 32'd7487
; 
32'd170241: dataIn1 = 32'd5156
; 
32'd170242: dataIn1 = 32'd6221
; 
32'd170243: dataIn1 = 32'd7399
; 
32'd170244: dataIn1 = 32'd7475
; 
32'd170245: dataIn1 = 32'd7480
; 
32'd170246: dataIn1 = 32'd7481
; 
32'd170247: dataIn1 = 32'd7484
; 
32'd170248: dataIn1 = 32'd6201
; 
32'd170249: dataIn1 = 32'd6211
; 
32'd170250: dataIn1 = 32'd7398
; 
32'd170251: dataIn1 = 32'd7431
; 
32'd170252: dataIn1 = 32'd7482
; 
32'd170253: dataIn1 = 32'd7483
; 
32'd170254: dataIn1 = 32'd7484
; 
32'd170255: dataIn1 = 32'd6211
; 
32'd170256: dataIn1 = 32'd6221
; 
32'd170257: dataIn1 = 32'd7433
; 
32'd170258: dataIn1 = 32'd7479
; 
32'd170259: dataIn1 = 32'd7482
; 
32'd170260: dataIn1 = 32'd7483
; 
32'd170261: dataIn1 = 32'd7484
; 
32'd170262: dataIn1 = 32'd6201
; 
32'd170263: dataIn1 = 32'd6221
; 
32'd170264: dataIn1 = 32'd7399
; 
32'd170265: dataIn1 = 32'd7481
; 
32'd170266: dataIn1 = 32'd7482
; 
32'd170267: dataIn1 = 32'd7483
; 
32'd170268: dataIn1 = 32'd7484
; 
32'd170269: dataIn1 = 32'd4896
; 
32'd170270: dataIn1 = 32'd6222
; 
32'd170271: dataIn1 = 32'd7477
; 
32'd170272: dataIn1 = 32'd7485
; 
32'd170273: dataIn1 = 32'd7486
; 
32'd170274: dataIn1 = 32'd7487
; 
32'd170275: dataIn1 = 32'd7488
; 
32'd170276: dataIn1 = 32'd4896
; 
32'd170277: dataIn1 = 32'd6202
; 
32'd170278: dataIn1 = 32'd7405
; 
32'd170279: dataIn1 = 32'd7485
; 
32'd170280: dataIn1 = 32'd7486
; 
32'd170281: dataIn1 = 32'd7487
; 
32'd170282: dataIn1 = 32'd7489
; 
32'd170283: dataIn1 = 32'd6202
; 
32'd170284: dataIn1 = 32'd6222
; 
32'd170285: dataIn1 = 32'd7406
; 
32'd170286: dataIn1 = 32'd7480
; 
32'd170287: dataIn1 = 32'd7485
; 
32'd170288: dataIn1 = 32'd7486
; 
32'd170289: dataIn1 = 32'd7487
; 
32'd170290: dataIn1 = 32'd2635
; 
32'd170291: dataIn1 = 32'd4896
; 
32'd170292: dataIn1 = 32'd7477
; 
32'd170293: dataIn1 = 32'd7485
; 
32'd170294: dataIn1 = 32'd7488
; 
32'd170295: dataIn1 = 32'd9616
; 
32'd170296: dataIn1 = 32'd9618
; 
32'd170297: dataIn1 = 32'd133
; 
32'd170298: dataIn1 = 32'd4896
; 
32'd170299: dataIn1 = 32'd7405
; 
32'd170300: dataIn1 = 32'd7486
; 
32'd170301: dataIn1 = 32'd7489
; 
32'd170302: dataIn1 = 32'd9604
; 
32'd170303: dataIn1 = 32'd9617
; 
32'd170304: dataIn1 = 32'd4897
; 
32'd170305: dataIn1 = 32'd6223
; 
32'd170306: dataIn1 = 32'd7476
; 
32'd170307: dataIn1 = 32'd7490
; 
32'd170308: dataIn1 = 32'd7491
; 
32'd170309: dataIn1 = 32'd7492
; 
32'd170310: dataIn1 = 32'd7493
; 
32'd170311: dataIn1 = 32'd6214
; 
32'd170312: dataIn1 = 32'd6223
; 
32'd170313: dataIn1 = 32'd7446
; 
32'd170314: dataIn1 = 32'd7478
; 
32'd170315: dataIn1 = 32'd7490
; 
32'd170316: dataIn1 = 32'd7491
; 
32'd170317: dataIn1 = 32'd7492
; 
32'd170318: dataIn1 = 32'd4897
; 
32'd170319: dataIn1 = 32'd6214
; 
32'd170320: dataIn1 = 32'd7448
; 
32'd170321: dataIn1 = 32'd7490
; 
32'd170322: dataIn1 = 32'd7491
; 
32'd170323: dataIn1 = 32'd7492
; 
32'd170324: dataIn1 = 32'd7494
; 
32'd170325: dataIn1 = 32'd2635
; 
32'd170326: dataIn1 = 32'd4897
; 
32'd170327: dataIn1 = 32'd7476
; 
32'd170328: dataIn1 = 32'd7490
; 
32'd170329: dataIn1 = 32'd7493
; 
32'd170330: dataIn1 = 32'd9614
; 
32'd170331: dataIn1 = 32'd9621
; 
32'd170332: dataIn1 = 32'd1107
; 
32'd170333: dataIn1 = 32'd4897
; 
32'd170334: dataIn1 = 32'd7448
; 
32'd170335: dataIn1 = 32'd7492
; 
32'd170336: dataIn1 = 32'd7494
; 
32'd170337: dataIn1 = 32'd9611
; 
32'd170338: dataIn1 = 32'd9622
; 
32'd170339: dataIn1 = 32'd6225
; 
32'd170340: dataIn1 = 32'd6226
; 
32'd170341: dataIn1 = 32'd7495
; 
32'd170342: dataIn1 = 32'd7496
; 
32'd170343: dataIn1 = 32'd7497
; 
32'd170344: dataIn1 = 32'd7498
; 
32'd170345: dataIn1 = 32'd7499
; 
32'd170346: dataIn1 = 32'd6224
; 
32'd170347: dataIn1 = 32'd6226
; 
32'd170348: dataIn1 = 32'd7495
; 
32'd170349: dataIn1 = 32'd7496
; 
32'd170350: dataIn1 = 32'd7497
; 
32'd170351: dataIn1 = 32'd7500
; 
32'd170352: dataIn1 = 32'd7501
; 
32'd170353: dataIn1 = 32'd6224
; 
32'd170354: dataIn1 = 32'd6225
; 
32'd170355: dataIn1 = 32'd7495
; 
32'd170356: dataIn1 = 32'd7496
; 
32'd170357: dataIn1 = 32'd7497
; 
32'd170358: dataIn1 = 32'd7502
; 
32'd170359: dataIn1 = 32'd7503
; 
32'd170360: dataIn1 = 32'd5163
; 
32'd170361: dataIn1 = 32'd6226
; 
32'd170362: dataIn1 = 32'd6751
; 
32'd170363: dataIn1 = 32'd7495
; 
32'd170364: dataIn1 = 32'd7498
; 
32'd170365: dataIn1 = 32'd7499
; 
32'd170366: dataIn1 = 32'd5163
; 
32'd170367: dataIn1 = 32'd6225
; 
32'd170368: dataIn1 = 32'd7495
; 
32'd170369: dataIn1 = 32'd7498
; 
32'd170370: dataIn1 = 32'd7499
; 
32'd170371: dataIn1 = 32'd7507
; 
32'd170372: dataIn1 = 32'd7510
; 
32'd170373: dataIn1 = 32'd5158
; 
32'd170374: dataIn1 = 32'd6226
; 
32'd170375: dataIn1 = 32'd6750
; 
32'd170376: dataIn1 = 32'd7496
; 
32'd170377: dataIn1 = 32'd7500
; 
32'd170378: dataIn1 = 32'd7501
; 
32'd170379: dataIn1 = 32'd5158
; 
32'd170380: dataIn1 = 32'd6224
; 
32'd170381: dataIn1 = 32'd7416
; 
32'd170382: dataIn1 = 32'd7496
; 
32'd170383: dataIn1 = 32'd7500
; 
32'd170384: dataIn1 = 32'd7501
; 
32'd170385: dataIn1 = 32'd7505
; 
32'd170386: dataIn1 = 32'd5161
; 
32'd170387: dataIn1 = 32'd6225
; 
32'd170388: dataIn1 = 32'd7441
; 
32'd170389: dataIn1 = 32'd7497
; 
32'd170390: dataIn1 = 32'd7502
; 
32'd170391: dataIn1 = 32'd7503
; 
32'd170392: dataIn1 = 32'd7509
; 
32'd170393: dataIn1 = 32'd5161
; 
32'd170394: dataIn1 = 32'd6224
; 
32'd170395: dataIn1 = 32'd7434
; 
32'd170396: dataIn1 = 32'd7497
; 
32'd170397: dataIn1 = 32'd7502
; 
32'd170398: dataIn1 = 32'd7503
; 
32'd170399: dataIn1 = 32'd7506
; 
32'd170400: dataIn1 = 32'd6206
; 
32'd170401: dataIn1 = 32'd6210
; 
32'd170402: dataIn1 = 32'd7415
; 
32'd170403: dataIn1 = 32'd7432
; 
32'd170404: dataIn1 = 32'd7504
; 
32'd170405: dataIn1 = 32'd7505
; 
32'd170406: dataIn1 = 32'd7506
; 
32'd170407: dataIn1 = 32'd6206
; 
32'd170408: dataIn1 = 32'd6224
; 
32'd170409: dataIn1 = 32'd7416
; 
32'd170410: dataIn1 = 32'd7501
; 
32'd170411: dataIn1 = 32'd7504
; 
32'd170412: dataIn1 = 32'd7505
; 
32'd170413: dataIn1 = 32'd7506
; 
32'd170414: dataIn1 = 32'd6210
; 
32'd170415: dataIn1 = 32'd6224
; 
32'd170416: dataIn1 = 32'd7434
; 
32'd170417: dataIn1 = 32'd7503
; 
32'd170418: dataIn1 = 32'd7504
; 
32'd170419: dataIn1 = 32'd7505
; 
32'd170420: dataIn1 = 32'd7506
; 
32'd170421: dataIn1 = 32'd6225
; 
32'd170422: dataIn1 = 32'd6227
; 
32'd170423: dataIn1 = 32'd7499
; 
32'd170424: dataIn1 = 32'd7507
; 
32'd170425: dataIn1 = 32'd7508
; 
32'd170426: dataIn1 = 32'd7509
; 
32'd170427: dataIn1 = 32'd7510
; 
32'd170428: dataIn1 = 32'd6212
; 
32'd170429: dataIn1 = 32'd6227
; 
32'd170430: dataIn1 = 32'd7440
; 
32'd170431: dataIn1 = 32'd7507
; 
32'd170432: dataIn1 = 32'd7508
; 
32'd170433: dataIn1 = 32'd7509
; 
32'd170434: dataIn1 = 32'd7511
; 
32'd170435: dataIn1 = 32'd6212
; 
32'd170436: dataIn1 = 32'd6225
; 
32'd170437: dataIn1 = 32'd7441
; 
32'd170438: dataIn1 = 32'd7502
; 
32'd170439: dataIn1 = 32'd7507
; 
32'd170440: dataIn1 = 32'd7508
; 
32'd170441: dataIn1 = 32'd7509
; 
32'd170442: dataIn1 = 32'd5163
; 
32'd170443: dataIn1 = 32'd6227
; 
32'd170444: dataIn1 = 32'd7499
; 
32'd170445: dataIn1 = 32'd7507
; 
32'd170446: dataIn1 = 32'd7510
; 
32'd170447: dataIn1 = 32'd8970
; 
32'd170448: dataIn1 = 32'd8973
; 
32'd170449: dataIn1 = 32'd2707
; 
32'd170450: dataIn1 = 32'd6227
; 
32'd170451: dataIn1 = 32'd7440
; 
32'd170452: dataIn1 = 32'd7508
; 
32'd170453: dataIn1 = 32'd7511
; 
32'd170454: dataIn1 = 32'd8949
; 
32'd170455: dataIn1 = 32'd8972
; 
32'd170456: dataIn1 = 32'd6229
; 
32'd170457: dataIn1 = 32'd6230
; 
32'd170458: dataIn1 = 32'd7512
; 
32'd170459: dataIn1 = 32'd7513
; 
32'd170460: dataIn1 = 32'd7514
; 
32'd170461: dataIn1 = 32'd7515
; 
32'd170462: dataIn1 = 32'd7516
; 
32'd170463: dataIn1 = 32'd6228
; 
32'd170464: dataIn1 = 32'd6230
; 
32'd170465: dataIn1 = 32'd7512
; 
32'd170466: dataIn1 = 32'd7513
; 
32'd170467: dataIn1 = 32'd7514
; 
32'd170468: dataIn1 = 32'd7517
; 
32'd170469: dataIn1 = 32'd7518
; 
32'd170470: dataIn1 = 32'd6228
; 
32'd170471: dataIn1 = 32'd6229
; 
32'd170472: dataIn1 = 32'd7512
; 
32'd170473: dataIn1 = 32'd7513
; 
32'd170474: dataIn1 = 32'd7514
; 
32'd170475: dataIn1 = 32'd7519
; 
32'd170476: dataIn1 = 32'd7520
; 
32'd170477: dataIn1 = 32'd5164
; 
32'd170478: dataIn1 = 32'd6230
; 
32'd170479: dataIn1 = 32'd7512
; 
32'd170480: dataIn1 = 32'd7515
; 
32'd170481: dataIn1 = 32'd7516
; 
32'd170482: dataIn1 = 32'd7535
; 
32'd170483: dataIn1 = 32'd7538
; 
32'd170484: dataIn1 = 32'd5164
; 
32'd170485: dataIn1 = 32'd6229
; 
32'd170486: dataIn1 = 32'd7512
; 
32'd170487: dataIn1 = 32'd7515
; 
32'd170488: dataIn1 = 32'd7516
; 
32'd170489: dataIn1 = 32'd7528
; 
32'd170490: dataIn1 = 32'd7531
; 
32'd170491: dataIn1 = 32'd5165
; 
32'd170492: dataIn1 = 32'd6230
; 
32'd170493: dataIn1 = 32'd7513
; 
32'd170494: dataIn1 = 32'd7517
; 
32'd170495: dataIn1 = 32'd7518
; 
32'd170496: dataIn1 = 32'd7536
; 
32'd170497: dataIn1 = 32'd7539
; 
32'd170498: dataIn1 = 32'd5165
; 
32'd170499: dataIn1 = 32'd6228
; 
32'd170500: dataIn1 = 32'd7513
; 
32'd170501: dataIn1 = 32'd7517
; 
32'd170502: dataIn1 = 32'd7518
; 
32'd170503: dataIn1 = 32'd7522
; 
32'd170504: dataIn1 = 32'd7526
; 
32'd170505: dataIn1 = 32'd5166
; 
32'd170506: dataIn1 = 32'd6229
; 
32'd170507: dataIn1 = 32'd7514
; 
32'd170508: dataIn1 = 32'd7519
; 
32'd170509: dataIn1 = 32'd7520
; 
32'd170510: dataIn1 = 32'd7530
; 
32'd170511: dataIn1 = 32'd7534
; 
32'd170512: dataIn1 = 32'd5166
; 
32'd170513: dataIn1 = 32'd6228
; 
32'd170514: dataIn1 = 32'd7514
; 
32'd170515: dataIn1 = 32'd7519
; 
32'd170516: dataIn1 = 32'd7520
; 
32'd170517: dataIn1 = 32'd7523
; 
32'd170518: dataIn1 = 32'd7527
; 
32'd170519: dataIn1 = 32'd6231
; 
32'd170520: dataIn1 = 32'd6232
; 
32'd170521: dataIn1 = 32'd7521
; 
32'd170522: dataIn1 = 32'd7522
; 
32'd170523: dataIn1 = 32'd7523
; 
32'd170524: dataIn1 = 32'd7524
; 
32'd170525: dataIn1 = 32'd7525
; 
32'd170526: dataIn1 = 32'd6228
; 
32'd170527: dataIn1 = 32'd6232
; 
32'd170528: dataIn1 = 32'd7518
; 
32'd170529: dataIn1 = 32'd7521
; 
32'd170530: dataIn1 = 32'd7522
; 
32'd170531: dataIn1 = 32'd7523
; 
32'd170532: dataIn1 = 32'd7526
; 
32'd170533: dataIn1 = 32'd6228
; 
32'd170534: dataIn1 = 32'd6231
; 
32'd170535: dataIn1 = 32'd7520
; 
32'd170536: dataIn1 = 32'd7521
; 
32'd170537: dataIn1 = 32'd7522
; 
32'd170538: dataIn1 = 32'd7523
; 
32'd170539: dataIn1 = 32'd7527
; 
32'd170540: dataIn1 = 32'd1108
; 
32'd170541: dataIn1 = 32'd6232
; 
32'd170542: dataIn1 = 32'd7521
; 
32'd170543: dataIn1 = 32'd7524
; 
32'd170544: dataIn1 = 32'd7525
; 
32'd170545: dataIn1 = 32'd7568
; 
32'd170546: dataIn1 = 32'd7571
; 
32'd170547: dataIn1 = 32'd1108
; 
32'd170548: dataIn1 = 32'd6231
; 
32'd170549: dataIn1 = 32'd7521
; 
32'd170550: dataIn1 = 32'd7524
; 
32'd170551: dataIn1 = 32'd7525
; 
32'd170552: dataIn1 = 32'd7590
; 
32'd170553: dataIn1 = 32'd7593
; 
32'd170554: dataIn1 = 32'd5165
; 
32'd170555: dataIn1 = 32'd6232
; 
32'd170556: dataIn1 = 32'd7518
; 
32'd170557: dataIn1 = 32'd7522
; 
32'd170558: dataIn1 = 32'd7526
; 
32'd170559: dataIn1 = 32'd7565
; 
32'd170560: dataIn1 = 32'd7569
; 
32'd170561: dataIn1 = 32'd5166
; 
32'd170562: dataIn1 = 32'd6231
; 
32'd170563: dataIn1 = 32'd7520
; 
32'd170564: dataIn1 = 32'd7523
; 
32'd170565: dataIn1 = 32'd7527
; 
32'd170566: dataIn1 = 32'd7589
; 
32'd170567: dataIn1 = 32'd7592
; 
32'd170568: dataIn1 = 32'd6229
; 
32'd170569: dataIn1 = 32'd6234
; 
32'd170570: dataIn1 = 32'd7516
; 
32'd170571: dataIn1 = 32'd7528
; 
32'd170572: dataIn1 = 32'd7529
; 
32'd170573: dataIn1 = 32'd7530
; 
32'd170574: dataIn1 = 32'd7531
; 
32'd170575: dataIn1 = 32'd6233
; 
32'd170576: dataIn1 = 32'd6234
; 
32'd170577: dataIn1 = 32'd7528
; 
32'd170578: dataIn1 = 32'd7529
; 
32'd170579: dataIn1 = 32'd7530
; 
32'd170580: dataIn1 = 32'd7532
; 
32'd170581: dataIn1 = 32'd7533
; 
32'd170582: dataIn1 = 32'd6229
; 
32'd170583: dataIn1 = 32'd6233
; 
32'd170584: dataIn1 = 32'd7519
; 
32'd170585: dataIn1 = 32'd7528
; 
32'd170586: dataIn1 = 32'd7529
; 
32'd170587: dataIn1 = 32'd7530
; 
32'd170588: dataIn1 = 32'd7534
; 
32'd170589: dataIn1 = 32'd5164
; 
32'd170590: dataIn1 = 32'd6234
; 
32'd170591: dataIn1 = 32'd7516
; 
32'd170592: dataIn1 = 32'd7528
; 
32'd170593: dataIn1 = 32'd7531
; 
32'd170594: dataIn1 = 32'd7546
; 
32'd170595: dataIn1 = 32'd7551
; 
32'd170596: dataIn1 = 32'd2708
; 
32'd170597: dataIn1 = 32'd6234
; 
32'd170598: dataIn1 = 32'd7529
; 
32'd170599: dataIn1 = 32'd7532
; 
32'd170600: dataIn1 = 32'd7533
; 
32'd170601: dataIn1 = 32'd7552
; 
32'd170602: dataIn1 = 32'd7554
; 
32'd170603: dataIn1 = 32'd2708
; 
32'd170604: dataIn1 = 32'd6233
; 
32'd170605: dataIn1 = 32'd7529
; 
32'd170606: dataIn1 = 32'd7532
; 
32'd170607: dataIn1 = 32'd7533
; 
32'd170608: dataIn1 = 32'd7596
; 
32'd170609: dataIn1 = 32'd7599
; 
32'd170610: dataIn1 = 32'd5166
; 
32'd170611: dataIn1 = 32'd6233
; 
32'd170612: dataIn1 = 32'd7519
; 
32'd170613: dataIn1 = 32'd7530
; 
32'd170614: dataIn1 = 32'd7534
; 
32'd170615: dataIn1 = 32'd7588
; 
32'd170616: dataIn1 = 32'd7597
; 
32'd170617: dataIn1 = 32'd6230
; 
32'd170618: dataIn1 = 32'd6236
; 
32'd170619: dataIn1 = 32'd7515
; 
32'd170620: dataIn1 = 32'd7535
; 
32'd170621: dataIn1 = 32'd7536
; 
32'd170622: dataIn1 = 32'd7537
; 
32'd170623: dataIn1 = 32'd7538
; 
32'd170624: dataIn1 = 32'd6230
; 
32'd170625: dataIn1 = 32'd6235
; 
32'd170626: dataIn1 = 32'd7517
; 
32'd170627: dataIn1 = 32'd7535
; 
32'd170628: dataIn1 = 32'd7536
; 
32'd170629: dataIn1 = 32'd7537
; 
32'd170630: dataIn1 = 32'd7539
; 
32'd170631: dataIn1 = 32'd6235
; 
32'd170632: dataIn1 = 32'd6236
; 
32'd170633: dataIn1 = 32'd7535
; 
32'd170634: dataIn1 = 32'd7536
; 
32'd170635: dataIn1 = 32'd7537
; 
32'd170636: dataIn1 = 32'd7540
; 
32'd170637: dataIn1 = 32'd7541
; 
32'd170638: dataIn1 = 32'd5164
; 
32'd170639: dataIn1 = 32'd6236
; 
32'd170640: dataIn1 = 32'd7515
; 
32'd170641: dataIn1 = 32'd7535
; 
32'd170642: dataIn1 = 32'd7538
; 
32'd170643: dataIn1 = 32'd7545
; 
32'd170644: dataIn1 = 32'd7556
; 
32'd170645: dataIn1 = 32'd5165
; 
32'd170646: dataIn1 = 32'd6235
; 
32'd170647: dataIn1 = 32'd7517
; 
32'd170648: dataIn1 = 32'd7536
; 
32'd170649: dataIn1 = 32'd7539
; 
32'd170650: dataIn1 = 32'd7564
; 
32'd170651: dataIn1 = 32'd7579
; 
32'd170652: dataIn1 = 32'd2706
; 
32'd170653: dataIn1 = 32'd6236
; 
32'd170654: dataIn1 = 32'd7385
; 
32'd170655: dataIn1 = 32'd7537
; 
32'd170656: dataIn1 = 32'd7540
; 
32'd170657: dataIn1 = 32'd7541
; 
32'd170658: dataIn1 = 32'd7558
; 
32'd170659: dataIn1 = 32'd2706
; 
32'd170660: dataIn1 = 32'd6235
; 
32'd170661: dataIn1 = 32'd7411
; 
32'd170662: dataIn1 = 32'd7537
; 
32'd170663: dataIn1 = 32'd7540
; 
32'd170664: dataIn1 = 32'd7541
; 
32'd170665: dataIn1 = 32'd7580
; 
32'd170666: dataIn1 = 32'd6238
; 
32'd170667: dataIn1 = 32'd6239
; 
32'd170668: dataIn1 = 32'd7542
; 
32'd170669: dataIn1 = 32'd7543
; 
32'd170670: dataIn1 = 32'd7544
; 
32'd170671: dataIn1 = 32'd7545
; 
32'd170672: dataIn1 = 32'd7546
; 
32'd170673: dataIn1 = 32'd6237
; 
32'd170674: dataIn1 = 32'd6239
; 
32'd170675: dataIn1 = 32'd7542
; 
32'd170676: dataIn1 = 32'd7543
; 
32'd170677: dataIn1 = 32'd7544
; 
32'd170678: dataIn1 = 32'd7547
; 
32'd170679: dataIn1 = 32'd7548
; 
32'd170680: dataIn1 = 32'd6237
; 
32'd170681: dataIn1 = 32'd6238
; 
32'd170682: dataIn1 = 32'd7542
; 
32'd170683: dataIn1 = 32'd7543
; 
32'd170684: dataIn1 = 32'd7544
; 
32'd170685: dataIn1 = 32'd7549
; 
32'd170686: dataIn1 = 32'd7550
; 
32'd170687: dataIn1 = 32'd5164
; 
32'd170688: dataIn1 = 32'd6239
; 
32'd170689: dataIn1 = 32'd7538
; 
32'd170690: dataIn1 = 32'd7542
; 
32'd170691: dataIn1 = 32'd7545
; 
32'd170692: dataIn1 = 32'd7546
; 
32'd170693: dataIn1 = 32'd7556
; 
32'd170694: dataIn1 = 32'd5164
; 
32'd170695: dataIn1 = 32'd6238
; 
32'd170696: dataIn1 = 32'd7531
; 
32'd170697: dataIn1 = 32'd7542
; 
32'd170698: dataIn1 = 32'd7545
; 
32'd170699: dataIn1 = 32'd7546
; 
32'd170700: dataIn1 = 32'd7551
; 
32'd170701: dataIn1 = 32'd5153
; 
32'd170702: dataIn1 = 32'd6239
; 
32'd170703: dataIn1 = 32'd7384
; 
32'd170704: dataIn1 = 32'd7543
; 
32'd170705: dataIn1 = 32'd7547
; 
32'd170706: dataIn1 = 32'd7548
; 
32'd170707: dataIn1 = 32'd7557
; 
32'd170708: dataIn1 = 32'd5153
; 
32'd170709: dataIn1 = 32'd6237
; 
32'd170710: dataIn1 = 32'd6753
; 
32'd170711: dataIn1 = 32'd7543
; 
32'd170712: dataIn1 = 32'd7547
; 
32'd170713: dataIn1 = 32'd7548
; 
32'd170714: dataIn1 = 32'd5167
; 
32'd170715: dataIn1 = 32'd6238
; 
32'd170716: dataIn1 = 32'd7544
; 
32'd170717: dataIn1 = 32'd7549
; 
32'd170718: dataIn1 = 32'd7550
; 
32'd170719: dataIn1 = 32'd7553
; 
32'd170720: dataIn1 = 32'd7555
; 
32'd170721: dataIn1 = 32'd5167
; 
32'd170722: dataIn1 = 32'd6237
; 
32'd170723: dataIn1 = 32'd6752
; 
32'd170724: dataIn1 = 32'd7544
; 
32'd170725: dataIn1 = 32'd7549
; 
32'd170726: dataIn1 = 32'd7550
; 
32'd170727: dataIn1 = 32'd6234
; 
32'd170728: dataIn1 = 32'd6238
; 
32'd170729: dataIn1 = 32'd7531
; 
32'd170730: dataIn1 = 32'd7546
; 
32'd170731: dataIn1 = 32'd7551
; 
32'd170732: dataIn1 = 32'd7552
; 
32'd170733: dataIn1 = 32'd7553
; 
32'd170734: dataIn1 = 32'd6234
; 
32'd170735: dataIn1 = 32'd6240
; 
32'd170736: dataIn1 = 32'd7532
; 
32'd170737: dataIn1 = 32'd7551
; 
32'd170738: dataIn1 = 32'd7552
; 
32'd170739: dataIn1 = 32'd7553
; 
32'd170740: dataIn1 = 32'd7554
; 
32'd170741: dataIn1 = 32'd6238
; 
32'd170742: dataIn1 = 32'd6240
; 
32'd170743: dataIn1 = 32'd7549
; 
32'd170744: dataIn1 = 32'd7551
; 
32'd170745: dataIn1 = 32'd7552
; 
32'd170746: dataIn1 = 32'd7553
; 
32'd170747: dataIn1 = 32'd7555
; 
32'd170748: dataIn1 = 32'd2708
; 
32'd170749: dataIn1 = 32'd6240
; 
32'd170750: dataIn1 = 32'd7532
; 
32'd170751: dataIn1 = 32'd7552
; 
32'd170752: dataIn1 = 32'd7554
; 
32'd170753: dataIn1 = 32'd8990
; 
32'd170754: dataIn1 = 32'd9023
; 
32'd170755: dataIn1 = 32'd5167
; 
32'd170756: dataIn1 = 32'd6240
; 
32'd170757: dataIn1 = 32'd7549
; 
32'd170758: dataIn1 = 32'd7553
; 
32'd170759: dataIn1 = 32'd7555
; 
32'd170760: dataIn1 = 32'd9022
; 
32'd170761: dataIn1 = 32'd9025
; 
32'd170762: dataIn1 = 32'd6236
; 
32'd170763: dataIn1 = 32'd6239
; 
32'd170764: dataIn1 = 32'd7538
; 
32'd170765: dataIn1 = 32'd7545
; 
32'd170766: dataIn1 = 32'd7556
; 
32'd170767: dataIn1 = 32'd7557
; 
32'd170768: dataIn1 = 32'd7558
; 
32'd170769: dataIn1 = 32'd6196
; 
32'd170770: dataIn1 = 32'd6239
; 
32'd170771: dataIn1 = 32'd7384
; 
32'd170772: dataIn1 = 32'd7547
; 
32'd170773: dataIn1 = 32'd7556
; 
32'd170774: dataIn1 = 32'd7557
; 
32'd170775: dataIn1 = 32'd7558
; 
32'd170776: dataIn1 = 32'd6196
; 
32'd170777: dataIn1 = 32'd6236
; 
32'd170778: dataIn1 = 32'd7385
; 
32'd170779: dataIn1 = 32'd7540
; 
32'd170780: dataIn1 = 32'd7556
; 
32'd170781: dataIn1 = 32'd7557
; 
32'd170782: dataIn1 = 32'd7558
; 
32'd170783: dataIn1 = 32'd6242
; 
32'd170784: dataIn1 = 32'd6243
; 
32'd170785: dataIn1 = 32'd7559
; 
32'd170786: dataIn1 = 32'd7560
; 
32'd170787: dataIn1 = 32'd7561
; 
32'd170788: dataIn1 = 32'd7562
; 
32'd170789: dataIn1 = 32'd7563
; 
32'd170790: dataIn1 = 32'd6241
; 
32'd170791: dataIn1 = 32'd6243
; 
32'd170792: dataIn1 = 32'd7559
; 
32'd170793: dataIn1 = 32'd7560
; 
32'd170794: dataIn1 = 32'd7561
; 
32'd170795: dataIn1 = 32'd7564
; 
32'd170796: dataIn1 = 32'd7565
; 
32'd170797: dataIn1 = 32'd6241
; 
32'd170798: dataIn1 = 32'd6242
; 
32'd170799: dataIn1 = 32'd7559
; 
32'd170800: dataIn1 = 32'd7560
; 
32'd170801: dataIn1 = 32'd7561
; 
32'd170802: dataIn1 = 32'd7566
; 
32'd170803: dataIn1 = 32'd7567
; 
32'd170804: dataIn1 = 32'd5155
; 
32'd170805: dataIn1 = 32'd6243
; 
32'd170806: dataIn1 = 32'd7410
; 
32'd170807: dataIn1 = 32'd7559
; 
32'd170808: dataIn1 = 32'd7562
; 
32'd170809: dataIn1 = 32'd7563
; 
32'd170810: dataIn1 = 32'd7578
; 
32'd170811: dataIn1 = 32'd5155
; 
32'd170812: dataIn1 = 32'd6242
; 
32'd170813: dataIn1 = 32'd7403
; 
32'd170814: dataIn1 = 32'd7559
; 
32'd170815: dataIn1 = 32'd7562
; 
32'd170816: dataIn1 = 32'd7563
; 
32'd170817: dataIn1 = 32'd7573
; 
32'd170818: dataIn1 = 32'd5165
; 
32'd170819: dataIn1 = 32'd6243
; 
32'd170820: dataIn1 = 32'd7539
; 
32'd170821: dataIn1 = 32'd7560
; 
32'd170822: dataIn1 = 32'd7564
; 
32'd170823: dataIn1 = 32'd7565
; 
32'd170824: dataIn1 = 32'd7579
; 
32'd170825: dataIn1 = 32'd5165
; 
32'd170826: dataIn1 = 32'd6241
; 
32'd170827: dataIn1 = 32'd7526
; 
32'd170828: dataIn1 = 32'd7560
; 
32'd170829: dataIn1 = 32'd7564
; 
32'd170830: dataIn1 = 32'd7565
; 
32'd170831: dataIn1 = 32'd7569
; 
32'd170832: dataIn1 = 32'd2640
; 
32'd170833: dataIn1 = 32'd6242
; 
32'd170834: dataIn1 = 32'd7561
; 
32'd170835: dataIn1 = 32'd7566
; 
32'd170836: dataIn1 = 32'd7567
; 
32'd170837: dataIn1 = 32'd7575
; 
32'd170838: dataIn1 = 32'd7577
; 
32'd170839: dataIn1 = 32'd2640
; 
32'd170840: dataIn1 = 32'd6241
; 
32'd170841: dataIn1 = 32'd7561
; 
32'd170842: dataIn1 = 32'd7566
; 
32'd170843: dataIn1 = 32'd7567
; 
32'd170844: dataIn1 = 32'd7570
; 
32'd170845: dataIn1 = 32'd7572
; 
32'd170846: dataIn1 = 32'd4916
; 
32'd170847: dataIn1 = 32'd6232
; 
32'd170848: dataIn1 = 32'd7524
; 
32'd170849: dataIn1 = 32'd7568
; 
32'd170850: dataIn1 = 32'd7569
; 
32'd170851: dataIn1 = 32'd7570
; 
32'd170852: dataIn1 = 32'd7571
; 
32'd170853: dataIn1 = 32'd6232
; 
32'd170854: dataIn1 = 32'd6241
; 
32'd170855: dataIn1 = 32'd7526
; 
32'd170856: dataIn1 = 32'd7565
; 
32'd170857: dataIn1 = 32'd7568
; 
32'd170858: dataIn1 = 32'd7569
; 
32'd170859: dataIn1 = 32'd7570
; 
32'd170860: dataIn1 = 32'd4916
; 
32'd170861: dataIn1 = 32'd6241
; 
32'd170862: dataIn1 = 32'd7567
; 
32'd170863: dataIn1 = 32'd7568
; 
32'd170864: dataIn1 = 32'd7569
; 
32'd170865: dataIn1 = 32'd7570
; 
32'd170866: dataIn1 = 32'd7572
; 
32'd170867: dataIn1 = 32'd1108
; 
32'd170868: dataIn1 = 32'd4916
; 
32'd170869: dataIn1 = 32'd7524
; 
32'd170870: dataIn1 = 32'd7568
; 
32'd170871: dataIn1 = 32'd7571
; 
32'd170872: dataIn1 = 32'd9623
; 
32'd170873: dataIn1 = 32'd9633
; 
32'd170874: dataIn1 = 32'd2640
; 
32'd170875: dataIn1 = 32'd4916
; 
32'd170876: dataIn1 = 32'd7567
; 
32'd170877: dataIn1 = 32'd7570
; 
32'd170878: dataIn1 = 32'd7572
; 
32'd170879: dataIn1 = 32'd9626
; 
32'd170880: dataIn1 = 32'd9634
; 
32'd170881: dataIn1 = 32'd6203
; 
32'd170882: dataIn1 = 32'd6242
; 
32'd170883: dataIn1 = 32'd7403
; 
32'd170884: dataIn1 = 32'd7563
; 
32'd170885: dataIn1 = 32'd7573
; 
32'd170886: dataIn1 = 32'd7574
; 
32'd170887: dataIn1 = 32'd7575
; 
32'd170888: dataIn1 = 32'd4915
; 
32'd170889: dataIn1 = 32'd6203
; 
32'd170890: dataIn1 = 32'd7404
; 
32'd170891: dataIn1 = 32'd7573
; 
32'd170892: dataIn1 = 32'd7574
; 
32'd170893: dataIn1 = 32'd7575
; 
32'd170894: dataIn1 = 32'd7576
; 
32'd170895: dataIn1 = 32'd4915
; 
32'd170896: dataIn1 = 32'd6242
; 
32'd170897: dataIn1 = 32'd7566
; 
32'd170898: dataIn1 = 32'd7573
; 
32'd170899: dataIn1 = 32'd7574
; 
32'd170900: dataIn1 = 32'd7575
; 
32'd170901: dataIn1 = 32'd7577
; 
32'd170902: dataIn1 = 32'd133
; 
32'd170903: dataIn1 = 32'd4915
; 
32'd170904: dataIn1 = 32'd7404
; 
32'd170905: dataIn1 = 32'd7574
; 
32'd170906: dataIn1 = 32'd7576
; 
32'd170907: dataIn1 = 32'd9603
; 
32'd170908: dataIn1 = 32'd9629
; 
32'd170909: dataIn1 = 32'd2640
; 
32'd170910: dataIn1 = 32'd4915
; 
32'd170911: dataIn1 = 32'd7566
; 
32'd170912: dataIn1 = 32'd7575
; 
32'd170913: dataIn1 = 32'd7577
; 
32'd170914: dataIn1 = 32'd9627
; 
32'd170915: dataIn1 = 32'd9631
; 
32'd170916: dataIn1 = 32'd6204
; 
32'd170917: dataIn1 = 32'd6243
; 
32'd170918: dataIn1 = 32'd7410
; 
32'd170919: dataIn1 = 32'd7562
; 
32'd170920: dataIn1 = 32'd7578
; 
32'd170921: dataIn1 = 32'd7579
; 
32'd170922: dataIn1 = 32'd7580
; 
32'd170923: dataIn1 = 32'd6235
; 
32'd170924: dataIn1 = 32'd6243
; 
32'd170925: dataIn1 = 32'd7539
; 
32'd170926: dataIn1 = 32'd7564
; 
32'd170927: dataIn1 = 32'd7578
; 
32'd170928: dataIn1 = 32'd7579
; 
32'd170929: dataIn1 = 32'd7580
; 
32'd170930: dataIn1 = 32'd6204
; 
32'd170931: dataIn1 = 32'd6235
; 
32'd170932: dataIn1 = 32'd7411
; 
32'd170933: dataIn1 = 32'd7541
; 
32'd170934: dataIn1 = 32'd7578
; 
32'd170935: dataIn1 = 32'd7579
; 
32'd170936: dataIn1 = 32'd7580
; 
32'd170937: dataIn1 = 32'd6245
; 
32'd170938: dataIn1 = 32'd6246
; 
32'd170939: dataIn1 = 32'd7581
; 
32'd170940: dataIn1 = 32'd7582
; 
32'd170941: dataIn1 = 32'd7583
; 
32'd170942: dataIn1 = 32'd7584
; 
32'd170943: dataIn1 = 32'd7585
; 
32'd170944: dataIn1 = 32'd6244
; 
32'd170945: dataIn1 = 32'd6246
; 
32'd170946: dataIn1 = 32'd7581
; 
32'd170947: dataIn1 = 32'd7582
; 
32'd170948: dataIn1 = 32'd7583
; 
32'd170949: dataIn1 = 32'd7586
; 
32'd170950: dataIn1 = 32'd7587
; 
32'd170951: dataIn1 = 32'd6244
; 
32'd170952: dataIn1 = 32'd6245
; 
32'd170953: dataIn1 = 32'd7581
; 
32'd170954: dataIn1 = 32'd7582
; 
32'd170955: dataIn1 = 32'd7583
; 
32'd170956: dataIn1 = 32'd7588
; 
32'd170957: dataIn1 = 32'd7589
; 
32'd170958: dataIn1 = 32'd5168
; 
32'd170959: dataIn1 = 32'd6246
; 
32'd170960: dataIn1 = 32'd7581
; 
32'd170961: dataIn1 = 32'd7584
; 
32'd170962: dataIn1 = 32'd7585
; 
32'd170963: dataIn1 = 32'd7600
; 
32'd170964: dataIn1 = 32'd7603
; 
32'd170965: dataIn1 = 32'd5168
; 
32'd170966: dataIn1 = 32'd6245
; 
32'd170967: dataIn1 = 32'd7581
; 
32'd170968: dataIn1 = 32'd7584
; 
32'd170969: dataIn1 = 32'd7585
; 
32'd170970: dataIn1 = 32'd7595
; 
32'd170971: dataIn1 = 32'd7598
; 
32'd170972: dataIn1 = 32'd2641
; 
32'd170973: dataIn1 = 32'd6246
; 
32'd170974: dataIn1 = 32'd7582
; 
32'd170975: dataIn1 = 32'd7586
; 
32'd170976: dataIn1 = 32'd7587
; 
32'd170977: dataIn1 = 32'd7601
; 
32'd170978: dataIn1 = 32'd7604
; 
32'd170979: dataIn1 = 32'd2641
; 
32'd170980: dataIn1 = 32'd6244
; 
32'd170981: dataIn1 = 32'd7582
; 
32'd170982: dataIn1 = 32'd7586
; 
32'd170983: dataIn1 = 32'd7587
; 
32'd170984: dataIn1 = 32'd7591
; 
32'd170985: dataIn1 = 32'd7594
; 
32'd170986: dataIn1 = 32'd5166
; 
32'd170987: dataIn1 = 32'd6245
; 
32'd170988: dataIn1 = 32'd7534
; 
32'd170989: dataIn1 = 32'd7583
; 
32'd170990: dataIn1 = 32'd7588
; 
32'd170991: dataIn1 = 32'd7589
; 
32'd170992: dataIn1 = 32'd7597
; 
32'd170993: dataIn1 = 32'd5166
; 
32'd170994: dataIn1 = 32'd6244
; 
32'd170995: dataIn1 = 32'd7527
; 
32'd170996: dataIn1 = 32'd7583
; 
32'd170997: dataIn1 = 32'd7588
; 
32'd170998: dataIn1 = 32'd7589
; 
32'd170999: dataIn1 = 32'd7592
; 
32'd171000: dataIn1 = 32'd4920
; 
32'd171001: dataIn1 = 32'd6231
; 
32'd171002: dataIn1 = 32'd7525
; 
32'd171003: dataIn1 = 32'd7590
; 
32'd171004: dataIn1 = 32'd7591
; 
32'd171005: dataIn1 = 32'd7592
; 
32'd171006: dataIn1 = 32'd7593
; 
32'd171007: dataIn1 = 32'd4920
; 
32'd171008: dataIn1 = 32'd6244
; 
32'd171009: dataIn1 = 32'd7587
; 
32'd171010: dataIn1 = 32'd7590
; 
32'd171011: dataIn1 = 32'd7591
; 
32'd171012: dataIn1 = 32'd7592
; 
32'd171013: dataIn1 = 32'd7594
; 
32'd171014: dataIn1 = 32'd6231
; 
32'd171015: dataIn1 = 32'd6244
; 
32'd171016: dataIn1 = 32'd7527
; 
32'd171017: dataIn1 = 32'd7589
; 
32'd171018: dataIn1 = 32'd7590
; 
32'd171019: dataIn1 = 32'd7591
; 
32'd171020: dataIn1 = 32'd7592
; 
32'd171021: dataIn1 = 32'd1108
; 
32'd171022: dataIn1 = 32'd4920
; 
32'd171023: dataIn1 = 32'd7525
; 
32'd171024: dataIn1 = 32'd7590
; 
32'd171025: dataIn1 = 32'd7593
; 
32'd171026: dataIn1 = 32'd9625
; 
32'd171027: dataIn1 = 32'd9639
; 
32'd171028: dataIn1 = 32'd2641
; 
32'd171029: dataIn1 = 32'd4920
; 
32'd171030: dataIn1 = 32'd7587
; 
32'd171031: dataIn1 = 32'd7591
; 
32'd171032: dataIn1 = 32'd7594
; 
32'd171033: dataIn1 = 32'd9637
; 
32'd171034: dataIn1 = 32'd9638
; 
32'd171035: dataIn1 = 32'd6245
; 
32'd171036: dataIn1 = 32'd6247
; 
32'd171037: dataIn1 = 32'd7585
; 
32'd171038: dataIn1 = 32'd7595
; 
32'd171039: dataIn1 = 32'd7596
; 
32'd171040: dataIn1 = 32'd7597
; 
32'd171041: dataIn1 = 32'd7598
; 
32'd171042: dataIn1 = 32'd6233
; 
32'd171043: dataIn1 = 32'd6247
; 
32'd171044: dataIn1 = 32'd7533
; 
32'd171045: dataIn1 = 32'd7595
; 
32'd171046: dataIn1 = 32'd7596
; 
32'd171047: dataIn1 = 32'd7597
; 
32'd171048: dataIn1 = 32'd7599
; 
32'd171049: dataIn1 = 32'd6233
; 
32'd171050: dataIn1 = 32'd6245
; 
32'd171051: dataIn1 = 32'd7534
; 
32'd171052: dataIn1 = 32'd7588
; 
32'd171053: dataIn1 = 32'd7595
; 
32'd171054: dataIn1 = 32'd7596
; 
32'd171055: dataIn1 = 32'd7597
; 
32'd171056: dataIn1 = 32'd5168
; 
32'd171057: dataIn1 = 32'd6247
; 
32'd171058: dataIn1 = 32'd7585
; 
32'd171059: dataIn1 = 32'd7595
; 
32'd171060: dataIn1 = 32'd7598
; 
32'd171061: dataIn1 = 32'd9006
; 
32'd171062: dataIn1 = 32'd9013
; 
32'd171063: dataIn1 = 32'd2708
; 
32'd171064: dataIn1 = 32'd6247
; 
32'd171065: dataIn1 = 32'd7533
; 
32'd171066: dataIn1 = 32'd7596
; 
32'd171067: dataIn1 = 32'd7599
; 
32'd171068: dataIn1 = 32'd8989
; 
32'd171069: dataIn1 = 32'd9012
; 
32'd171070: dataIn1 = 32'd6246
; 
32'd171071: dataIn1 = 32'd6248
; 
32'd171072: dataIn1 = 32'd7584
; 
32'd171073: dataIn1 = 32'd7600
; 
32'd171074: dataIn1 = 32'd7601
; 
32'd171075: dataIn1 = 32'd7602
; 
32'd171076: dataIn1 = 32'd7603
; 
32'd171077: dataIn1 = 32'd4921
; 
32'd171078: dataIn1 = 32'd6246
; 
32'd171079: dataIn1 = 32'd7586
; 
32'd171080: dataIn1 = 32'd7600
; 
32'd171081: dataIn1 = 32'd7601
; 
32'd171082: dataIn1 = 32'd7602
; 
32'd171083: dataIn1 = 32'd7604
; 
32'd171084: dataIn1 = 32'd4921
; 
32'd171085: dataIn1 = 32'd6248
; 
32'd171086: dataIn1 = 32'd7600
; 
32'd171087: dataIn1 = 32'd7601
; 
32'd171088: dataIn1 = 32'd7602
; 
32'd171089: dataIn1 = 32'd7605
; 
32'd171090: dataIn1 = 32'd7606
; 
32'd171091: dataIn1 = 32'd5168
; 
32'd171092: dataIn1 = 32'd6248
; 
32'd171093: dataIn1 = 32'd7584
; 
32'd171094: dataIn1 = 32'd7600
; 
32'd171095: dataIn1 = 32'd7603
; 
32'd171096: dataIn1 = 32'd9007
; 
32'd171097: dataIn1 = 32'd9010
; 
32'd171098: dataIn1 = 32'd2641
; 
32'd171099: dataIn1 = 32'd4921
; 
32'd171100: dataIn1 = 32'd7586
; 
32'd171101: dataIn1 = 32'd7601
; 
32'd171102: dataIn1 = 32'd7604
; 
32'd171103: dataIn1 = 32'd9636
; 
32'd171104: dataIn1 = 32'd9641
; 
32'd171105: dataIn1 = 32'd7
; 
32'd171106: dataIn1 = 32'd6248
; 
32'd171107: dataIn1 = 32'd7602
; 
32'd171108: dataIn1 = 32'd7605
; 
32'd171109: dataIn1 = 32'd7606
; 
32'd171110: dataIn1 = 32'd7713
; 
32'd171111: dataIn1 = 32'd9008
; 
32'd171112: dataIn1 = 32'd7
; 
32'd171113: dataIn1 = 32'd4921
; 
32'd171114: dataIn1 = 32'd7602
; 
32'd171115: dataIn1 = 32'd7605
; 
32'd171116: dataIn1 = 32'd7606
; 
32'd171117: dataIn1 = 32'd9607
; 
32'd171118: dataIn1 = 32'd9643
; 
32'd171119: dataIn1 = 32'd6250
; 
32'd171120: dataIn1 = 32'd6251
; 
32'd171121: dataIn1 = 32'd7607
; 
32'd171122: dataIn1 = 32'd7608
; 
32'd171123: dataIn1 = 32'd7609
; 
32'd171124: dataIn1 = 32'd7610
; 
32'd171125: dataIn1 = 32'd7611
; 
32'd171126: dataIn1 = 32'd6249
; 
32'd171127: dataIn1 = 32'd6251
; 
32'd171128: dataIn1 = 32'd7607
; 
32'd171129: dataIn1 = 32'd7608
; 
32'd171130: dataIn1 = 32'd7609
; 
32'd171131: dataIn1 = 32'd7612
; 
32'd171132: dataIn1 = 32'd7613
; 
32'd171133: dataIn1 = 32'd6249
; 
32'd171134: dataIn1 = 32'd6250
; 
32'd171135: dataIn1 = 32'd7607
; 
32'd171136: dataIn1 = 32'd7608
; 
32'd171137: dataIn1 = 32'd7609
; 
32'd171138: dataIn1 = 32'd7614
; 
32'd171139: dataIn1 = 32'd7615
; 
32'd171140: dataIn1 = 32'd5169
; 
32'd171141: dataIn1 = 32'd6251
; 
32'd171142: dataIn1 = 32'd7607
; 
32'd171143: dataIn1 = 32'd7610
; 
32'd171144: dataIn1 = 32'd7611
; 
32'd171145: dataIn1 = 32'd7623
; 
32'd171146: dataIn1 = 32'd7626
; 
32'd171147: dataIn1 = 32'd5169
; 
32'd171148: dataIn1 = 32'd6250
; 
32'd171149: dataIn1 = 32'd6755
; 
32'd171150: dataIn1 = 32'd7607
; 
32'd171151: dataIn1 = 32'd7610
; 
32'd171152: dataIn1 = 32'd7611
; 
32'd171153: dataIn1 = 32'd5170
; 
32'd171154: dataIn1 = 32'd6251
; 
32'd171155: dataIn1 = 32'd7608
; 
32'd171156: dataIn1 = 32'd7612
; 
32'd171157: dataIn1 = 32'd7613
; 
32'd171158: dataIn1 = 32'd7624
; 
32'd171159: dataIn1 = 32'd7627
; 
32'd171160: dataIn1 = 32'd5170
; 
32'd171161: dataIn1 = 32'd6249
; 
32'd171162: dataIn1 = 32'd7608
; 
32'd171163: dataIn1 = 32'd7612
; 
32'd171164: dataIn1 = 32'd7613
; 
32'd171165: dataIn1 = 32'd7617
; 
32'd171166: dataIn1 = 32'd7621
; 
32'd171167: dataIn1 = 32'd5171
; 
32'd171168: dataIn1 = 32'd6250
; 
32'd171169: dataIn1 = 32'd6754
; 
32'd171170: dataIn1 = 32'd7609
; 
32'd171171: dataIn1 = 32'd7614
; 
32'd171172: dataIn1 = 32'd7615
; 
32'd171173: dataIn1 = 32'd5171
; 
32'd171174: dataIn1 = 32'd6249
; 
32'd171175: dataIn1 = 32'd7609
; 
32'd171176: dataIn1 = 32'd7614
; 
32'd171177: dataIn1 = 32'd7615
; 
32'd171178: dataIn1 = 32'd7618
; 
32'd171179: dataIn1 = 32'd7622
; 
32'd171180: dataIn1 = 32'd6252
; 
32'd171181: dataIn1 = 32'd6253
; 
32'd171182: dataIn1 = 32'd7616
; 
32'd171183: dataIn1 = 32'd7617
; 
32'd171184: dataIn1 = 32'd7618
; 
32'd171185: dataIn1 = 32'd7619
; 
32'd171186: dataIn1 = 32'd7620
; 
32'd171187: dataIn1 = 32'd6249
; 
32'd171188: dataIn1 = 32'd6253
; 
32'd171189: dataIn1 = 32'd7613
; 
32'd171190: dataIn1 = 32'd7616
; 
32'd171191: dataIn1 = 32'd7617
; 
32'd171192: dataIn1 = 32'd7618
; 
32'd171193: dataIn1 = 32'd7621
; 
32'd171194: dataIn1 = 32'd6249
; 
32'd171195: dataIn1 = 32'd6252
; 
32'd171196: dataIn1 = 32'd7615
; 
32'd171197: dataIn1 = 32'd7616
; 
32'd171198: dataIn1 = 32'd7617
; 
32'd171199: dataIn1 = 32'd7618
; 
32'd171200: dataIn1 = 32'd7622
; 
32'd171201: dataIn1 = 32'd2709
; 
32'd171202: dataIn1 = 32'd6253
; 
32'd171203: dataIn1 = 32'd7616
; 
32'd171204: dataIn1 = 32'd7619
; 
32'd171205: dataIn1 = 32'd7620
; 
32'd171206: dataIn1 = 32'd7646
; 
32'd171207: dataIn1 = 32'd7649
; 
32'd171208: dataIn1 = 32'd2709
; 
32'd171209: dataIn1 = 32'd6252
; 
32'd171210: dataIn1 = 32'd7616
; 
32'd171211: dataIn1 = 32'd7619
; 
32'd171212: dataIn1 = 32'd7620
; 
32'd171213: dataIn1 = 32'd7663
; 
32'd171214: dataIn1 = 32'd7666
; 
32'd171215: dataIn1 = 32'd5170
; 
32'd171216: dataIn1 = 32'd6253
; 
32'd171217: dataIn1 = 32'd7613
; 
32'd171218: dataIn1 = 32'd7617
; 
32'd171219: dataIn1 = 32'd7621
; 
32'd171220: dataIn1 = 32'd7643
; 
32'd171221: dataIn1 = 32'd7647
; 
32'd171222: dataIn1 = 32'd5171
; 
32'd171223: dataIn1 = 32'd6252
; 
32'd171224: dataIn1 = 32'd7615
; 
32'd171225: dataIn1 = 32'd7618
; 
32'd171226: dataIn1 = 32'd7622
; 
32'd171227: dataIn1 = 32'd7665
; 
32'd171228: dataIn1 = 32'd7669
; 
32'd171229: dataIn1 = 32'd6251
; 
32'd171230: dataIn1 = 32'd6255
; 
32'd171231: dataIn1 = 32'd7610
; 
32'd171232: dataIn1 = 32'd7623
; 
32'd171233: dataIn1 = 32'd7624
; 
32'd171234: dataIn1 = 32'd7625
; 
32'd171235: dataIn1 = 32'd7626
; 
32'd171236: dataIn1 = 32'd6251
; 
32'd171237: dataIn1 = 32'd6254
; 
32'd171238: dataIn1 = 32'd7612
; 
32'd171239: dataIn1 = 32'd7623
; 
32'd171240: dataIn1 = 32'd7624
; 
32'd171241: dataIn1 = 32'd7625
; 
32'd171242: dataIn1 = 32'd7627
; 
32'd171243: dataIn1 = 32'd6254
; 
32'd171244: dataIn1 = 32'd6255
; 
32'd171245: dataIn1 = 32'd7623
; 
32'd171246: dataIn1 = 32'd7624
; 
32'd171247: dataIn1 = 32'd7625
; 
32'd171248: dataIn1 = 32'd7628
; 
32'd171249: dataIn1 = 32'd7629
; 
32'd171250: dataIn1 = 32'd5169
; 
32'd171251: dataIn1 = 32'd6255
; 
32'd171252: dataIn1 = 32'd7610
; 
32'd171253: dataIn1 = 32'd7623
; 
32'd171254: dataIn1 = 32'd7626
; 
32'd171255: dataIn1 = 32'd7630
; 
32'd171256: dataIn1 = 32'd7633
; 
32'd171257: dataIn1 = 32'd5170
; 
32'd171258: dataIn1 = 32'd6254
; 
32'd171259: dataIn1 = 32'd7612
; 
32'd171260: dataIn1 = 32'd7624
; 
32'd171261: dataIn1 = 32'd7627
; 
32'd171262: dataIn1 = 32'd7642
; 
32'd171263: dataIn1 = 32'd7659
; 
32'd171264: dataIn1 = 32'd2711
; 
32'd171265: dataIn1 = 32'd6255
; 
32'd171266: dataIn1 = 32'd7625
; 
32'd171267: dataIn1 = 32'd7628
; 
32'd171268: dataIn1 = 32'd7629
; 
32'd171269: dataIn1 = 32'd7632
; 
32'd171270: dataIn1 = 32'd7636
; 
32'd171271: dataIn1 = 32'd2711
; 
32'd171272: dataIn1 = 32'd6254
; 
32'd171273: dataIn1 = 32'd7625
; 
32'd171274: dataIn1 = 32'd7628
; 
32'd171275: dataIn1 = 32'd7629
; 
32'd171276: dataIn1 = 32'd7660
; 
32'd171277: dataIn1 = 32'd7662
; 
32'd171278: dataIn1 = 32'd6255
; 
32'd171279: dataIn1 = 32'd6257
; 
32'd171280: dataIn1 = 32'd7626
; 
32'd171281: dataIn1 = 32'd7630
; 
32'd171282: dataIn1 = 32'd7631
; 
32'd171283: dataIn1 = 32'd7632
; 
32'd171284: dataIn1 = 32'd7633
; 
32'd171285: dataIn1 = 32'd6256
; 
32'd171286: dataIn1 = 32'd6257
; 
32'd171287: dataIn1 = 32'd7630
; 
32'd171288: dataIn1 = 32'd7631
; 
32'd171289: dataIn1 = 32'd7632
; 
32'd171290: dataIn1 = 32'd7634
; 
32'd171291: dataIn1 = 32'd7635
; 
32'd171292: dataIn1 = 32'd6255
; 
32'd171293: dataIn1 = 32'd6256
; 
32'd171294: dataIn1 = 32'd7628
; 
32'd171295: dataIn1 = 32'd7630
; 
32'd171296: dataIn1 = 32'd7631
; 
32'd171297: dataIn1 = 32'd7632
; 
32'd171298: dataIn1 = 32'd7636
; 
32'd171299: dataIn1 = 32'd5169
; 
32'd171300: dataIn1 = 32'd6257
; 
32'd171301: dataIn1 = 32'd6757
; 
32'd171302: dataIn1 = 32'd7626
; 
32'd171303: dataIn1 = 32'd7630
; 
32'd171304: dataIn1 = 32'd7633
; 
32'd171305: dataIn1 = 32'd5172
; 
32'd171306: dataIn1 = 32'd6257
; 
32'd171307: dataIn1 = 32'd6756
; 
32'd171308: dataIn1 = 32'd7631
; 
32'd171309: dataIn1 = 32'd7634
; 
32'd171310: dataIn1 = 32'd7635
; 
32'd171311: dataIn1 = 32'd5172
; 
32'd171312: dataIn1 = 32'd6256
; 
32'd171313: dataIn1 = 32'd7631
; 
32'd171314: dataIn1 = 32'd7634
; 
32'd171315: dataIn1 = 32'd7635
; 
32'd171316: dataIn1 = 32'd7800
; 
32'd171317: dataIn1 = 32'd7810
; 
32'd171318: dataIn1 = 32'd2711
; 
32'd171319: dataIn1 = 32'd6256
; 
32'd171320: dataIn1 = 32'd7628
; 
32'd171321: dataIn1 = 32'd7632
; 
32'd171322: dataIn1 = 32'd7636
; 
32'd171323: dataIn1 = 32'd7793
; 
32'd171324: dataIn1 = 32'd7811
; 
32'd171325: dataIn1 = 32'd6259
; 
32'd171326: dataIn1 = 32'd6260
; 
32'd171327: dataIn1 = 32'd7637
; 
32'd171328: dataIn1 = 32'd7638
; 
32'd171329: dataIn1 = 32'd7639
; 
32'd171330: dataIn1 = 32'd7640
; 
32'd171331: dataIn1 = 32'd7641
; 
32'd171332: dataIn1 = 32'd6258
; 
32'd171333: dataIn1 = 32'd6260
; 
32'd171334: dataIn1 = 32'd7637
; 
32'd171335: dataIn1 = 32'd7638
; 
32'd171336: dataIn1 = 32'd7639
; 
32'd171337: dataIn1 = 32'd7642
; 
32'd171338: dataIn1 = 32'd7643
; 
32'd171339: dataIn1 = 32'd6258
; 
32'd171340: dataIn1 = 32'd6259
; 
32'd171341: dataIn1 = 32'd7637
; 
32'd171342: dataIn1 = 32'd7638
; 
32'd171343: dataIn1 = 32'd7639
; 
32'd171344: dataIn1 = 32'd7644
; 
32'd171345: dataIn1 = 32'd7645
; 
32'd171346: dataIn1 = 32'd5174
; 
32'd171347: dataIn1 = 32'd6260
; 
32'd171348: dataIn1 = 32'd7637
; 
32'd171349: dataIn1 = 32'd7640
; 
32'd171350: dataIn1 = 32'd7641
; 
32'd171351: dataIn1 = 32'd7658
; 
32'd171352: dataIn1 = 32'd7661
; 
32'd171353: dataIn1 = 32'd5174
; 
32'd171354: dataIn1 = 32'd6259
; 
32'd171355: dataIn1 = 32'd7637
; 
32'd171356: dataIn1 = 32'd7640
; 
32'd171357: dataIn1 = 32'd7641
; 
32'd171358: dataIn1 = 32'd7651
; 
32'd171359: dataIn1 = 32'd7654
; 
32'd171360: dataIn1 = 32'd5170
; 
32'd171361: dataIn1 = 32'd6260
; 
32'd171362: dataIn1 = 32'd7627
; 
32'd171363: dataIn1 = 32'd7638
; 
32'd171364: dataIn1 = 32'd7642
; 
32'd171365: dataIn1 = 32'd7643
; 
32'd171366: dataIn1 = 32'd7659
; 
32'd171367: dataIn1 = 32'd5170
; 
32'd171368: dataIn1 = 32'd6258
; 
32'd171369: dataIn1 = 32'd7621
; 
32'd171370: dataIn1 = 32'd7638
; 
32'd171371: dataIn1 = 32'd7642
; 
32'd171372: dataIn1 = 32'd7643
; 
32'd171373: dataIn1 = 32'd7647
; 
32'd171374: dataIn1 = 32'd5175
; 
32'd171375: dataIn1 = 32'd6259
; 
32'd171376: dataIn1 = 32'd7639
; 
32'd171377: dataIn1 = 32'd7644
; 
32'd171378: dataIn1 = 32'd7645
; 
32'd171379: dataIn1 = 32'd7653
; 
32'd171380: dataIn1 = 32'd7657
; 
32'd171381: dataIn1 = 32'd5175
; 
32'd171382: dataIn1 = 32'd6258
; 
32'd171383: dataIn1 = 32'd7639
; 
32'd171384: dataIn1 = 32'd7644
; 
32'd171385: dataIn1 = 32'd7645
; 
32'd171386: dataIn1 = 32'd7648
; 
32'd171387: dataIn1 = 32'd7650
; 
32'd171388: dataIn1 = 32'd6253
; 
32'd171389: dataIn1 = 32'd6261
; 
32'd171390: dataIn1 = 32'd7619
; 
32'd171391: dataIn1 = 32'd7646
; 
32'd171392: dataIn1 = 32'd7647
; 
32'd171393: dataIn1 = 32'd7648
; 
32'd171394: dataIn1 = 32'd7649
; 
32'd171395: dataIn1 = 32'd6253
; 
32'd171396: dataIn1 = 32'd6258
; 
32'd171397: dataIn1 = 32'd7621
; 
32'd171398: dataIn1 = 32'd7643
; 
32'd171399: dataIn1 = 32'd7646
; 
32'd171400: dataIn1 = 32'd7647
; 
32'd171401: dataIn1 = 32'd7648
; 
32'd171402: dataIn1 = 32'd6258
; 
32'd171403: dataIn1 = 32'd6261
; 
32'd171404: dataIn1 = 32'd7645
; 
32'd171405: dataIn1 = 32'd7646
; 
32'd171406: dataIn1 = 32'd7647
; 
32'd171407: dataIn1 = 32'd7648
; 
32'd171408: dataIn1 = 32'd7650
; 
32'd171409: dataIn1 = 32'd2709
; 
32'd171410: dataIn1 = 32'd6261
; 
32'd171411: dataIn1 = 32'd7619
; 
32'd171412: dataIn1 = 32'd7646
; 
32'd171413: dataIn1 = 32'd7649
; 
32'd171414: dataIn1 = 32'd7682
; 
32'd171415: dataIn1 = 32'd7735
; 
32'd171416: dataIn1 = 32'd5175
; 
32'd171417: dataIn1 = 32'd6261
; 
32'd171418: dataIn1 = 32'd7645
; 
32'd171419: dataIn1 = 32'd7648
; 
32'd171420: dataIn1 = 32'd7650
; 
32'd171421: dataIn1 = 32'd7734
; 
32'd171422: dataIn1 = 32'd7737
; 
32'd171423: dataIn1 = 32'd6259
; 
32'd171424: dataIn1 = 32'd6263
; 
32'd171425: dataIn1 = 32'd7641
; 
32'd171426: dataIn1 = 32'd7651
; 
32'd171427: dataIn1 = 32'd7652
; 
32'd171428: dataIn1 = 32'd7653
; 
32'd171429: dataIn1 = 32'd7654
; 
32'd171430: dataIn1 = 32'd6262
; 
32'd171431: dataIn1 = 32'd6263
; 
32'd171432: dataIn1 = 32'd7651
; 
32'd171433: dataIn1 = 32'd7652
; 
32'd171434: dataIn1 = 32'd7653
; 
32'd171435: dataIn1 = 32'd7655
; 
32'd171436: dataIn1 = 32'd7656
; 
32'd171437: dataIn1 = 32'd6259
; 
32'd171438: dataIn1 = 32'd6262
; 
32'd171439: dataIn1 = 32'd7644
; 
32'd171440: dataIn1 = 32'd7651
; 
32'd171441: dataIn1 = 32'd7652
; 
32'd171442: dataIn1 = 32'd7653
; 
32'd171443: dataIn1 = 32'd7657
; 
32'd171444: dataIn1 = 32'd5174
; 
32'd171445: dataIn1 = 32'd6263
; 
32'd171446: dataIn1 = 32'd7641
; 
32'd171447: dataIn1 = 32'd7651
; 
32'd171448: dataIn1 = 32'd7654
; 
32'd171449: dataIn1 = 32'd7816
; 
32'd171450: dataIn1 = 32'd7826
; 
32'd171451: dataIn1 = 32'd136
; 
32'd171452: dataIn1 = 32'd6263
; 
32'd171453: dataIn1 = 32'd7652
; 
32'd171454: dataIn1 = 32'd7655
; 
32'd171455: dataIn1 = 32'd7656
; 
32'd171456: dataIn1 = 32'd7827
; 
32'd171457: dataIn1 = 32'd7829
; 
32'd171458: dataIn1 = 32'd136
; 
32'd171459: dataIn1 = 32'd6262
; 
32'd171460: dataIn1 = 32'd7652
; 
32'd171461: dataIn1 = 32'd7655
; 
32'd171462: dataIn1 = 32'd7656
; 
32'd171463: dataIn1 = 32'd7739
; 
32'd171464: dataIn1 = 32'd7742
; 
32'd171465: dataIn1 = 32'd5175
; 
32'd171466: dataIn1 = 32'd6262
; 
32'd171467: dataIn1 = 32'd7644
; 
32'd171468: dataIn1 = 32'd7653
; 
32'd171469: dataIn1 = 32'd7657
; 
32'd171470: dataIn1 = 32'd7733
; 
32'd171471: dataIn1 = 32'd7740
; 
32'd171472: dataIn1 = 32'd6260
; 
32'd171473: dataIn1 = 32'd6264
; 
32'd171474: dataIn1 = 32'd7640
; 
32'd171475: dataIn1 = 32'd7658
; 
32'd171476: dataIn1 = 32'd7659
; 
32'd171477: dataIn1 = 32'd7660
; 
32'd171478: dataIn1 = 32'd7661
; 
32'd171479: dataIn1 = 32'd6254
; 
32'd171480: dataIn1 = 32'd6260
; 
32'd171481: dataIn1 = 32'd7627
; 
32'd171482: dataIn1 = 32'd7642
; 
32'd171483: dataIn1 = 32'd7658
; 
32'd171484: dataIn1 = 32'd7659
; 
32'd171485: dataIn1 = 32'd7660
; 
32'd171486: dataIn1 = 32'd6254
; 
32'd171487: dataIn1 = 32'd6264
; 
32'd171488: dataIn1 = 32'd7629
; 
32'd171489: dataIn1 = 32'd7658
; 
32'd171490: dataIn1 = 32'd7659
; 
32'd171491: dataIn1 = 32'd7660
; 
32'd171492: dataIn1 = 32'd7662
; 
32'd171493: dataIn1 = 32'd5174
; 
32'd171494: dataIn1 = 32'd6264
; 
32'd171495: dataIn1 = 32'd7640
; 
32'd171496: dataIn1 = 32'd7658
; 
32'd171497: dataIn1 = 32'd7661
; 
32'd171498: dataIn1 = 32'd7815
; 
32'd171499: dataIn1 = 32'd7831
; 
32'd171500: dataIn1 = 32'd2711
; 
32'd171501: dataIn1 = 32'd6264
; 
32'd171502: dataIn1 = 32'd7629
; 
32'd171503: dataIn1 = 32'd7660
; 
32'd171504: dataIn1 = 32'd7662
; 
32'd171505: dataIn1 = 32'd7794
; 
32'd171506: dataIn1 = 32'd7833
; 
32'd171507: dataIn1 = 32'd6252
; 
32'd171508: dataIn1 = 32'd6266
; 
32'd171509: dataIn1 = 32'd7620
; 
32'd171510: dataIn1 = 32'd7663
; 
32'd171511: dataIn1 = 32'd7664
; 
32'd171512: dataIn1 = 32'd7665
; 
32'd171513: dataIn1 = 32'd7666
; 
32'd171514: dataIn1 = 32'd6265
; 
32'd171515: dataIn1 = 32'd6266
; 
32'd171516: dataIn1 = 32'd7663
; 
32'd171517: dataIn1 = 32'd7664
; 
32'd171518: dataIn1 = 32'd7665
; 
32'd171519: dataIn1 = 32'd7667
; 
32'd171520: dataIn1 = 32'd7668
; 
32'd171521: dataIn1 = 32'd6252
; 
32'd171522: dataIn1 = 32'd6265
; 
32'd171523: dataIn1 = 32'd7622
; 
32'd171524: dataIn1 = 32'd7663
; 
32'd171525: dataIn1 = 32'd7664
; 
32'd171526: dataIn1 = 32'd7665
; 
32'd171527: dataIn1 = 32'd7669
; 
32'd171528: dataIn1 = 32'd2709
; 
32'd171529: dataIn1 = 32'd6266
; 
32'd171530: dataIn1 = 32'd7620
; 
32'd171531: dataIn1 = 32'd7663
; 
32'd171532: dataIn1 = 32'd7666
; 
32'd171533: dataIn1 = 32'd7683
; 
32'd171534: dataIn1 = 32'd7757
; 
32'd171535: dataIn1 = 32'd5177
; 
32'd171536: dataIn1 = 32'd6266
; 
32'd171537: dataIn1 = 32'd7664
; 
32'd171538: dataIn1 = 32'd7667
; 
32'd171539: dataIn1 = 32'd7668
; 
32'd171540: dataIn1 = 32'd7754
; 
32'd171541: dataIn1 = 32'd7758
; 
32'd171542: dataIn1 = 32'd5177
; 
32'd171543: dataIn1 = 32'd6265
; 
32'd171544: dataIn1 = 32'd6759
; 
32'd171545: dataIn1 = 32'd7664
; 
32'd171546: dataIn1 = 32'd7667
; 
32'd171547: dataIn1 = 32'd7668
; 
32'd171548: dataIn1 = 32'd5171
; 
32'd171549: dataIn1 = 32'd6265
; 
32'd171550: dataIn1 = 32'd6758
; 
32'd171551: dataIn1 = 32'd7622
; 
32'd171552: dataIn1 = 32'd7665
; 
32'd171553: dataIn1 = 32'd7669
; 
32'd171554: dataIn1 = 32'd6268
; 
32'd171555: dataIn1 = 32'd6269
; 
32'd171556: dataIn1 = 32'd7670
; 
32'd171557: dataIn1 = 32'd7671
; 
32'd171558: dataIn1 = 32'd7672
; 
32'd171559: dataIn1 = 32'd7673
; 
32'd171560: dataIn1 = 32'd7674
; 
32'd171561: dataIn1 = 32'd6267
; 
32'd171562: dataIn1 = 32'd6269
; 
32'd171563: dataIn1 = 32'd7670
; 
32'd171564: dataIn1 = 32'd7671
; 
32'd171565: dataIn1 = 32'd7672
; 
32'd171566: dataIn1 = 32'd7675
; 
32'd171567: dataIn1 = 32'd7676
; 
32'd171568: dataIn1 = 32'd6267
; 
32'd171569: dataIn1 = 32'd6268
; 
32'd171570: dataIn1 = 32'd7670
; 
32'd171571: dataIn1 = 32'd7671
; 
32'd171572: dataIn1 = 32'd7672
; 
32'd171573: dataIn1 = 32'd7677
; 
32'd171574: dataIn1 = 32'd7678
; 
32'd171575: dataIn1 = 32'd5178
; 
32'd171576: dataIn1 = 32'd6269
; 
32'd171577: dataIn1 = 32'd7670
; 
32'd171578: dataIn1 = 32'd7673
; 
32'd171579: dataIn1 = 32'd7674
; 
32'd171580: dataIn1 = 32'd7693
; 
32'd171581: dataIn1 = 32'd7696
; 
32'd171582: dataIn1 = 32'd5178
; 
32'd171583: dataIn1 = 32'd6268
; 
32'd171584: dataIn1 = 32'd7670
; 
32'd171585: dataIn1 = 32'd7673
; 
32'd171586: dataIn1 = 32'd7674
; 
32'd171587: dataIn1 = 32'd7686
; 
32'd171588: dataIn1 = 32'd7689
; 
32'd171589: dataIn1 = 32'd5179
; 
32'd171590: dataIn1 = 32'd6269
; 
32'd171591: dataIn1 = 32'd7671
; 
32'd171592: dataIn1 = 32'd7675
; 
32'd171593: dataIn1 = 32'd7676
; 
32'd171594: dataIn1 = 32'd7694
; 
32'd171595: dataIn1 = 32'd7697
; 
32'd171596: dataIn1 = 32'd5179
; 
32'd171597: dataIn1 = 32'd6267
; 
32'd171598: dataIn1 = 32'd7671
; 
32'd171599: dataIn1 = 32'd7675
; 
32'd171600: dataIn1 = 32'd7676
; 
32'd171601: dataIn1 = 32'd7680
; 
32'd171602: dataIn1 = 32'd7684
; 
32'd171603: dataIn1 = 32'd5180
; 
32'd171604: dataIn1 = 32'd6268
; 
32'd171605: dataIn1 = 32'd7672
; 
32'd171606: dataIn1 = 32'd7677
; 
32'd171607: dataIn1 = 32'd7678
; 
32'd171608: dataIn1 = 32'd7688
; 
32'd171609: dataIn1 = 32'd7692
; 
32'd171610: dataIn1 = 32'd5180
; 
32'd171611: dataIn1 = 32'd6267
; 
32'd171612: dataIn1 = 32'd7672
; 
32'd171613: dataIn1 = 32'd7677
; 
32'd171614: dataIn1 = 32'd7678
; 
32'd171615: dataIn1 = 32'd7681
; 
32'd171616: dataIn1 = 32'd7685
; 
32'd171617: dataIn1 = 32'd6270
; 
32'd171618: dataIn1 = 32'd6271
; 
32'd171619: dataIn1 = 32'd7679
; 
32'd171620: dataIn1 = 32'd7680
; 
32'd171621: dataIn1 = 32'd7681
; 
32'd171622: dataIn1 = 32'd7682
; 
32'd171623: dataIn1 = 32'd7683
; 
32'd171624: dataIn1 = 32'd6267
; 
32'd171625: dataIn1 = 32'd6271
; 
32'd171626: dataIn1 = 32'd7676
; 
32'd171627: dataIn1 = 32'd7679
; 
32'd171628: dataIn1 = 32'd7680
; 
32'd171629: dataIn1 = 32'd7681
; 
32'd171630: dataIn1 = 32'd7684
; 
32'd171631: dataIn1 = 32'd6267
; 
32'd171632: dataIn1 = 32'd6270
; 
32'd171633: dataIn1 = 32'd7678
; 
32'd171634: dataIn1 = 32'd7679
; 
32'd171635: dataIn1 = 32'd7680
; 
32'd171636: dataIn1 = 32'd7681
; 
32'd171637: dataIn1 = 32'd7685
; 
32'd171638: dataIn1 = 32'd2709
; 
32'd171639: dataIn1 = 32'd6271
; 
32'd171640: dataIn1 = 32'd7649
; 
32'd171641: dataIn1 = 32'd7679
; 
32'd171642: dataIn1 = 32'd7682
; 
32'd171643: dataIn1 = 32'd7683
; 
32'd171644: dataIn1 = 32'd7735
; 
32'd171645: dataIn1 = 32'd2709
; 
32'd171646: dataIn1 = 32'd6270
; 
32'd171647: dataIn1 = 32'd7666
; 
32'd171648: dataIn1 = 32'd7679
; 
32'd171649: dataIn1 = 32'd7682
; 
32'd171650: dataIn1 = 32'd7683
; 
32'd171651: dataIn1 = 32'd7757
; 
32'd171652: dataIn1 = 32'd5179
; 
32'd171653: dataIn1 = 32'd6271
; 
32'd171654: dataIn1 = 32'd7676
; 
32'd171655: dataIn1 = 32'd7680
; 
32'd171656: dataIn1 = 32'd7684
; 
32'd171657: dataIn1 = 32'd7732
; 
32'd171658: dataIn1 = 32'd7736
; 
32'd171659: dataIn1 = 32'd5180
; 
32'd171660: dataIn1 = 32'd6270
; 
32'd171661: dataIn1 = 32'd7678
; 
32'd171662: dataIn1 = 32'd7681
; 
32'd171663: dataIn1 = 32'd7685
; 
32'd171664: dataIn1 = 32'd7756
; 
32'd171665: dataIn1 = 32'd7759
; 
32'd171666: dataIn1 = 32'd6268
; 
32'd171667: dataIn1 = 32'd6273
; 
32'd171668: dataIn1 = 32'd7674
; 
32'd171669: dataIn1 = 32'd7686
; 
32'd171670: dataIn1 = 32'd7687
; 
32'd171671: dataIn1 = 32'd7688
; 
32'd171672: dataIn1 = 32'd7689
; 
32'd171673: dataIn1 = 32'd6272
; 
32'd171674: dataIn1 = 32'd6273
; 
32'd171675: dataIn1 = 32'd7686
; 
32'd171676: dataIn1 = 32'd7687
; 
32'd171677: dataIn1 = 32'd7688
; 
32'd171678: dataIn1 = 32'd7690
; 
32'd171679: dataIn1 = 32'd7691
; 
32'd171680: dataIn1 = 32'd6268
; 
32'd171681: dataIn1 = 32'd6272
; 
32'd171682: dataIn1 = 32'd7677
; 
32'd171683: dataIn1 = 32'd7686
; 
32'd171684: dataIn1 = 32'd7687
; 
32'd171685: dataIn1 = 32'd7688
; 
32'd171686: dataIn1 = 32'd7692
; 
32'd171687: dataIn1 = 32'd5178
; 
32'd171688: dataIn1 = 32'd6273
; 
32'd171689: dataIn1 = 32'd7674
; 
32'd171690: dataIn1 = 32'd7686
; 
32'd171691: dataIn1 = 32'd7689
; 
32'd171692: dataIn1 = 32'd7704
; 
32'd171693: dataIn1 = 32'd7716
; 
32'd171694: dataIn1 = 32'd2712
; 
32'd171695: dataIn1 = 32'd6273
; 
32'd171696: dataIn1 = 32'd7687
; 
32'd171697: dataIn1 = 32'd7690
; 
32'd171698: dataIn1 = 32'd7691
; 
32'd171699: dataIn1 = 32'd7717
; 
32'd171700: dataIn1 = 32'd7719
; 
32'd171701: dataIn1 = 32'd2712
; 
32'd171702: dataIn1 = 32'd6272
; 
32'd171703: dataIn1 = 32'd7687
; 
32'd171704: dataIn1 = 32'd7690
; 
32'd171705: dataIn1 = 32'd7691
; 
32'd171706: dataIn1 = 32'd7761
; 
32'd171707: dataIn1 = 32'd7764
; 
32'd171708: dataIn1 = 32'd5180
; 
32'd171709: dataIn1 = 32'd6272
; 
32'd171710: dataIn1 = 32'd7677
; 
32'd171711: dataIn1 = 32'd7688
; 
32'd171712: dataIn1 = 32'd7692
; 
32'd171713: dataIn1 = 32'd7755
; 
32'd171714: dataIn1 = 32'd7762
; 
32'd171715: dataIn1 = 32'd6269
; 
32'd171716: dataIn1 = 32'd6275
; 
32'd171717: dataIn1 = 32'd7673
; 
32'd171718: dataIn1 = 32'd7693
; 
32'd171719: dataIn1 = 32'd7694
; 
32'd171720: dataIn1 = 32'd7695
; 
32'd171721: dataIn1 = 32'd7696
; 
32'd171722: dataIn1 = 32'd6269
; 
32'd171723: dataIn1 = 32'd6274
; 
32'd171724: dataIn1 = 32'd7675
; 
32'd171725: dataIn1 = 32'd7693
; 
32'd171726: dataIn1 = 32'd7694
; 
32'd171727: dataIn1 = 32'd7695
; 
32'd171728: dataIn1 = 32'd7697
; 
32'd171729: dataIn1 = 32'd6274
; 
32'd171730: dataIn1 = 32'd6275
; 
32'd171731: dataIn1 = 32'd7693
; 
32'd171732: dataIn1 = 32'd7694
; 
32'd171733: dataIn1 = 32'd7695
; 
32'd171734: dataIn1 = 32'd7698
; 
32'd171735: dataIn1 = 32'd7699
; 
32'd171736: dataIn1 = 32'd5178
; 
32'd171737: dataIn1 = 32'd6275
; 
32'd171738: dataIn1 = 32'd7673
; 
32'd171739: dataIn1 = 32'd7693
; 
32'd171740: dataIn1 = 32'd7696
; 
32'd171741: dataIn1 = 32'd7703
; 
32'd171742: dataIn1 = 32'd7721
; 
32'd171743: dataIn1 = 32'd5179
; 
32'd171744: dataIn1 = 32'd6274
; 
32'd171745: dataIn1 = 32'd7675
; 
32'd171746: dataIn1 = 32'd7694
; 
32'd171747: dataIn1 = 32'd7697
; 
32'd171748: dataIn1 = 32'd7731
; 
32'd171749: dataIn1 = 32'd7744
; 
32'd171750: dataIn1 = 32'd1109
; 
32'd171751: dataIn1 = 32'd6275
; 
32'd171752: dataIn1 = 32'd7695
; 
32'd171753: dataIn1 = 32'd7698
; 
32'd171754: dataIn1 = 32'd7699
; 
32'd171755: dataIn1 = 32'd7723
; 
32'd171756: dataIn1 = 32'd7725
; 
32'd171757: dataIn1 = 32'd1109
; 
32'd171758: dataIn1 = 32'd6274
; 
32'd171759: dataIn1 = 32'd7695
; 
32'd171760: dataIn1 = 32'd7698
; 
32'd171761: dataIn1 = 32'd7699
; 
32'd171762: dataIn1 = 32'd7745
; 
32'd171763: dataIn1 = 32'd7747
; 
32'd171764: dataIn1 = 32'd6277
; 
32'd171765: dataIn1 = 32'd6278
; 
32'd171766: dataIn1 = 32'd7700
; 
32'd171767: dataIn1 = 32'd7701
; 
32'd171768: dataIn1 = 32'd7702
; 
32'd171769: dataIn1 = 32'd7703
; 
32'd171770: dataIn1 = 32'd7704
; 
32'd171771: dataIn1 = 32'd6276
; 
32'd171772: dataIn1 = 32'd6278
; 
32'd171773: dataIn1 = 32'd7700
; 
32'd171774: dataIn1 = 32'd7701
; 
32'd171775: dataIn1 = 32'd7702
; 
32'd171776: dataIn1 = 32'd7705
; 
32'd171777: dataIn1 = 32'd7706
; 
32'd171778: dataIn1 = 32'd6276
; 
32'd171779: dataIn1 = 32'd6277
; 
32'd171780: dataIn1 = 32'd7700
; 
32'd171781: dataIn1 = 32'd7701
; 
32'd171782: dataIn1 = 32'd7702
; 
32'd171783: dataIn1 = 32'd7707
; 
32'd171784: dataIn1 = 32'd7708
; 
32'd171785: dataIn1 = 32'd5178
; 
32'd171786: dataIn1 = 32'd6278
; 
32'd171787: dataIn1 = 32'd7696
; 
32'd171788: dataIn1 = 32'd7700
; 
32'd171789: dataIn1 = 32'd7703
; 
32'd171790: dataIn1 = 32'd7704
; 
32'd171791: dataIn1 = 32'd7721
; 
32'd171792: dataIn1 = 32'd5178
; 
32'd171793: dataIn1 = 32'd6277
; 
32'd171794: dataIn1 = 32'd7689
; 
32'd171795: dataIn1 = 32'd7700
; 
32'd171796: dataIn1 = 32'd7703
; 
32'd171797: dataIn1 = 32'd7704
; 
32'd171798: dataIn1 = 32'd7716
; 
32'd171799: dataIn1 = 32'd2646
; 
32'd171800: dataIn1 = 32'd6278
; 
32'd171801: dataIn1 = 32'd7701
; 
32'd171802: dataIn1 = 32'd7705
; 
32'd171803: dataIn1 = 32'd7706
; 
32'd171804: dataIn1 = 32'd7722
; 
32'd171805: dataIn1 = 32'd7724
; 
32'd171806: dataIn1 = 32'd2646
; 
32'd171807: dataIn1 = 32'd6276
; 
32'd171808: dataIn1 = 32'd7701
; 
32'd171809: dataIn1 = 32'd7705
; 
32'd171810: dataIn1 = 32'd7706
; 
32'd171811: dataIn1 = 32'd7710
; 
32'd171812: dataIn1 = 32'd7714
; 
32'd171813: dataIn1 = 32'd5181
; 
32'd171814: dataIn1 = 32'd6277
; 
32'd171815: dataIn1 = 32'd7702
; 
32'd171816: dataIn1 = 32'd7707
; 
32'd171817: dataIn1 = 32'd7708
; 
32'd171818: dataIn1 = 32'd7718
; 
32'd171819: dataIn1 = 32'd7720
; 
32'd171820: dataIn1 = 32'd5181
; 
32'd171821: dataIn1 = 32'd6276
; 
32'd171822: dataIn1 = 32'd7702
; 
32'd171823: dataIn1 = 32'd7707
; 
32'd171824: dataIn1 = 32'd7708
; 
32'd171825: dataIn1 = 32'd7711
; 
32'd171826: dataIn1 = 32'd7715
; 
32'd171827: dataIn1 = 32'd4939
; 
32'd171828: dataIn1 = 32'd6279
; 
32'd171829: dataIn1 = 32'd7709
; 
32'd171830: dataIn1 = 32'd7710
; 
32'd171831: dataIn1 = 32'd7711
; 
32'd171832: dataIn1 = 32'd7712
; 
32'd171833: dataIn1 = 32'd7713
; 
32'd171834: dataIn1 = 32'd4939
; 
32'd171835: dataIn1 = 32'd6276
; 
32'd171836: dataIn1 = 32'd7706
; 
32'd171837: dataIn1 = 32'd7709
; 
32'd171838: dataIn1 = 32'd7710
; 
32'd171839: dataIn1 = 32'd7711
; 
32'd171840: dataIn1 = 32'd7714
; 
32'd171841: dataIn1 = 32'd6276
; 
32'd171842: dataIn1 = 32'd6279
; 
32'd171843: dataIn1 = 32'd7708
; 
32'd171844: dataIn1 = 32'd7709
; 
32'd171845: dataIn1 = 32'd7710
; 
32'd171846: dataIn1 = 32'd7711
; 
32'd171847: dataIn1 = 32'd7715
; 
32'd171848: dataIn1 = 32'd7
; 
32'd171849: dataIn1 = 32'd4939
; 
32'd171850: dataIn1 = 32'd7709
; 
32'd171851: dataIn1 = 32'd7712
; 
32'd171852: dataIn1 = 32'd7713
; 
32'd171853: dataIn1 = 32'd9605
; 
32'd171854: dataIn1 = 32'd9660
; 
32'd171855: dataIn1 = 32'd7
; 
32'd171856: dataIn1 = 32'd6279
; 
32'd171857: dataIn1 = 32'd7605
; 
32'd171858: dataIn1 = 32'd7709
; 
32'd171859: dataIn1 = 32'd7712
; 
32'd171860: dataIn1 = 32'd7713
; 
32'd171861: dataIn1 = 32'd9008
; 
32'd171862: dataIn1 = 32'd2646
; 
32'd171863: dataIn1 = 32'd4939
; 
32'd171864: dataIn1 = 32'd7706
; 
32'd171865: dataIn1 = 32'd7710
; 
32'd171866: dataIn1 = 32'd7714
; 
32'd171867: dataIn1 = 32'd9658
; 
32'd171868: dataIn1 = 32'd9659
; 
32'd171869: dataIn1 = 32'd5181
; 
32'd171870: dataIn1 = 32'd6279
; 
32'd171871: dataIn1 = 32'd7708
; 
32'd171872: dataIn1 = 32'd7711
; 
32'd171873: dataIn1 = 32'd7715
; 
32'd171874: dataIn1 = 32'd9005
; 
32'd171875: dataIn1 = 32'd9009
; 
32'd171876: dataIn1 = 32'd6273
; 
32'd171877: dataIn1 = 32'd6277
; 
32'd171878: dataIn1 = 32'd7689
; 
32'd171879: dataIn1 = 32'd7704
; 
32'd171880: dataIn1 = 32'd7716
; 
32'd171881: dataIn1 = 32'd7717
; 
32'd171882: dataIn1 = 32'd7718
; 
32'd171883: dataIn1 = 32'd6273
; 
32'd171884: dataIn1 = 32'd6280
; 
32'd171885: dataIn1 = 32'd7690
; 
32'd171886: dataIn1 = 32'd7716
; 
32'd171887: dataIn1 = 32'd7717
; 
32'd171888: dataIn1 = 32'd7718
; 
32'd171889: dataIn1 = 32'd7719
; 
32'd171890: dataIn1 = 32'd6277
; 
32'd171891: dataIn1 = 32'd6280
; 
32'd171892: dataIn1 = 32'd7707
; 
32'd171893: dataIn1 = 32'd7716
; 
32'd171894: dataIn1 = 32'd7717
; 
32'd171895: dataIn1 = 32'd7718
; 
32'd171896: dataIn1 = 32'd7720
; 
32'd171897: dataIn1 = 32'd2712
; 
32'd171898: dataIn1 = 32'd6280
; 
32'd171899: dataIn1 = 32'd7690
; 
32'd171900: dataIn1 = 32'd7717
; 
32'd171901: dataIn1 = 32'd7719
; 
32'd171902: dataIn1 = 32'd8997
; 
32'd171903: dataIn1 = 32'd9016
; 
32'd171904: dataIn1 = 32'd5181
; 
32'd171905: dataIn1 = 32'd6280
; 
32'd171906: dataIn1 = 32'd7707
; 
32'd171907: dataIn1 = 32'd7718
; 
32'd171908: dataIn1 = 32'd7720
; 
32'd171909: dataIn1 = 32'd9004
; 
32'd171910: dataIn1 = 32'd9015
; 
32'd171911: dataIn1 = 32'd6275
; 
32'd171912: dataIn1 = 32'd6278
; 
32'd171913: dataIn1 = 32'd7696
; 
32'd171914: dataIn1 = 32'd7703
; 
32'd171915: dataIn1 = 32'd7721
; 
32'd171916: dataIn1 = 32'd7722
; 
32'd171917: dataIn1 = 32'd7723
; 
32'd171918: dataIn1 = 32'd4940
; 
32'd171919: dataIn1 = 32'd6278
; 
32'd171920: dataIn1 = 32'd7705
; 
32'd171921: dataIn1 = 32'd7721
; 
32'd171922: dataIn1 = 32'd7722
; 
32'd171923: dataIn1 = 32'd7723
; 
32'd171924: dataIn1 = 32'd7724
; 
32'd171925: dataIn1 = 32'd4940
; 
32'd171926: dataIn1 = 32'd6275
; 
32'd171927: dataIn1 = 32'd7698
; 
32'd171928: dataIn1 = 32'd7721
; 
32'd171929: dataIn1 = 32'd7722
; 
32'd171930: dataIn1 = 32'd7723
; 
32'd171931: dataIn1 = 32'd7725
; 
32'd171932: dataIn1 = 32'd2646
; 
32'd171933: dataIn1 = 32'd4940
; 
32'd171934: dataIn1 = 32'd7705
; 
32'd171935: dataIn1 = 32'd7722
; 
32'd171936: dataIn1 = 32'd7724
; 
32'd171937: dataIn1 = 32'd9657
; 
32'd171938: dataIn1 = 32'd9662
; 
32'd171939: dataIn1 = 32'd1109
; 
32'd171940: dataIn1 = 32'd4940
; 
32'd171941: dataIn1 = 32'd7698
; 
32'd171942: dataIn1 = 32'd7723
; 
32'd171943: dataIn1 = 32'd7725
; 
32'd171944: dataIn1 = 32'd9645
; 
32'd171945: dataIn1 = 32'd9664
; 
32'd171946: dataIn1 = 32'd6282
; 
32'd171947: dataIn1 = 32'd6283
; 
32'd171948: dataIn1 = 32'd7726
; 
32'd171949: dataIn1 = 32'd7727
; 
32'd171950: dataIn1 = 32'd7728
; 
32'd171951: dataIn1 = 32'd7729
; 
32'd171952: dataIn1 = 32'd7730
; 
32'd171953: dataIn1 = 32'd6281
; 
32'd171954: dataIn1 = 32'd6283
; 
32'd171955: dataIn1 = 32'd7726
; 
32'd171956: dataIn1 = 32'd7727
; 
32'd171957: dataIn1 = 32'd7728
; 
32'd171958: dataIn1 = 32'd7731
; 
32'd171959: dataIn1 = 32'd7732
; 
32'd171960: dataIn1 = 32'd6281
; 
32'd171961: dataIn1 = 32'd6282
; 
32'd171962: dataIn1 = 32'd7726
; 
32'd171963: dataIn1 = 32'd7727
; 
32'd171964: dataIn1 = 32'd7728
; 
32'd171965: dataIn1 = 32'd7733
; 
32'd171966: dataIn1 = 32'd7734
; 
32'd171967: dataIn1 = 32'd2645
; 
32'd171968: dataIn1 = 32'd6283
; 
32'd171969: dataIn1 = 32'd7726
; 
32'd171970: dataIn1 = 32'd7729
; 
32'd171971: dataIn1 = 32'd7730
; 
32'd171972: dataIn1 = 32'd7743
; 
32'd171973: dataIn1 = 32'd7746
; 
32'd171974: dataIn1 = 32'd2645
; 
32'd171975: dataIn1 = 32'd6282
; 
32'd171976: dataIn1 = 32'd7726
; 
32'd171977: dataIn1 = 32'd7729
; 
32'd171978: dataIn1 = 32'd7730
; 
32'd171979: dataIn1 = 32'd7738
; 
32'd171980: dataIn1 = 32'd7741
; 
32'd171981: dataIn1 = 32'd5179
; 
32'd171982: dataIn1 = 32'd6283
; 
32'd171983: dataIn1 = 32'd7697
; 
32'd171984: dataIn1 = 32'd7727
; 
32'd171985: dataIn1 = 32'd7731
; 
32'd171986: dataIn1 = 32'd7732
; 
32'd171987: dataIn1 = 32'd7744
; 
32'd171988: dataIn1 = 32'd5179
; 
32'd171989: dataIn1 = 32'd6281
; 
32'd171990: dataIn1 = 32'd7684
; 
32'd171991: dataIn1 = 32'd7727
; 
32'd171992: dataIn1 = 32'd7731
; 
32'd171993: dataIn1 = 32'd7732
; 
32'd171994: dataIn1 = 32'd7736
; 
32'd171995: dataIn1 = 32'd5175
; 
32'd171996: dataIn1 = 32'd6282
; 
32'd171997: dataIn1 = 32'd7657
; 
32'd171998: dataIn1 = 32'd7728
; 
32'd171999: dataIn1 = 32'd7733
; 
32'd172000: dataIn1 = 32'd7734
; 
32'd172001: dataIn1 = 32'd7740
; 
32'd172002: dataIn1 = 32'd5175
; 
32'd172003: dataIn1 = 32'd6281
; 
32'd172004: dataIn1 = 32'd7650
; 
32'd172005: dataIn1 = 32'd7728
; 
32'd172006: dataIn1 = 32'd7733
; 
32'd172007: dataIn1 = 32'd7734
; 
32'd172008: dataIn1 = 32'd7737
; 
32'd172009: dataIn1 = 32'd6261
; 
32'd172010: dataIn1 = 32'd6271
; 
32'd172011: dataIn1 = 32'd7649
; 
32'd172012: dataIn1 = 32'd7682
; 
32'd172013: dataIn1 = 32'd7735
; 
32'd172014: dataIn1 = 32'd7736
; 
32'd172015: dataIn1 = 32'd7737
; 
32'd172016: dataIn1 = 32'd6271
; 
32'd172017: dataIn1 = 32'd6281
; 
32'd172018: dataIn1 = 32'd7684
; 
32'd172019: dataIn1 = 32'd7732
; 
32'd172020: dataIn1 = 32'd7735
; 
32'd172021: dataIn1 = 32'd7736
; 
32'd172022: dataIn1 = 32'd7737
; 
32'd172023: dataIn1 = 32'd6261
; 
32'd172024: dataIn1 = 32'd6281
; 
32'd172025: dataIn1 = 32'd7650
; 
32'd172026: dataIn1 = 32'd7734
; 
32'd172027: dataIn1 = 32'd7735
; 
32'd172028: dataIn1 = 32'd7736
; 
32'd172029: dataIn1 = 32'd7737
; 
32'd172030: dataIn1 = 32'd4934
; 
32'd172031: dataIn1 = 32'd6282
; 
32'd172032: dataIn1 = 32'd7730
; 
32'd172033: dataIn1 = 32'd7738
; 
32'd172034: dataIn1 = 32'd7739
; 
32'd172035: dataIn1 = 32'd7740
; 
32'd172036: dataIn1 = 32'd7741
; 
32'd172037: dataIn1 = 32'd4934
; 
32'd172038: dataIn1 = 32'd6262
; 
32'd172039: dataIn1 = 32'd7656
; 
32'd172040: dataIn1 = 32'd7738
; 
32'd172041: dataIn1 = 32'd7739
; 
32'd172042: dataIn1 = 32'd7740
; 
32'd172043: dataIn1 = 32'd7742
; 
32'd172044: dataIn1 = 32'd6262
; 
32'd172045: dataIn1 = 32'd6282
; 
32'd172046: dataIn1 = 32'd7657
; 
32'd172047: dataIn1 = 32'd7733
; 
32'd172048: dataIn1 = 32'd7738
; 
32'd172049: dataIn1 = 32'd7739
; 
32'd172050: dataIn1 = 32'd7740
; 
32'd172051: dataIn1 = 32'd2645
; 
32'd172052: dataIn1 = 32'd4934
; 
32'd172053: dataIn1 = 32'd7730
; 
32'd172054: dataIn1 = 32'd7738
; 
32'd172055: dataIn1 = 32'd7741
; 
32'd172056: dataIn1 = 32'd9649
; 
32'd172057: dataIn1 = 32'd9651
; 
32'd172058: dataIn1 = 32'd136
; 
32'd172059: dataIn1 = 32'd4934
; 
32'd172060: dataIn1 = 32'd7656
; 
32'd172061: dataIn1 = 32'd7739
; 
32'd172062: dataIn1 = 32'd7742
; 
32'd172063: dataIn1 = 32'd9610
; 
32'd172064: dataIn1 = 32'd9650
; 
32'd172065: dataIn1 = 32'd4935
; 
32'd172066: dataIn1 = 32'd6283
; 
32'd172067: dataIn1 = 32'd7729
; 
32'd172068: dataIn1 = 32'd7743
; 
32'd172069: dataIn1 = 32'd7744
; 
32'd172070: dataIn1 = 32'd7745
; 
32'd172071: dataIn1 = 32'd7746
; 
32'd172072: dataIn1 = 32'd6274
; 
32'd172073: dataIn1 = 32'd6283
; 
32'd172074: dataIn1 = 32'd7697
; 
32'd172075: dataIn1 = 32'd7731
; 
32'd172076: dataIn1 = 32'd7743
; 
32'd172077: dataIn1 = 32'd7744
; 
32'd172078: dataIn1 = 32'd7745
; 
32'd172079: dataIn1 = 32'd4935
; 
32'd172080: dataIn1 = 32'd6274
; 
32'd172081: dataIn1 = 32'd7699
; 
32'd172082: dataIn1 = 32'd7743
; 
32'd172083: dataIn1 = 32'd7744
; 
32'd172084: dataIn1 = 32'd7745
; 
32'd172085: dataIn1 = 32'd7747
; 
32'd172086: dataIn1 = 32'd2645
; 
32'd172087: dataIn1 = 32'd4935
; 
32'd172088: dataIn1 = 32'd7729
; 
32'd172089: dataIn1 = 32'd7743
; 
32'd172090: dataIn1 = 32'd7746
; 
32'd172091: dataIn1 = 32'd9647
; 
32'd172092: dataIn1 = 32'd9654
; 
32'd172093: dataIn1 = 32'd1109
; 
32'd172094: dataIn1 = 32'd4935
; 
32'd172095: dataIn1 = 32'd7699
; 
32'd172096: dataIn1 = 32'd7745
; 
32'd172097: dataIn1 = 32'd7747
; 
32'd172098: dataIn1 = 32'd9644
; 
32'd172099: dataIn1 = 32'd9655
; 
32'd172100: dataIn1 = 32'd6285
; 
32'd172101: dataIn1 = 32'd6286
; 
32'd172102: dataIn1 = 32'd7748
; 
32'd172103: dataIn1 = 32'd7749
; 
32'd172104: dataIn1 = 32'd7750
; 
32'd172105: dataIn1 = 32'd7751
; 
32'd172106: dataIn1 = 32'd7752
; 
32'd172107: dataIn1 = 32'd6284
; 
32'd172108: dataIn1 = 32'd6286
; 
32'd172109: dataIn1 = 32'd7748
; 
32'd172110: dataIn1 = 32'd7749
; 
32'd172111: dataIn1 = 32'd7750
; 
32'd172112: dataIn1 = 32'd7753
; 
32'd172113: dataIn1 = 32'd7754
; 
32'd172114: dataIn1 = 32'd6284
; 
32'd172115: dataIn1 = 32'd6285
; 
32'd172116: dataIn1 = 32'd7748
; 
32'd172117: dataIn1 = 32'd7749
; 
32'd172118: dataIn1 = 32'd7750
; 
32'd172119: dataIn1 = 32'd7755
; 
32'd172120: dataIn1 = 32'd7756
; 
32'd172121: dataIn1 = 32'd5182
; 
32'd172122: dataIn1 = 32'd6286
; 
32'd172123: dataIn1 = 32'd6761
; 
32'd172124: dataIn1 = 32'd7748
; 
32'd172125: dataIn1 = 32'd7751
; 
32'd172126: dataIn1 = 32'd7752
; 
32'd172127: dataIn1 = 32'd5182
; 
32'd172128: dataIn1 = 32'd6285
; 
32'd172129: dataIn1 = 32'd7748
; 
32'd172130: dataIn1 = 32'd7751
; 
32'd172131: dataIn1 = 32'd7752
; 
32'd172132: dataIn1 = 32'd7760
; 
32'd172133: dataIn1 = 32'd7763
; 
32'd172134: dataIn1 = 32'd5177
; 
32'd172135: dataIn1 = 32'd6286
; 
32'd172136: dataIn1 = 32'd6760
; 
32'd172137: dataIn1 = 32'd7749
; 
32'd172138: dataIn1 = 32'd7753
; 
32'd172139: dataIn1 = 32'd7754
; 
32'd172140: dataIn1 = 32'd5177
; 
32'd172141: dataIn1 = 32'd6284
; 
32'd172142: dataIn1 = 32'd7667
; 
32'd172143: dataIn1 = 32'd7749
; 
32'd172144: dataIn1 = 32'd7753
; 
32'd172145: dataIn1 = 32'd7754
; 
32'd172146: dataIn1 = 32'd7758
; 
32'd172147: dataIn1 = 32'd5180
; 
32'd172148: dataIn1 = 32'd6285
; 
32'd172149: dataIn1 = 32'd7692
; 
32'd172150: dataIn1 = 32'd7750
; 
32'd172151: dataIn1 = 32'd7755
; 
32'd172152: dataIn1 = 32'd7756
; 
32'd172153: dataIn1 = 32'd7762
; 
32'd172154: dataIn1 = 32'd5180
; 
32'd172155: dataIn1 = 32'd6284
; 
32'd172156: dataIn1 = 32'd7685
; 
32'd172157: dataIn1 = 32'd7750
; 
32'd172158: dataIn1 = 32'd7755
; 
32'd172159: dataIn1 = 32'd7756
; 
32'd172160: dataIn1 = 32'd7759
; 
32'd172161: dataIn1 = 32'd6266
; 
32'd172162: dataIn1 = 32'd6270
; 
32'd172163: dataIn1 = 32'd7666
; 
32'd172164: dataIn1 = 32'd7683
; 
32'd172165: dataIn1 = 32'd7757
; 
32'd172166: dataIn1 = 32'd7758
; 
32'd172167: dataIn1 = 32'd7759
; 
32'd172168: dataIn1 = 32'd6266
; 
32'd172169: dataIn1 = 32'd6284
; 
32'd172170: dataIn1 = 32'd7667
; 
32'd172171: dataIn1 = 32'd7754
; 
32'd172172: dataIn1 = 32'd7757
; 
32'd172173: dataIn1 = 32'd7758
; 
32'd172174: dataIn1 = 32'd7759
; 
32'd172175: dataIn1 = 32'd6270
; 
32'd172176: dataIn1 = 32'd6284
; 
32'd172177: dataIn1 = 32'd7685
; 
32'd172178: dataIn1 = 32'd7756
; 
32'd172179: dataIn1 = 32'd7757
; 
32'd172180: dataIn1 = 32'd7758
; 
32'd172181: dataIn1 = 32'd7759
; 
32'd172182: dataIn1 = 32'd6285
; 
32'd172183: dataIn1 = 32'd6287
; 
32'd172184: dataIn1 = 32'd7752
; 
32'd172185: dataIn1 = 32'd7760
; 
32'd172186: dataIn1 = 32'd7761
; 
32'd172187: dataIn1 = 32'd7762
; 
32'd172188: dataIn1 = 32'd7763
; 
32'd172189: dataIn1 = 32'd6272
; 
32'd172190: dataIn1 = 32'd6287
; 
32'd172191: dataIn1 = 32'd7691
; 
32'd172192: dataIn1 = 32'd7760
; 
32'd172193: dataIn1 = 32'd7761
; 
32'd172194: dataIn1 = 32'd7762
; 
32'd172195: dataIn1 = 32'd7764
; 
32'd172196: dataIn1 = 32'd6272
; 
32'd172197: dataIn1 = 32'd6285
; 
32'd172198: dataIn1 = 32'd7692
; 
32'd172199: dataIn1 = 32'd7755
; 
32'd172200: dataIn1 = 32'd7760
; 
32'd172201: dataIn1 = 32'd7761
; 
32'd172202: dataIn1 = 32'd7762
; 
32'd172203: dataIn1 = 32'd5182
; 
32'd172204: dataIn1 = 32'd6287
; 
32'd172205: dataIn1 = 32'd7752
; 
32'd172206: dataIn1 = 32'd7760
; 
32'd172207: dataIn1 = 32'd7763
; 
32'd172208: dataIn1 = 32'd9017
; 
32'd172209: dataIn1 = 32'd9020
; 
32'd172210: dataIn1 = 32'd2712
; 
32'd172211: dataIn1 = 32'd6287
; 
32'd172212: dataIn1 = 32'd7691
; 
32'd172213: dataIn1 = 32'd7761
; 
32'd172214: dataIn1 = 32'd7764
; 
32'd172215: dataIn1 = 32'd8998
; 
32'd172216: dataIn1 = 32'd9019
; 
32'd172217: dataIn1 = 32'd6289
; 
32'd172218: dataIn1 = 32'd6290
; 
32'd172219: dataIn1 = 32'd7765
; 
32'd172220: dataIn1 = 32'd7766
; 
32'd172221: dataIn1 = 32'd7767
; 
32'd172222: dataIn1 = 32'd7768
; 
32'd172223: dataIn1 = 32'd7769
; 
32'd172224: dataIn1 = 32'd6288
; 
32'd172225: dataIn1 = 32'd6290
; 
32'd172226: dataIn1 = 32'd7765
; 
32'd172227: dataIn1 = 32'd7766
; 
32'd172228: dataIn1 = 32'd7767
; 
32'd172229: dataIn1 = 32'd7770
; 
32'd172230: dataIn1 = 32'd7771
; 
32'd172231: dataIn1 = 32'd6288
; 
32'd172232: dataIn1 = 32'd6289
; 
32'd172233: dataIn1 = 32'd7765
; 
32'd172234: dataIn1 = 32'd7766
; 
32'd172235: dataIn1 = 32'd7767
; 
32'd172236: dataIn1 = 32'd7772
; 
32'd172237: dataIn1 = 32'd7773
; 
32'd172238: dataIn1 = 32'd5183
; 
32'd172239: dataIn1 = 32'd6290
; 
32'd172240: dataIn1 = 32'd7765
; 
32'd172241: dataIn1 = 32'd7768
; 
32'd172242: dataIn1 = 32'd7769
; 
32'd172243: dataIn1 = 32'd7788
; 
32'd172244: dataIn1 = 32'd7791
; 
32'd172245: dataIn1 = 32'd5183
; 
32'd172246: dataIn1 = 32'd6289
; 
32'd172247: dataIn1 = 32'd7765
; 
32'd172248: dataIn1 = 32'd7768
; 
32'd172249: dataIn1 = 32'd7769
; 
32'd172250: dataIn1 = 32'd7781
; 
32'd172251: dataIn1 = 32'd7784
; 
32'd172252: dataIn1 = 32'd5184
; 
32'd172253: dataIn1 = 32'd6290
; 
32'd172254: dataIn1 = 32'd7766
; 
32'd172255: dataIn1 = 32'd7770
; 
32'd172256: dataIn1 = 32'd7771
; 
32'd172257: dataIn1 = 32'd7789
; 
32'd172258: dataIn1 = 32'd7792
; 
32'd172259: dataIn1 = 32'd5184
; 
32'd172260: dataIn1 = 32'd6288
; 
32'd172261: dataIn1 = 32'd7766
; 
32'd172262: dataIn1 = 32'd7770
; 
32'd172263: dataIn1 = 32'd7771
; 
32'd172264: dataIn1 = 32'd7775
; 
32'd172265: dataIn1 = 32'd7779
; 
32'd172266: dataIn1 = 32'd5185
; 
32'd172267: dataIn1 = 32'd6289
; 
32'd172268: dataIn1 = 32'd7767
; 
32'd172269: dataIn1 = 32'd7772
; 
32'd172270: dataIn1 = 32'd7773
; 
32'd172271: dataIn1 = 32'd7783
; 
32'd172272: dataIn1 = 32'd7787
; 
32'd172273: dataIn1 = 32'd5185
; 
32'd172274: dataIn1 = 32'd6288
; 
32'd172275: dataIn1 = 32'd7767
; 
32'd172276: dataIn1 = 32'd7772
; 
32'd172277: dataIn1 = 32'd7773
; 
32'd172278: dataIn1 = 32'd7776
; 
32'd172279: dataIn1 = 32'd7780
; 
32'd172280: dataIn1 = 32'd6291
; 
32'd172281: dataIn1 = 32'd6292
; 
32'd172282: dataIn1 = 32'd7774
; 
32'd172283: dataIn1 = 32'd7775
; 
32'd172284: dataIn1 = 32'd7776
; 
32'd172285: dataIn1 = 32'd7777
; 
32'd172286: dataIn1 = 32'd7778
; 
32'd172287: dataIn1 = 32'd6288
; 
32'd172288: dataIn1 = 32'd6292
; 
32'd172289: dataIn1 = 32'd7771
; 
32'd172290: dataIn1 = 32'd7774
; 
32'd172291: dataIn1 = 32'd7775
; 
32'd172292: dataIn1 = 32'd7776
; 
32'd172293: dataIn1 = 32'd7779
; 
32'd172294: dataIn1 = 32'd6288
; 
32'd172295: dataIn1 = 32'd6291
; 
32'd172296: dataIn1 = 32'd7773
; 
32'd172297: dataIn1 = 32'd7774
; 
32'd172298: dataIn1 = 32'd7775
; 
32'd172299: dataIn1 = 32'd7776
; 
32'd172300: dataIn1 = 32'd7780
; 
32'd172301: dataIn1 = 32'd1110
; 
32'd172302: dataIn1 = 32'd6292
; 
32'd172303: dataIn1 = 32'd7774
; 
32'd172304: dataIn1 = 32'd7777
; 
32'd172305: dataIn1 = 32'd7778
; 
32'd172306: dataIn1 = 32'd7821
; 
32'd172307: dataIn1 = 32'd7824
; 
32'd172308: dataIn1 = 32'd1110
; 
32'd172309: dataIn1 = 32'd6291
; 
32'd172310: dataIn1 = 32'd7774
; 
32'd172311: dataIn1 = 32'd7777
; 
32'd172312: dataIn1 = 32'd7778
; 
32'd172313: dataIn1 = 32'd7843
; 
32'd172314: dataIn1 = 32'd7846
; 
32'd172315: dataIn1 = 32'd5184
; 
32'd172316: dataIn1 = 32'd6292
; 
32'd172317: dataIn1 = 32'd7771
; 
32'd172318: dataIn1 = 32'd7775
; 
32'd172319: dataIn1 = 32'd7779
; 
32'd172320: dataIn1 = 32'd7818
; 
32'd172321: dataIn1 = 32'd7822
; 
32'd172322: dataIn1 = 32'd5185
; 
32'd172323: dataIn1 = 32'd6291
; 
32'd172324: dataIn1 = 32'd7773
; 
32'd172325: dataIn1 = 32'd7776
; 
32'd172326: dataIn1 = 32'd7780
; 
32'd172327: dataIn1 = 32'd7842
; 
32'd172328: dataIn1 = 32'd7845
; 
32'd172329: dataIn1 = 32'd6289
; 
32'd172330: dataIn1 = 32'd6294
; 
32'd172331: dataIn1 = 32'd7769
; 
32'd172332: dataIn1 = 32'd7781
; 
32'd172333: dataIn1 = 32'd7782
; 
32'd172334: dataIn1 = 32'd7783
; 
32'd172335: dataIn1 = 32'd7784
; 
32'd172336: dataIn1 = 32'd6293
; 
32'd172337: dataIn1 = 32'd6294
; 
32'd172338: dataIn1 = 32'd7781
; 
32'd172339: dataIn1 = 32'd7782
; 
32'd172340: dataIn1 = 32'd7783
; 
32'd172341: dataIn1 = 32'd7785
; 
32'd172342: dataIn1 = 32'd7786
; 
32'd172343: dataIn1 = 32'd6289
; 
32'd172344: dataIn1 = 32'd6293
; 
32'd172345: dataIn1 = 32'd7772
; 
32'd172346: dataIn1 = 32'd7781
; 
32'd172347: dataIn1 = 32'd7782
; 
32'd172348: dataIn1 = 32'd7783
; 
32'd172349: dataIn1 = 32'd7787
; 
32'd172350: dataIn1 = 32'd5183
; 
32'd172351: dataIn1 = 32'd6294
; 
32'd172352: dataIn1 = 32'd7769
; 
32'd172353: dataIn1 = 32'd7781
; 
32'd172354: dataIn1 = 32'd7784
; 
32'd172355: dataIn1 = 32'd7799
; 
32'd172356: dataIn1 = 32'd7804
; 
32'd172357: dataIn1 = 32'd2713
; 
32'd172358: dataIn1 = 32'd6294
; 
32'd172359: dataIn1 = 32'd7782
; 
32'd172360: dataIn1 = 32'd7785
; 
32'd172361: dataIn1 = 32'd7786
; 
32'd172362: dataIn1 = 32'd7805
; 
32'd172363: dataIn1 = 32'd7807
; 
32'd172364: dataIn1 = 32'd2713
; 
32'd172365: dataIn1 = 32'd6293
; 
32'd172366: dataIn1 = 32'd7782
; 
32'd172367: dataIn1 = 32'd7785
; 
32'd172368: dataIn1 = 32'd7786
; 
32'd172369: dataIn1 = 32'd7849
; 
32'd172370: dataIn1 = 32'd7852
; 
32'd172371: dataIn1 = 32'd5185
; 
32'd172372: dataIn1 = 32'd6293
; 
32'd172373: dataIn1 = 32'd7772
; 
32'd172374: dataIn1 = 32'd7783
; 
32'd172375: dataIn1 = 32'd7787
; 
32'd172376: dataIn1 = 32'd7841
; 
32'd172377: dataIn1 = 32'd7850
; 
32'd172378: dataIn1 = 32'd6290
; 
32'd172379: dataIn1 = 32'd6296
; 
32'd172380: dataIn1 = 32'd7768
; 
32'd172381: dataIn1 = 32'd7788
; 
32'd172382: dataIn1 = 32'd7789
; 
32'd172383: dataIn1 = 32'd7790
; 
32'd172384: dataIn1 = 32'd7791
; 
32'd172385: dataIn1 = 32'd6290
; 
32'd172386: dataIn1 = 32'd6295
; 
32'd172387: dataIn1 = 32'd7770
; 
32'd172388: dataIn1 = 32'd7788
; 
32'd172389: dataIn1 = 32'd7789
; 
32'd172390: dataIn1 = 32'd7790
; 
32'd172391: dataIn1 = 32'd7792
; 
32'd172392: dataIn1 = 32'd6295
; 
32'd172393: dataIn1 = 32'd6296
; 
32'd172394: dataIn1 = 32'd7788
; 
32'd172395: dataIn1 = 32'd7789
; 
32'd172396: dataIn1 = 32'd7790
; 
32'd172397: dataIn1 = 32'd7793
; 
32'd172398: dataIn1 = 32'd7794
; 
32'd172399: dataIn1 = 32'd5183
; 
32'd172400: dataIn1 = 32'd6296
; 
32'd172401: dataIn1 = 32'd7768
; 
32'd172402: dataIn1 = 32'd7788
; 
32'd172403: dataIn1 = 32'd7791
; 
32'd172404: dataIn1 = 32'd7798
; 
32'd172405: dataIn1 = 32'd7809
; 
32'd172406: dataIn1 = 32'd5184
; 
32'd172407: dataIn1 = 32'd6295
; 
32'd172408: dataIn1 = 32'd7770
; 
32'd172409: dataIn1 = 32'd7789
; 
32'd172410: dataIn1 = 32'd7792
; 
32'd172411: dataIn1 = 32'd7817
; 
32'd172412: dataIn1 = 32'd7832
; 
32'd172413: dataIn1 = 32'd2711
; 
32'd172414: dataIn1 = 32'd6296
; 
32'd172415: dataIn1 = 32'd7636
; 
32'd172416: dataIn1 = 32'd7790
; 
32'd172417: dataIn1 = 32'd7793
; 
32'd172418: dataIn1 = 32'd7794
; 
32'd172419: dataIn1 = 32'd7811
; 
32'd172420: dataIn1 = 32'd2711
; 
32'd172421: dataIn1 = 32'd6295
; 
32'd172422: dataIn1 = 32'd7662
; 
32'd172423: dataIn1 = 32'd7790
; 
32'd172424: dataIn1 = 32'd7793
; 
32'd172425: dataIn1 = 32'd7794
; 
32'd172426: dataIn1 = 32'd7833
; 
32'd172427: dataIn1 = 32'd6298
; 
32'd172428: dataIn1 = 32'd6299
; 
32'd172429: dataIn1 = 32'd7795
; 
32'd172430: dataIn1 = 32'd7796
; 
32'd172431: dataIn1 = 32'd7797
; 
32'd172432: dataIn1 = 32'd7798
; 
32'd172433: dataIn1 = 32'd7799
; 
32'd172434: dataIn1 = 32'd6297
; 
32'd172435: dataIn1 = 32'd6299
; 
32'd172436: dataIn1 = 32'd7795
; 
32'd172437: dataIn1 = 32'd7796
; 
32'd172438: dataIn1 = 32'd7797
; 
32'd172439: dataIn1 = 32'd7800
; 
32'd172440: dataIn1 = 32'd7801
; 
32'd172441: dataIn1 = 32'd6297
; 
32'd172442: dataIn1 = 32'd6298
; 
32'd172443: dataIn1 = 32'd7795
; 
32'd172444: dataIn1 = 32'd7796
; 
32'd172445: dataIn1 = 32'd7797
; 
32'd172446: dataIn1 = 32'd7802
; 
32'd172447: dataIn1 = 32'd7803
; 
32'd172448: dataIn1 = 32'd5183
; 
32'd172449: dataIn1 = 32'd6299
; 
32'd172450: dataIn1 = 32'd7791
; 
32'd172451: dataIn1 = 32'd7795
; 
32'd172452: dataIn1 = 32'd7798
; 
32'd172453: dataIn1 = 32'd7799
; 
32'd172454: dataIn1 = 32'd7809
; 
32'd172455: dataIn1 = 32'd5183
; 
32'd172456: dataIn1 = 32'd6298
; 
32'd172457: dataIn1 = 32'd7784
; 
32'd172458: dataIn1 = 32'd7795
; 
32'd172459: dataIn1 = 32'd7798
; 
32'd172460: dataIn1 = 32'd7799
; 
32'd172461: dataIn1 = 32'd7804
; 
32'd172462: dataIn1 = 32'd5172
; 
32'd172463: dataIn1 = 32'd6299
; 
32'd172464: dataIn1 = 32'd7635
; 
32'd172465: dataIn1 = 32'd7796
; 
32'd172466: dataIn1 = 32'd7800
; 
32'd172467: dataIn1 = 32'd7801
; 
32'd172468: dataIn1 = 32'd7810
; 
32'd172469: dataIn1 = 32'd5172
; 
32'd172470: dataIn1 = 32'd6297
; 
32'd172471: dataIn1 = 32'd6763
; 
32'd172472: dataIn1 = 32'd7796
; 
32'd172473: dataIn1 = 32'd7800
; 
32'd172474: dataIn1 = 32'd7801
; 
32'd172475: dataIn1 = 32'd5186
; 
32'd172476: dataIn1 = 32'd6298
; 
32'd172477: dataIn1 = 32'd7797
; 
32'd172478: dataIn1 = 32'd7802
; 
32'd172479: dataIn1 = 32'd7803
; 
32'd172480: dataIn1 = 32'd7806
; 
32'd172481: dataIn1 = 32'd7808
; 
32'd172482: dataIn1 = 32'd5186
; 
32'd172483: dataIn1 = 32'd6297
; 
32'd172484: dataIn1 = 32'd6762
; 
32'd172485: dataIn1 = 32'd7797
; 
32'd172486: dataIn1 = 32'd7802
; 
32'd172487: dataIn1 = 32'd7803
; 
32'd172488: dataIn1 = 32'd6294
; 
32'd172489: dataIn1 = 32'd6298
; 
32'd172490: dataIn1 = 32'd7784
; 
32'd172491: dataIn1 = 32'd7799
; 
32'd172492: dataIn1 = 32'd7804
; 
32'd172493: dataIn1 = 32'd7805
; 
32'd172494: dataIn1 = 32'd7806
; 
32'd172495: dataIn1 = 32'd6294
; 
32'd172496: dataIn1 = 32'd6300
; 
32'd172497: dataIn1 = 32'd7785
; 
32'd172498: dataIn1 = 32'd7804
; 
32'd172499: dataIn1 = 32'd7805
; 
32'd172500: dataIn1 = 32'd7806
; 
32'd172501: dataIn1 = 32'd7807
; 
32'd172502: dataIn1 = 32'd6298
; 
32'd172503: dataIn1 = 32'd6300
; 
32'd172504: dataIn1 = 32'd7802
; 
32'd172505: dataIn1 = 32'd7804
; 
32'd172506: dataIn1 = 32'd7805
; 
32'd172507: dataIn1 = 32'd7806
; 
32'd172508: dataIn1 = 32'd7808
; 
32'd172509: dataIn1 = 32'd2713
; 
32'd172510: dataIn1 = 32'd6300
; 
32'd172511: dataIn1 = 32'd7785
; 
32'd172512: dataIn1 = 32'd7805
; 
32'd172513: dataIn1 = 32'd7807
; 
32'd172514: dataIn1 = 32'd9042
; 
32'd172515: dataIn1 = 32'd9075
; 
32'd172516: dataIn1 = 32'd5186
; 
32'd172517: dataIn1 = 32'd6300
; 
32'd172518: dataIn1 = 32'd7802
; 
32'd172519: dataIn1 = 32'd7806
; 
32'd172520: dataIn1 = 32'd7808
; 
32'd172521: dataIn1 = 32'd9074
; 
32'd172522: dataIn1 = 32'd9077
; 
32'd172523: dataIn1 = 32'd6296
; 
32'd172524: dataIn1 = 32'd6299
; 
32'd172525: dataIn1 = 32'd7791
; 
32'd172526: dataIn1 = 32'd7798
; 
32'd172527: dataIn1 = 32'd7809
; 
32'd172528: dataIn1 = 32'd7810
; 
32'd172529: dataIn1 = 32'd7811
; 
32'd172530: dataIn1 = 32'd6256
; 
32'd172531: dataIn1 = 32'd6299
; 
32'd172532: dataIn1 = 32'd7635
; 
32'd172533: dataIn1 = 32'd7800
; 
32'd172534: dataIn1 = 32'd7809
; 
32'd172535: dataIn1 = 32'd7810
; 
32'd172536: dataIn1 = 32'd7811
; 
32'd172537: dataIn1 = 32'd6256
; 
32'd172538: dataIn1 = 32'd6296
; 
32'd172539: dataIn1 = 32'd7636
; 
32'd172540: dataIn1 = 32'd7793
; 
32'd172541: dataIn1 = 32'd7809
; 
32'd172542: dataIn1 = 32'd7810
; 
32'd172543: dataIn1 = 32'd7811
; 
32'd172544: dataIn1 = 32'd6302
; 
32'd172545: dataIn1 = 32'd6303
; 
32'd172546: dataIn1 = 32'd7812
; 
32'd172547: dataIn1 = 32'd7813
; 
32'd172548: dataIn1 = 32'd7814
; 
32'd172549: dataIn1 = 32'd7815
; 
32'd172550: dataIn1 = 32'd7816
; 
32'd172551: dataIn1 = 32'd6301
; 
32'd172552: dataIn1 = 32'd6303
; 
32'd172553: dataIn1 = 32'd7812
; 
32'd172554: dataIn1 = 32'd7813
; 
32'd172555: dataIn1 = 32'd7814
; 
32'd172556: dataIn1 = 32'd7817
; 
32'd172557: dataIn1 = 32'd7818
; 
32'd172558: dataIn1 = 32'd6301
; 
32'd172559: dataIn1 = 32'd6302
; 
32'd172560: dataIn1 = 32'd7812
; 
32'd172561: dataIn1 = 32'd7813
; 
32'd172562: dataIn1 = 32'd7814
; 
32'd172563: dataIn1 = 32'd7819
; 
32'd172564: dataIn1 = 32'd7820
; 
32'd172565: dataIn1 = 32'd5174
; 
32'd172566: dataIn1 = 32'd6303
; 
32'd172567: dataIn1 = 32'd7661
; 
32'd172568: dataIn1 = 32'd7812
; 
32'd172569: dataIn1 = 32'd7815
; 
32'd172570: dataIn1 = 32'd7816
; 
32'd172571: dataIn1 = 32'd7831
; 
32'd172572: dataIn1 = 32'd5174
; 
32'd172573: dataIn1 = 32'd6302
; 
32'd172574: dataIn1 = 32'd7654
; 
32'd172575: dataIn1 = 32'd7812
; 
32'd172576: dataIn1 = 32'd7815
; 
32'd172577: dataIn1 = 32'd7816
; 
32'd172578: dataIn1 = 32'd7826
; 
32'd172579: dataIn1 = 32'd5184
; 
32'd172580: dataIn1 = 32'd6303
; 
32'd172581: dataIn1 = 32'd7792
; 
32'd172582: dataIn1 = 32'd7813
; 
32'd172583: dataIn1 = 32'd7817
; 
32'd172584: dataIn1 = 32'd7818
; 
32'd172585: dataIn1 = 32'd7832
; 
32'd172586: dataIn1 = 32'd5184
; 
32'd172587: dataIn1 = 32'd6301
; 
32'd172588: dataIn1 = 32'd7779
; 
32'd172589: dataIn1 = 32'd7813
; 
32'd172590: dataIn1 = 32'd7817
; 
32'd172591: dataIn1 = 32'd7818
; 
32'd172592: dataIn1 = 32'd7822
; 
32'd172593: dataIn1 = 32'd2650
; 
32'd172594: dataIn1 = 32'd6302
; 
32'd172595: dataIn1 = 32'd7814
; 
32'd172596: dataIn1 = 32'd7819
; 
32'd172597: dataIn1 = 32'd7820
; 
32'd172598: dataIn1 = 32'd7828
; 
32'd172599: dataIn1 = 32'd7830
; 
32'd172600: dataIn1 = 32'd2650
; 
32'd172601: dataIn1 = 32'd6301
; 
32'd172602: dataIn1 = 32'd7814
; 
32'd172603: dataIn1 = 32'd7819
; 
32'd172604: dataIn1 = 32'd7820
; 
32'd172605: dataIn1 = 32'd7823
; 
32'd172606: dataIn1 = 32'd7825
; 
32'd172607: dataIn1 = 32'd4954
; 
32'd172608: dataIn1 = 32'd6292
; 
32'd172609: dataIn1 = 32'd7777
; 
32'd172610: dataIn1 = 32'd7821
; 
32'd172611: dataIn1 = 32'd7822
; 
32'd172612: dataIn1 = 32'd7823
; 
32'd172613: dataIn1 = 32'd7824
; 
32'd172614: dataIn1 = 32'd6292
; 
32'd172615: dataIn1 = 32'd6301
; 
32'd172616: dataIn1 = 32'd7779
; 
32'd172617: dataIn1 = 32'd7818
; 
32'd172618: dataIn1 = 32'd7821
; 
32'd172619: dataIn1 = 32'd7822
; 
32'd172620: dataIn1 = 32'd7823
; 
32'd172621: dataIn1 = 32'd4954
; 
32'd172622: dataIn1 = 32'd6301
; 
32'd172623: dataIn1 = 32'd7820
; 
32'd172624: dataIn1 = 32'd7821
; 
32'd172625: dataIn1 = 32'd7822
; 
32'd172626: dataIn1 = 32'd7823
; 
32'd172627: dataIn1 = 32'd7825
; 
32'd172628: dataIn1 = 32'd1110
; 
32'd172629: dataIn1 = 32'd4947
; 
32'd172630: dataIn1 = 32'd4954
; 
32'd172631: dataIn1 = 32'd7777
; 
32'd172632: dataIn1 = 32'd7821
; 
32'd172633: dataIn1 = 32'd7824
; 
32'd172634: dataIn1 = 32'd2650
; 
32'd172635: dataIn1 = 32'd4951
; 
32'd172636: dataIn1 = 32'd4954
; 
32'd172637: dataIn1 = 32'd7820
; 
32'd172638: dataIn1 = 32'd7823
; 
32'd172639: dataIn1 = 32'd7825
; 
32'd172640: dataIn1 = 32'd6263
; 
32'd172641: dataIn1 = 32'd6302
; 
32'd172642: dataIn1 = 32'd7654
; 
32'd172643: dataIn1 = 32'd7816
; 
32'd172644: dataIn1 = 32'd7826
; 
32'd172645: dataIn1 = 32'd7827
; 
32'd172646: dataIn1 = 32'd7828
; 
32'd172647: dataIn1 = 32'd4953
; 
32'd172648: dataIn1 = 32'd6263
; 
32'd172649: dataIn1 = 32'd7655
; 
32'd172650: dataIn1 = 32'd7826
; 
32'd172651: dataIn1 = 32'd7827
; 
32'd172652: dataIn1 = 32'd7828
; 
32'd172653: dataIn1 = 32'd7829
; 
32'd172654: dataIn1 = 32'd4953
; 
32'd172655: dataIn1 = 32'd6302
; 
32'd172656: dataIn1 = 32'd7819
; 
32'd172657: dataIn1 = 32'd7826
; 
32'd172658: dataIn1 = 32'd7827
; 
32'd172659: dataIn1 = 32'd7828
; 
32'd172660: dataIn1 = 32'd7830
; 
32'd172661: dataIn1 = 32'd136
; 
32'd172662: dataIn1 = 32'd4953
; 
32'd172663: dataIn1 = 32'd7655
; 
32'd172664: dataIn1 = 32'd7827
; 
32'd172665: dataIn1 = 32'd7829
; 
32'd172666: dataIn1 = 32'd9609
; 
32'd172667: dataIn1 = 32'd9665
; 
32'd172668: dataIn1 = 32'd2650
; 
32'd172669: dataIn1 = 32'd4953
; 
32'd172670: dataIn1 = 32'd7819
; 
32'd172671: dataIn1 = 32'd7828
; 
32'd172672: dataIn1 = 32'd7830
; 
32'd172673: dataIn1 = 32'd9667
; 
32'd172674: dataIn1 = 32'd9764
; 
32'd172675: dataIn1 = 32'd6264
; 
32'd172676: dataIn1 = 32'd6303
; 
32'd172677: dataIn1 = 32'd7661
; 
32'd172678: dataIn1 = 32'd7815
; 
32'd172679: dataIn1 = 32'd7831
; 
32'd172680: dataIn1 = 32'd7832
; 
32'd172681: dataIn1 = 32'd7833
; 
32'd172682: dataIn1 = 32'd6295
; 
32'd172683: dataIn1 = 32'd6303
; 
32'd172684: dataIn1 = 32'd7792
; 
32'd172685: dataIn1 = 32'd7817
; 
32'd172686: dataIn1 = 32'd7831
; 
32'd172687: dataIn1 = 32'd7832
; 
32'd172688: dataIn1 = 32'd7833
; 
32'd172689: dataIn1 = 32'd6264
; 
32'd172690: dataIn1 = 32'd6295
; 
32'd172691: dataIn1 = 32'd7662
; 
32'd172692: dataIn1 = 32'd7794
; 
32'd172693: dataIn1 = 32'd7831
; 
32'd172694: dataIn1 = 32'd7832
; 
32'd172695: dataIn1 = 32'd7833
; 
32'd172696: dataIn1 = 32'd6305
; 
32'd172697: dataIn1 = 32'd6306
; 
32'd172698: dataIn1 = 32'd7834
; 
32'd172699: dataIn1 = 32'd7835
; 
32'd172700: dataIn1 = 32'd7836
; 
32'd172701: dataIn1 = 32'd7837
; 
32'd172702: dataIn1 = 32'd7838
; 
32'd172703: dataIn1 = 32'd6304
; 
32'd172704: dataIn1 = 32'd6306
; 
32'd172705: dataIn1 = 32'd7834
; 
32'd172706: dataIn1 = 32'd7835
; 
32'd172707: dataIn1 = 32'd7836
; 
32'd172708: dataIn1 = 32'd7839
; 
32'd172709: dataIn1 = 32'd7840
; 
32'd172710: dataIn1 = 32'd6304
; 
32'd172711: dataIn1 = 32'd6305
; 
32'd172712: dataIn1 = 32'd7834
; 
32'd172713: dataIn1 = 32'd7835
; 
32'd172714: dataIn1 = 32'd7836
; 
32'd172715: dataIn1 = 32'd7841
; 
32'd172716: dataIn1 = 32'd7842
; 
32'd172717: dataIn1 = 32'd5187
; 
32'd172718: dataIn1 = 32'd6306
; 
32'd172719: dataIn1 = 32'd7834
; 
32'd172720: dataIn1 = 32'd7837
; 
32'd172721: dataIn1 = 32'd7838
; 
32'd172722: dataIn1 = 32'd7853
; 
32'd172723: dataIn1 = 32'd7856
; 
32'd172724: dataIn1 = 32'd5187
; 
32'd172725: dataIn1 = 32'd6305
; 
32'd172726: dataIn1 = 32'd7834
; 
32'd172727: dataIn1 = 32'd7837
; 
32'd172728: dataIn1 = 32'd7838
; 
32'd172729: dataIn1 = 32'd7848
; 
32'd172730: dataIn1 = 32'd7851
; 
32'd172731: dataIn1 = 32'd2651
; 
32'd172732: dataIn1 = 32'd6306
; 
32'd172733: dataIn1 = 32'd7835
; 
32'd172734: dataIn1 = 32'd7839
; 
32'd172735: dataIn1 = 32'd7840
; 
32'd172736: dataIn1 = 32'd7854
; 
32'd172737: dataIn1 = 32'd7857
; 
32'd172738: dataIn1 = 32'd2651
; 
32'd172739: dataIn1 = 32'd6304
; 
32'd172740: dataIn1 = 32'd7835
; 
32'd172741: dataIn1 = 32'd7839
; 
32'd172742: dataIn1 = 32'd7840
; 
32'd172743: dataIn1 = 32'd7844
; 
32'd172744: dataIn1 = 32'd7847
; 
32'd172745: dataIn1 = 32'd5185
; 
32'd172746: dataIn1 = 32'd6305
; 
32'd172747: dataIn1 = 32'd7787
; 
32'd172748: dataIn1 = 32'd7836
; 
32'd172749: dataIn1 = 32'd7841
; 
32'd172750: dataIn1 = 32'd7842
; 
32'd172751: dataIn1 = 32'd7850
; 
32'd172752: dataIn1 = 32'd5185
; 
32'd172753: dataIn1 = 32'd6304
; 
32'd172754: dataIn1 = 32'd7780
; 
32'd172755: dataIn1 = 32'd7836
; 
32'd172756: dataIn1 = 32'd7841
; 
32'd172757: dataIn1 = 32'd7842
; 
32'd172758: dataIn1 = 32'd7845
; 
32'd172759: dataIn1 = 32'd4958
; 
32'd172760: dataIn1 = 32'd6291
; 
32'd172761: dataIn1 = 32'd7778
; 
32'd172762: dataIn1 = 32'd7843
; 
32'd172763: dataIn1 = 32'd7844
; 
32'd172764: dataIn1 = 32'd7845
; 
32'd172765: dataIn1 = 32'd7846
; 
32'd172766: dataIn1 = 32'd4958
; 
32'd172767: dataIn1 = 32'd6304
; 
32'd172768: dataIn1 = 32'd7840
; 
32'd172769: dataIn1 = 32'd7843
; 
32'd172770: dataIn1 = 32'd7844
; 
32'd172771: dataIn1 = 32'd7845
; 
32'd172772: dataIn1 = 32'd7847
; 
32'd172773: dataIn1 = 32'd6291
; 
32'd172774: dataIn1 = 32'd6304
; 
32'd172775: dataIn1 = 32'd7780
; 
32'd172776: dataIn1 = 32'd7842
; 
32'd172777: dataIn1 = 32'd7843
; 
32'd172778: dataIn1 = 32'd7844
; 
32'd172779: dataIn1 = 32'd7845
; 
32'd172780: dataIn1 = 32'd1110
; 
32'd172781: dataIn1 = 32'd4946
; 
32'd172782: dataIn1 = 32'd4958
; 
32'd172783: dataIn1 = 32'd7778
; 
32'd172784: dataIn1 = 32'd7843
; 
32'd172785: dataIn1 = 32'd7846
; 
32'd172786: dataIn1 = 32'd2651
; 
32'd172787: dataIn1 = 32'd4956
; 
32'd172788: dataIn1 = 32'd4958
; 
32'd172789: dataIn1 = 32'd7840
; 
32'd172790: dataIn1 = 32'd7844
; 
32'd172791: dataIn1 = 32'd7847
; 
32'd172792: dataIn1 = 32'd6305
; 
32'd172793: dataIn1 = 32'd6307
; 
32'd172794: dataIn1 = 32'd7838
; 
32'd172795: dataIn1 = 32'd7848
; 
32'd172796: dataIn1 = 32'd7849
; 
32'd172797: dataIn1 = 32'd7850
; 
32'd172798: dataIn1 = 32'd7851
; 
32'd172799: dataIn1 = 32'd6293
; 
32'd172800: dataIn1 = 32'd6307
; 
32'd172801: dataIn1 = 32'd7786
; 
32'd172802: dataIn1 = 32'd7848
; 
32'd172803: dataIn1 = 32'd7849
; 
32'd172804: dataIn1 = 32'd7850
; 
32'd172805: dataIn1 = 32'd7852
; 
32'd172806: dataIn1 = 32'd6293
; 
32'd172807: dataIn1 = 32'd6305
; 
32'd172808: dataIn1 = 32'd7787
; 
32'd172809: dataIn1 = 32'd7841
; 
32'd172810: dataIn1 = 32'd7848
; 
32'd172811: dataIn1 = 32'd7849
; 
32'd172812: dataIn1 = 32'd7850
; 
32'd172813: dataIn1 = 32'd5187
; 
32'd172814: dataIn1 = 32'd6307
; 
32'd172815: dataIn1 = 32'd7838
; 
32'd172816: dataIn1 = 32'd7848
; 
32'd172817: dataIn1 = 32'd7851
; 
32'd172818: dataIn1 = 32'd9058
; 
32'd172819: dataIn1 = 32'd9065
; 
32'd172820: dataIn1 = 32'd2713
; 
32'd172821: dataIn1 = 32'd6307
; 
32'd172822: dataIn1 = 32'd7786
; 
32'd172823: dataIn1 = 32'd7849
; 
32'd172824: dataIn1 = 32'd7852
; 
32'd172825: dataIn1 = 32'd9041
; 
32'd172826: dataIn1 = 32'd9064
; 
32'd172827: dataIn1 = 32'd6306
; 
32'd172828: dataIn1 = 32'd6308
; 
32'd172829: dataIn1 = 32'd7837
; 
32'd172830: dataIn1 = 32'd7853
; 
32'd172831: dataIn1 = 32'd7854
; 
32'd172832: dataIn1 = 32'd7855
; 
32'd172833: dataIn1 = 32'd7856
; 
32'd172834: dataIn1 = 32'd4959
; 
32'd172835: dataIn1 = 32'd6306
; 
32'd172836: dataIn1 = 32'd7839
; 
32'd172837: dataIn1 = 32'd7853
; 
32'd172838: dataIn1 = 32'd7854
; 
32'd172839: dataIn1 = 32'd7855
; 
32'd172840: dataIn1 = 32'd7857
; 
32'd172841: dataIn1 = 32'd4959
; 
32'd172842: dataIn1 = 32'd6308
; 
32'd172843: dataIn1 = 32'd7853
; 
32'd172844: dataIn1 = 32'd7854
; 
32'd172845: dataIn1 = 32'd7855
; 
32'd172846: dataIn1 = 32'd7858
; 
32'd172847: dataIn1 = 32'd7859
; 
32'd172848: dataIn1 = 32'd5187
; 
32'd172849: dataIn1 = 32'd6308
; 
32'd172850: dataIn1 = 32'd7837
; 
32'd172851: dataIn1 = 32'd7853
; 
32'd172852: dataIn1 = 32'd7856
; 
32'd172853: dataIn1 = 32'd9059
; 
32'd172854: dataIn1 = 32'd9062
; 
32'd172855: dataIn1 = 32'd2651
; 
32'd172856: dataIn1 = 32'd4957
; 
32'd172857: dataIn1 = 32'd4959
; 
32'd172858: dataIn1 = 32'd7839
; 
32'd172859: dataIn1 = 32'd7854
; 
32'd172860: dataIn1 = 32'd7857
; 
32'd172861: dataIn1 = 32'd8
; 
32'd172862: dataIn1 = 32'd6308
; 
32'd172863: dataIn1 = 32'd7855
; 
32'd172864: dataIn1 = 32'd7858
; 
32'd172865: dataIn1 = 32'd7859
; 
32'd172866: dataIn1 = 32'd7966
; 
32'd172867: dataIn1 = 32'd9060
; 
32'd172868: dataIn1 = 32'd8
; 
32'd172869: dataIn1 = 32'd4716
; 
32'd172870: dataIn1 = 32'd4959
; 
32'd172871: dataIn1 = 32'd7855
; 
32'd172872: dataIn1 = 32'd7858
; 
32'd172873: dataIn1 = 32'd7859
; 
32'd172874: dataIn1 = 32'd6310
; 
32'd172875: dataIn1 = 32'd6311
; 
32'd172876: dataIn1 = 32'd7860
; 
32'd172877: dataIn1 = 32'd7861
; 
32'd172878: dataIn1 = 32'd7862
; 
32'd172879: dataIn1 = 32'd7863
; 
32'd172880: dataIn1 = 32'd7864
; 
32'd172881: dataIn1 = 32'd6309
; 
32'd172882: dataIn1 = 32'd6311
; 
32'd172883: dataIn1 = 32'd7860
; 
32'd172884: dataIn1 = 32'd7861
; 
32'd172885: dataIn1 = 32'd7862
; 
32'd172886: dataIn1 = 32'd7865
; 
32'd172887: dataIn1 = 32'd7866
; 
32'd172888: dataIn1 = 32'd6309
; 
32'd172889: dataIn1 = 32'd6310
; 
32'd172890: dataIn1 = 32'd7860
; 
32'd172891: dataIn1 = 32'd7861
; 
32'd172892: dataIn1 = 32'd7862
; 
32'd172893: dataIn1 = 32'd7867
; 
32'd172894: dataIn1 = 32'd7868
; 
32'd172895: dataIn1 = 32'd5188
; 
32'd172896: dataIn1 = 32'd6311
; 
32'd172897: dataIn1 = 32'd7860
; 
32'd172898: dataIn1 = 32'd7863
; 
32'd172899: dataIn1 = 32'd7864
; 
32'd172900: dataIn1 = 32'd7876
; 
32'd172901: dataIn1 = 32'd7879
; 
32'd172902: dataIn1 = 32'd5188
; 
32'd172903: dataIn1 = 32'd6310
; 
32'd172904: dataIn1 = 32'd6315
; 
32'd172905: dataIn1 = 32'd7860
; 
32'd172906: dataIn1 = 32'd7863
; 
32'd172907: dataIn1 = 32'd7864
; 
32'd172908: dataIn1 = 32'd5189
; 
32'd172909: dataIn1 = 32'd6311
; 
32'd172910: dataIn1 = 32'd7861
; 
32'd172911: dataIn1 = 32'd7865
; 
32'd172912: dataIn1 = 32'd7866
; 
32'd172913: dataIn1 = 32'd7877
; 
32'd172914: dataIn1 = 32'd7880
; 
32'd172915: dataIn1 = 32'd5189
; 
32'd172916: dataIn1 = 32'd6309
; 
32'd172917: dataIn1 = 32'd7861
; 
32'd172918: dataIn1 = 32'd7865
; 
32'd172919: dataIn1 = 32'd7866
; 
32'd172920: dataIn1 = 32'd7870
; 
32'd172921: dataIn1 = 32'd7874
; 
32'd172922: dataIn1 = 32'd5190
; 
32'd172923: dataIn1 = 32'd6310
; 
32'd172924: dataIn1 = 32'd6314
; 
32'd172925: dataIn1 = 32'd7862
; 
32'd172926: dataIn1 = 32'd7867
; 
32'd172927: dataIn1 = 32'd7868
; 
32'd172928: dataIn1 = 32'd5190
; 
32'd172929: dataIn1 = 32'd6309
; 
32'd172930: dataIn1 = 32'd7862
; 
32'd172931: dataIn1 = 32'd7867
; 
32'd172932: dataIn1 = 32'd7868
; 
32'd172933: dataIn1 = 32'd7871
; 
32'd172934: dataIn1 = 32'd7875
; 
32'd172935: dataIn1 = 32'd6312
; 
32'd172936: dataIn1 = 32'd6313
; 
32'd172937: dataIn1 = 32'd7869
; 
32'd172938: dataIn1 = 32'd7870
; 
32'd172939: dataIn1 = 32'd7871
; 
32'd172940: dataIn1 = 32'd7872
; 
32'd172941: dataIn1 = 32'd7873
; 
32'd172942: dataIn1 = 32'd6309
; 
32'd172943: dataIn1 = 32'd6313
; 
32'd172944: dataIn1 = 32'd7866
; 
32'd172945: dataIn1 = 32'd7869
; 
32'd172946: dataIn1 = 32'd7870
; 
32'd172947: dataIn1 = 32'd7871
; 
32'd172948: dataIn1 = 32'd7874
; 
32'd172949: dataIn1 = 32'd6309
; 
32'd172950: dataIn1 = 32'd6312
; 
32'd172951: dataIn1 = 32'd7868
; 
32'd172952: dataIn1 = 32'd7869
; 
32'd172953: dataIn1 = 32'd7870
; 
32'd172954: dataIn1 = 32'd7871
; 
32'd172955: dataIn1 = 32'd7875
; 
32'd172956: dataIn1 = 32'd2714
; 
32'd172957: dataIn1 = 32'd6313
; 
32'd172958: dataIn1 = 32'd7869
; 
32'd172959: dataIn1 = 32'd7872
; 
32'd172960: dataIn1 = 32'd7873
; 
32'd172961: dataIn1 = 32'd7899
; 
32'd172962: dataIn1 = 32'd7902
; 
32'd172963: dataIn1 = 32'd2714
; 
32'd172964: dataIn1 = 32'd6312
; 
32'd172965: dataIn1 = 32'd7869
; 
32'd172966: dataIn1 = 32'd7872
; 
32'd172967: dataIn1 = 32'd7873
; 
32'd172968: dataIn1 = 32'd7916
; 
32'd172969: dataIn1 = 32'd7919
; 
32'd172970: dataIn1 = 32'd5189
; 
32'd172971: dataIn1 = 32'd6313
; 
32'd172972: dataIn1 = 32'd7866
; 
32'd172973: dataIn1 = 32'd7870
; 
32'd172974: dataIn1 = 32'd7874
; 
32'd172975: dataIn1 = 32'd7896
; 
32'd172976: dataIn1 = 32'd7900
; 
32'd172977: dataIn1 = 32'd5190
; 
32'd172978: dataIn1 = 32'd6312
; 
32'd172979: dataIn1 = 32'd7868
; 
32'd172980: dataIn1 = 32'd7871
; 
32'd172981: dataIn1 = 32'd7875
; 
32'd172982: dataIn1 = 32'd7918
; 
32'd172983: dataIn1 = 32'd7922
; 
32'd172984: dataIn1 = 32'd6311
; 
32'd172985: dataIn1 = 32'd6317
; 
32'd172986: dataIn1 = 32'd7863
; 
32'd172987: dataIn1 = 32'd7876
; 
32'd172988: dataIn1 = 32'd7877
; 
32'd172989: dataIn1 = 32'd7878
; 
32'd172990: dataIn1 = 32'd7879
; 
32'd172991: dataIn1 = 32'd6311
; 
32'd172992: dataIn1 = 32'd6316
; 
32'd172993: dataIn1 = 32'd7865
; 
32'd172994: dataIn1 = 32'd7876
; 
32'd172995: dataIn1 = 32'd7877
; 
32'd172996: dataIn1 = 32'd7878
; 
32'd172997: dataIn1 = 32'd7880
; 
32'd172998: dataIn1 = 32'd6316
; 
32'd172999: dataIn1 = 32'd6317
; 
32'd173000: dataIn1 = 32'd7876
; 
32'd173001: dataIn1 = 32'd7877
; 
32'd173002: dataIn1 = 32'd7878
; 
32'd173003: dataIn1 = 32'd7881
; 
32'd173004: dataIn1 = 32'd7882
; 
32'd173005: dataIn1 = 32'd5188
; 
32'd173006: dataIn1 = 32'd6317
; 
32'd173007: dataIn1 = 32'd7863
; 
32'd173008: dataIn1 = 32'd7876
; 
32'd173009: dataIn1 = 32'd7879
; 
32'd173010: dataIn1 = 32'd7883
; 
32'd173011: dataIn1 = 32'd7886
; 
32'd173012: dataIn1 = 32'd5189
; 
32'd173013: dataIn1 = 32'd6316
; 
32'd173014: dataIn1 = 32'd7865
; 
32'd173015: dataIn1 = 32'd7877
; 
32'd173016: dataIn1 = 32'd7880
; 
32'd173017: dataIn1 = 32'd7895
; 
32'd173018: dataIn1 = 32'd7912
; 
32'd173019: dataIn1 = 32'd2716
; 
32'd173020: dataIn1 = 32'd6317
; 
32'd173021: dataIn1 = 32'd7878
; 
32'd173022: dataIn1 = 32'd7881
; 
32'd173023: dataIn1 = 32'd7882
; 
32'd173024: dataIn1 = 32'd7885
; 
32'd173025: dataIn1 = 32'd7889
; 
32'd173026: dataIn1 = 32'd2716
; 
32'd173027: dataIn1 = 32'd6316
; 
32'd173028: dataIn1 = 32'd7878
; 
32'd173029: dataIn1 = 32'd7881
; 
32'd173030: dataIn1 = 32'd7882
; 
32'd173031: dataIn1 = 32'd7913
; 
32'd173032: dataIn1 = 32'd7915
; 
32'd173033: dataIn1 = 32'd6317
; 
32'd173034: dataIn1 = 32'd6324
; 
32'd173035: dataIn1 = 32'd7879
; 
32'd173036: dataIn1 = 32'd7883
; 
32'd173037: dataIn1 = 32'd7884
; 
32'd173038: dataIn1 = 32'd7885
; 
32'd173039: dataIn1 = 32'd7886
; 
32'd173040: dataIn1 = 32'd6323
; 
32'd173041: dataIn1 = 32'd6324
; 
32'd173042: dataIn1 = 32'd7883
; 
32'd173043: dataIn1 = 32'd7884
; 
32'd173044: dataIn1 = 32'd7885
; 
32'd173045: dataIn1 = 32'd7887
; 
32'd173046: dataIn1 = 32'd7888
; 
32'd173047: dataIn1 = 32'd6317
; 
32'd173048: dataIn1 = 32'd6323
; 
32'd173049: dataIn1 = 32'd7881
; 
32'd173050: dataIn1 = 32'd7883
; 
32'd173051: dataIn1 = 32'd7884
; 
32'd173052: dataIn1 = 32'd7885
; 
32'd173053: dataIn1 = 32'd7889
; 
32'd173054: dataIn1 = 32'd5188
; 
32'd173055: dataIn1 = 32'd6322
; 
32'd173056: dataIn1 = 32'd6324
; 
32'd173057: dataIn1 = 32'd7879
; 
32'd173058: dataIn1 = 32'd7883
; 
32'd173059: dataIn1 = 32'd7886
; 
32'd173060: dataIn1 = 32'd5191
; 
32'd173061: dataIn1 = 32'd6318
; 
32'd173062: dataIn1 = 32'd6324
; 
32'd173063: dataIn1 = 32'd7884
; 
32'd173064: dataIn1 = 32'd7887
; 
32'd173065: dataIn1 = 32'd7888
; 
32'd173066: dataIn1 = 32'd5191
; 
32'd173067: dataIn1 = 32'd6323
; 
32'd173068: dataIn1 = 32'd7884
; 
32'd173069: dataIn1 = 32'd7887
; 
32'd173070: dataIn1 = 32'd7888
; 
32'd173071: dataIn1 = 32'd8053
; 
32'd173072: dataIn1 = 32'd8063
; 
32'd173073: dataIn1 = 32'd2716
; 
32'd173074: dataIn1 = 32'd6323
; 
32'd173075: dataIn1 = 32'd7881
; 
32'd173076: dataIn1 = 32'd7885
; 
32'd173077: dataIn1 = 32'd7889
; 
32'd173078: dataIn1 = 32'd8046
; 
32'd173079: dataIn1 = 32'd8064
; 
32'd173080: dataIn1 = 32'd6326
; 
32'd173081: dataIn1 = 32'd6327
; 
32'd173082: dataIn1 = 32'd7890
; 
32'd173083: dataIn1 = 32'd7891
; 
32'd173084: dataIn1 = 32'd7892
; 
32'd173085: dataIn1 = 32'd7893
; 
32'd173086: dataIn1 = 32'd7894
; 
32'd173087: dataIn1 = 32'd6325
; 
32'd173088: dataIn1 = 32'd6327
; 
32'd173089: dataIn1 = 32'd7890
; 
32'd173090: dataIn1 = 32'd7891
; 
32'd173091: dataIn1 = 32'd7892
; 
32'd173092: dataIn1 = 32'd7895
; 
32'd173093: dataIn1 = 32'd7896
; 
32'd173094: dataIn1 = 32'd6325
; 
32'd173095: dataIn1 = 32'd6326
; 
32'd173096: dataIn1 = 32'd7890
; 
32'd173097: dataIn1 = 32'd7891
; 
32'd173098: dataIn1 = 32'd7892
; 
32'd173099: dataIn1 = 32'd7897
; 
32'd173100: dataIn1 = 32'd7898
; 
32'd173101: dataIn1 = 32'd5193
; 
32'd173102: dataIn1 = 32'd6327
; 
32'd173103: dataIn1 = 32'd7890
; 
32'd173104: dataIn1 = 32'd7893
; 
32'd173105: dataIn1 = 32'd7894
; 
32'd173106: dataIn1 = 32'd7911
; 
32'd173107: dataIn1 = 32'd7914
; 
32'd173108: dataIn1 = 32'd5193
; 
32'd173109: dataIn1 = 32'd6326
; 
32'd173110: dataIn1 = 32'd7890
; 
32'd173111: dataIn1 = 32'd7893
; 
32'd173112: dataIn1 = 32'd7894
; 
32'd173113: dataIn1 = 32'd7904
; 
32'd173114: dataIn1 = 32'd7907
; 
32'd173115: dataIn1 = 32'd5189
; 
32'd173116: dataIn1 = 32'd6327
; 
32'd173117: dataIn1 = 32'd7880
; 
32'd173118: dataIn1 = 32'd7891
; 
32'd173119: dataIn1 = 32'd7895
; 
32'd173120: dataIn1 = 32'd7896
; 
32'd173121: dataIn1 = 32'd7912
; 
32'd173122: dataIn1 = 32'd5189
; 
32'd173123: dataIn1 = 32'd6325
; 
32'd173124: dataIn1 = 32'd7874
; 
32'd173125: dataIn1 = 32'd7891
; 
32'd173126: dataIn1 = 32'd7895
; 
32'd173127: dataIn1 = 32'd7896
; 
32'd173128: dataIn1 = 32'd7900
; 
32'd173129: dataIn1 = 32'd5194
; 
32'd173130: dataIn1 = 32'd6326
; 
32'd173131: dataIn1 = 32'd7892
; 
32'd173132: dataIn1 = 32'd7897
; 
32'd173133: dataIn1 = 32'd7898
; 
32'd173134: dataIn1 = 32'd7906
; 
32'd173135: dataIn1 = 32'd7910
; 
32'd173136: dataIn1 = 32'd5194
; 
32'd173137: dataIn1 = 32'd6325
; 
32'd173138: dataIn1 = 32'd7892
; 
32'd173139: dataIn1 = 32'd7897
; 
32'd173140: dataIn1 = 32'd7898
; 
32'd173141: dataIn1 = 32'd7901
; 
32'd173142: dataIn1 = 32'd7903
; 
32'd173143: dataIn1 = 32'd6313
; 
32'd173144: dataIn1 = 32'd6328
; 
32'd173145: dataIn1 = 32'd7872
; 
32'd173146: dataIn1 = 32'd7899
; 
32'd173147: dataIn1 = 32'd7900
; 
32'd173148: dataIn1 = 32'd7901
; 
32'd173149: dataIn1 = 32'd7902
; 
32'd173150: dataIn1 = 32'd6313
; 
32'd173151: dataIn1 = 32'd6325
; 
32'd173152: dataIn1 = 32'd7874
; 
32'd173153: dataIn1 = 32'd7896
; 
32'd173154: dataIn1 = 32'd7899
; 
32'd173155: dataIn1 = 32'd7900
; 
32'd173156: dataIn1 = 32'd7901
; 
32'd173157: dataIn1 = 32'd6325
; 
32'd173158: dataIn1 = 32'd6328
; 
32'd173159: dataIn1 = 32'd7898
; 
32'd173160: dataIn1 = 32'd7899
; 
32'd173161: dataIn1 = 32'd7900
; 
32'd173162: dataIn1 = 32'd7901
; 
32'd173163: dataIn1 = 32'd7903
; 
32'd173164: dataIn1 = 32'd2714
; 
32'd173165: dataIn1 = 32'd6328
; 
32'd173166: dataIn1 = 32'd7872
; 
32'd173167: dataIn1 = 32'd7899
; 
32'd173168: dataIn1 = 32'd7902
; 
32'd173169: dataIn1 = 32'd7935
; 
32'd173170: dataIn1 = 32'd7988
; 
32'd173171: dataIn1 = 32'd5194
; 
32'd173172: dataIn1 = 32'd6328
; 
32'd173173: dataIn1 = 32'd7898
; 
32'd173174: dataIn1 = 32'd7901
; 
32'd173175: dataIn1 = 32'd7903
; 
32'd173176: dataIn1 = 32'd7987
; 
32'd173177: dataIn1 = 32'd7990
; 
32'd173178: dataIn1 = 32'd6326
; 
32'd173179: dataIn1 = 32'd6330
; 
32'd173180: dataIn1 = 32'd7894
; 
32'd173181: dataIn1 = 32'd7904
; 
32'd173182: dataIn1 = 32'd7905
; 
32'd173183: dataIn1 = 32'd7906
; 
32'd173184: dataIn1 = 32'd7907
; 
32'd173185: dataIn1 = 32'd6329
; 
32'd173186: dataIn1 = 32'd6330
; 
32'd173187: dataIn1 = 32'd7904
; 
32'd173188: dataIn1 = 32'd7905
; 
32'd173189: dataIn1 = 32'd7906
; 
32'd173190: dataIn1 = 32'd7908
; 
32'd173191: dataIn1 = 32'd7909
; 
32'd173192: dataIn1 = 32'd6326
; 
32'd173193: dataIn1 = 32'd6329
; 
32'd173194: dataIn1 = 32'd7897
; 
32'd173195: dataIn1 = 32'd7904
; 
32'd173196: dataIn1 = 32'd7905
; 
32'd173197: dataIn1 = 32'd7906
; 
32'd173198: dataIn1 = 32'd7910
; 
32'd173199: dataIn1 = 32'd5193
; 
32'd173200: dataIn1 = 32'd6330
; 
32'd173201: dataIn1 = 32'd7894
; 
32'd173202: dataIn1 = 32'd7904
; 
32'd173203: dataIn1 = 32'd7907
; 
32'd173204: dataIn1 = 32'd8069
; 
32'd173205: dataIn1 = 32'd8079
; 
32'd173206: dataIn1 = 32'd139
; 
32'd173207: dataIn1 = 32'd6330
; 
32'd173208: dataIn1 = 32'd7905
; 
32'd173209: dataIn1 = 32'd7908
; 
32'd173210: dataIn1 = 32'd7909
; 
32'd173211: dataIn1 = 32'd8080
; 
32'd173212: dataIn1 = 32'd8082
; 
32'd173213: dataIn1 = 32'd139
; 
32'd173214: dataIn1 = 32'd6329
; 
32'd173215: dataIn1 = 32'd7905
; 
32'd173216: dataIn1 = 32'd7908
; 
32'd173217: dataIn1 = 32'd7909
; 
32'd173218: dataIn1 = 32'd7992
; 
32'd173219: dataIn1 = 32'd7995
; 
32'd173220: dataIn1 = 32'd5194
; 
32'd173221: dataIn1 = 32'd6329
; 
32'd173222: dataIn1 = 32'd7897
; 
32'd173223: dataIn1 = 32'd7906
; 
32'd173224: dataIn1 = 32'd7910
; 
32'd173225: dataIn1 = 32'd7986
; 
32'd173226: dataIn1 = 32'd7993
; 
32'd173227: dataIn1 = 32'd6327
; 
32'd173228: dataIn1 = 32'd6331
; 
32'd173229: dataIn1 = 32'd7893
; 
32'd173230: dataIn1 = 32'd7911
; 
32'd173231: dataIn1 = 32'd7912
; 
32'd173232: dataIn1 = 32'd7913
; 
32'd173233: dataIn1 = 32'd7914
; 
32'd173234: dataIn1 = 32'd6316
; 
32'd173235: dataIn1 = 32'd6327
; 
32'd173236: dataIn1 = 32'd7880
; 
32'd173237: dataIn1 = 32'd7895
; 
32'd173238: dataIn1 = 32'd7911
; 
32'd173239: dataIn1 = 32'd7912
; 
32'd173240: dataIn1 = 32'd7913
; 
32'd173241: dataIn1 = 32'd6316
; 
32'd173242: dataIn1 = 32'd6331
; 
32'd173243: dataIn1 = 32'd7882
; 
32'd173244: dataIn1 = 32'd7911
; 
32'd173245: dataIn1 = 32'd7912
; 
32'd173246: dataIn1 = 32'd7913
; 
32'd173247: dataIn1 = 32'd7915
; 
32'd173248: dataIn1 = 32'd5193
; 
32'd173249: dataIn1 = 32'd6331
; 
32'd173250: dataIn1 = 32'd7893
; 
32'd173251: dataIn1 = 32'd7911
; 
32'd173252: dataIn1 = 32'd7914
; 
32'd173253: dataIn1 = 32'd8068
; 
32'd173254: dataIn1 = 32'd8084
; 
32'd173255: dataIn1 = 32'd2716
; 
32'd173256: dataIn1 = 32'd6331
; 
32'd173257: dataIn1 = 32'd7882
; 
32'd173258: dataIn1 = 32'd7913
; 
32'd173259: dataIn1 = 32'd7915
; 
32'd173260: dataIn1 = 32'd8047
; 
32'd173261: dataIn1 = 32'd8086
; 
32'd173262: dataIn1 = 32'd6312
; 
32'd173263: dataIn1 = 32'd6333
; 
32'd173264: dataIn1 = 32'd7873
; 
32'd173265: dataIn1 = 32'd7916
; 
32'd173266: dataIn1 = 32'd7917
; 
32'd173267: dataIn1 = 32'd7918
; 
32'd173268: dataIn1 = 32'd7919
; 
32'd173269: dataIn1 = 32'd6332
; 
32'd173270: dataIn1 = 32'd6333
; 
32'd173271: dataIn1 = 32'd7916
; 
32'd173272: dataIn1 = 32'd7917
; 
32'd173273: dataIn1 = 32'd7918
; 
32'd173274: dataIn1 = 32'd7920
; 
32'd173275: dataIn1 = 32'd7921
; 
32'd173276: dataIn1 = 32'd6312
; 
32'd173277: dataIn1 = 32'd6332
; 
32'd173278: dataIn1 = 32'd7875
; 
32'd173279: dataIn1 = 32'd7916
; 
32'd173280: dataIn1 = 32'd7917
; 
32'd173281: dataIn1 = 32'd7918
; 
32'd173282: dataIn1 = 32'd7922
; 
32'd173283: dataIn1 = 32'd2714
; 
32'd173284: dataIn1 = 32'd6333
; 
32'd173285: dataIn1 = 32'd7873
; 
32'd173286: dataIn1 = 32'd7916
; 
32'd173287: dataIn1 = 32'd7919
; 
32'd173288: dataIn1 = 32'd7936
; 
32'd173289: dataIn1 = 32'd8010
; 
32'd173290: dataIn1 = 32'd5196
; 
32'd173291: dataIn1 = 32'd6333
; 
32'd173292: dataIn1 = 32'd7917
; 
32'd173293: dataIn1 = 32'd7920
; 
32'd173294: dataIn1 = 32'd7921
; 
32'd173295: dataIn1 = 32'd8007
; 
32'd173296: dataIn1 = 32'd8011
; 
32'd173297: dataIn1 = 32'd5196
; 
32'd173298: dataIn1 = 32'd6332
; 
32'd173299: dataIn1 = 32'd6338
; 
32'd173300: dataIn1 = 32'd7917
; 
32'd173301: dataIn1 = 32'd7920
; 
32'd173302: dataIn1 = 32'd7921
; 
32'd173303: dataIn1 = 32'd5190
; 
32'd173304: dataIn1 = 32'd6332
; 
32'd173305: dataIn1 = 32'd6334
; 
32'd173306: dataIn1 = 32'd7875
; 
32'd173307: dataIn1 = 32'd7918
; 
32'd173308: dataIn1 = 32'd7922
; 
32'd173309: dataIn1 = 32'd6340
; 
32'd173310: dataIn1 = 32'd6341
; 
32'd173311: dataIn1 = 32'd7923
; 
32'd173312: dataIn1 = 32'd7924
; 
32'd173313: dataIn1 = 32'd7925
; 
32'd173314: dataIn1 = 32'd7926
; 
32'd173315: dataIn1 = 32'd7927
; 
32'd173316: dataIn1 = 32'd6339
; 
32'd173317: dataIn1 = 32'd6341
; 
32'd173318: dataIn1 = 32'd7923
; 
32'd173319: dataIn1 = 32'd7924
; 
32'd173320: dataIn1 = 32'd7925
; 
32'd173321: dataIn1 = 32'd7928
; 
32'd173322: dataIn1 = 32'd7929
; 
32'd173323: dataIn1 = 32'd6339
; 
32'd173324: dataIn1 = 32'd6340
; 
32'd173325: dataIn1 = 32'd7923
; 
32'd173326: dataIn1 = 32'd7924
; 
32'd173327: dataIn1 = 32'd7925
; 
32'd173328: dataIn1 = 32'd7930
; 
32'd173329: dataIn1 = 32'd7931
; 
32'd173330: dataIn1 = 32'd5197
; 
32'd173331: dataIn1 = 32'd6341
; 
32'd173332: dataIn1 = 32'd7923
; 
32'd173333: dataIn1 = 32'd7926
; 
32'd173334: dataIn1 = 32'd7927
; 
32'd173335: dataIn1 = 32'd7946
; 
32'd173336: dataIn1 = 32'd7949
; 
32'd173337: dataIn1 = 32'd5197
; 
32'd173338: dataIn1 = 32'd6340
; 
32'd173339: dataIn1 = 32'd7923
; 
32'd173340: dataIn1 = 32'd7926
; 
32'd173341: dataIn1 = 32'd7927
; 
32'd173342: dataIn1 = 32'd7939
; 
32'd173343: dataIn1 = 32'd7942
; 
32'd173344: dataIn1 = 32'd5198
; 
32'd173345: dataIn1 = 32'd6341
; 
32'd173346: dataIn1 = 32'd7924
; 
32'd173347: dataIn1 = 32'd7928
; 
32'd173348: dataIn1 = 32'd7929
; 
32'd173349: dataIn1 = 32'd7947
; 
32'd173350: dataIn1 = 32'd7950
; 
32'd173351: dataIn1 = 32'd5198
; 
32'd173352: dataIn1 = 32'd6339
; 
32'd173353: dataIn1 = 32'd7924
; 
32'd173354: dataIn1 = 32'd7928
; 
32'd173355: dataIn1 = 32'd7929
; 
32'd173356: dataIn1 = 32'd7933
; 
32'd173357: dataIn1 = 32'd7937
; 
32'd173358: dataIn1 = 32'd5199
; 
32'd173359: dataIn1 = 32'd6340
; 
32'd173360: dataIn1 = 32'd7925
; 
32'd173361: dataIn1 = 32'd7930
; 
32'd173362: dataIn1 = 32'd7931
; 
32'd173363: dataIn1 = 32'd7941
; 
32'd173364: dataIn1 = 32'd7945
; 
32'd173365: dataIn1 = 32'd5199
; 
32'd173366: dataIn1 = 32'd6339
; 
32'd173367: dataIn1 = 32'd7925
; 
32'd173368: dataIn1 = 32'd7930
; 
32'd173369: dataIn1 = 32'd7931
; 
32'd173370: dataIn1 = 32'd7934
; 
32'd173371: dataIn1 = 32'd7938
; 
32'd173372: dataIn1 = 32'd6342
; 
32'd173373: dataIn1 = 32'd6343
; 
32'd173374: dataIn1 = 32'd7932
; 
32'd173375: dataIn1 = 32'd7933
; 
32'd173376: dataIn1 = 32'd7934
; 
32'd173377: dataIn1 = 32'd7935
; 
32'd173378: dataIn1 = 32'd7936
; 
32'd173379: dataIn1 = 32'd6339
; 
32'd173380: dataIn1 = 32'd6343
; 
32'd173381: dataIn1 = 32'd7929
; 
32'd173382: dataIn1 = 32'd7932
; 
32'd173383: dataIn1 = 32'd7933
; 
32'd173384: dataIn1 = 32'd7934
; 
32'd173385: dataIn1 = 32'd7937
; 
32'd173386: dataIn1 = 32'd6339
; 
32'd173387: dataIn1 = 32'd6342
; 
32'd173388: dataIn1 = 32'd7931
; 
32'd173389: dataIn1 = 32'd7932
; 
32'd173390: dataIn1 = 32'd7933
; 
32'd173391: dataIn1 = 32'd7934
; 
32'd173392: dataIn1 = 32'd7938
; 
32'd173393: dataIn1 = 32'd2714
; 
32'd173394: dataIn1 = 32'd6343
; 
32'd173395: dataIn1 = 32'd7902
; 
32'd173396: dataIn1 = 32'd7932
; 
32'd173397: dataIn1 = 32'd7935
; 
32'd173398: dataIn1 = 32'd7936
; 
32'd173399: dataIn1 = 32'd7988
; 
32'd173400: dataIn1 = 32'd2714
; 
32'd173401: dataIn1 = 32'd6342
; 
32'd173402: dataIn1 = 32'd7919
; 
32'd173403: dataIn1 = 32'd7932
; 
32'd173404: dataIn1 = 32'd7935
; 
32'd173405: dataIn1 = 32'd7936
; 
32'd173406: dataIn1 = 32'd8010
; 
32'd173407: dataIn1 = 32'd5198
; 
32'd173408: dataIn1 = 32'd6343
; 
32'd173409: dataIn1 = 32'd7929
; 
32'd173410: dataIn1 = 32'd7933
; 
32'd173411: dataIn1 = 32'd7937
; 
32'd173412: dataIn1 = 32'd7985
; 
32'd173413: dataIn1 = 32'd7989
; 
32'd173414: dataIn1 = 32'd5199
; 
32'd173415: dataIn1 = 32'd6342
; 
32'd173416: dataIn1 = 32'd7931
; 
32'd173417: dataIn1 = 32'd7934
; 
32'd173418: dataIn1 = 32'd7938
; 
32'd173419: dataIn1 = 32'd8009
; 
32'd173420: dataIn1 = 32'd8012
; 
32'd173421: dataIn1 = 32'd6340
; 
32'd173422: dataIn1 = 32'd6345
; 
32'd173423: dataIn1 = 32'd7927
; 
32'd173424: dataIn1 = 32'd7939
; 
32'd173425: dataIn1 = 32'd7940
; 
32'd173426: dataIn1 = 32'd7941
; 
32'd173427: dataIn1 = 32'd7942
; 
32'd173428: dataIn1 = 32'd6344
; 
32'd173429: dataIn1 = 32'd6345
; 
32'd173430: dataIn1 = 32'd7939
; 
32'd173431: dataIn1 = 32'd7940
; 
32'd173432: dataIn1 = 32'd7941
; 
32'd173433: dataIn1 = 32'd7943
; 
32'd173434: dataIn1 = 32'd7944
; 
32'd173435: dataIn1 = 32'd6340
; 
32'd173436: dataIn1 = 32'd6344
; 
32'd173437: dataIn1 = 32'd7930
; 
32'd173438: dataIn1 = 32'd7939
; 
32'd173439: dataIn1 = 32'd7940
; 
32'd173440: dataIn1 = 32'd7941
; 
32'd173441: dataIn1 = 32'd7945
; 
32'd173442: dataIn1 = 32'd5197
; 
32'd173443: dataIn1 = 32'd6345
; 
32'd173444: dataIn1 = 32'd7927
; 
32'd173445: dataIn1 = 32'd7939
; 
32'd173446: dataIn1 = 32'd7942
; 
32'd173447: dataIn1 = 32'd7957
; 
32'd173448: dataIn1 = 32'd7969
; 
32'd173449: dataIn1 = 32'd2717
; 
32'd173450: dataIn1 = 32'd6345
; 
32'd173451: dataIn1 = 32'd7940
; 
32'd173452: dataIn1 = 32'd7943
; 
32'd173453: dataIn1 = 32'd7944
; 
32'd173454: dataIn1 = 32'd7970
; 
32'd173455: dataIn1 = 32'd7972
; 
32'd173456: dataIn1 = 32'd2717
; 
32'd173457: dataIn1 = 32'd6344
; 
32'd173458: dataIn1 = 32'd7940
; 
32'd173459: dataIn1 = 32'd7943
; 
32'd173460: dataIn1 = 32'd7944
; 
32'd173461: dataIn1 = 32'd8014
; 
32'd173462: dataIn1 = 32'd8017
; 
32'd173463: dataIn1 = 32'd5199
; 
32'd173464: dataIn1 = 32'd6344
; 
32'd173465: dataIn1 = 32'd7930
; 
32'd173466: dataIn1 = 32'd7941
; 
32'd173467: dataIn1 = 32'd7945
; 
32'd173468: dataIn1 = 32'd8008
; 
32'd173469: dataIn1 = 32'd8015
; 
32'd173470: dataIn1 = 32'd6341
; 
32'd173471: dataIn1 = 32'd6347
; 
32'd173472: dataIn1 = 32'd7926
; 
32'd173473: dataIn1 = 32'd7946
; 
32'd173474: dataIn1 = 32'd7947
; 
32'd173475: dataIn1 = 32'd7948
; 
32'd173476: dataIn1 = 32'd7949
; 
32'd173477: dataIn1 = 32'd6341
; 
32'd173478: dataIn1 = 32'd6346
; 
32'd173479: dataIn1 = 32'd7928
; 
32'd173480: dataIn1 = 32'd7946
; 
32'd173481: dataIn1 = 32'd7947
; 
32'd173482: dataIn1 = 32'd7948
; 
32'd173483: dataIn1 = 32'd7950
; 
32'd173484: dataIn1 = 32'd6346
; 
32'd173485: dataIn1 = 32'd6347
; 
32'd173486: dataIn1 = 32'd7946
; 
32'd173487: dataIn1 = 32'd7947
; 
32'd173488: dataIn1 = 32'd7948
; 
32'd173489: dataIn1 = 32'd7951
; 
32'd173490: dataIn1 = 32'd7952
; 
32'd173491: dataIn1 = 32'd5197
; 
32'd173492: dataIn1 = 32'd6347
; 
32'd173493: dataIn1 = 32'd7926
; 
32'd173494: dataIn1 = 32'd7946
; 
32'd173495: dataIn1 = 32'd7949
; 
32'd173496: dataIn1 = 32'd7956
; 
32'd173497: dataIn1 = 32'd7974
; 
32'd173498: dataIn1 = 32'd5198
; 
32'd173499: dataIn1 = 32'd6346
; 
32'd173500: dataIn1 = 32'd7928
; 
32'd173501: dataIn1 = 32'd7947
; 
32'd173502: dataIn1 = 32'd7950
; 
32'd173503: dataIn1 = 32'd7984
; 
32'd173504: dataIn1 = 32'd7997
; 
32'd173505: dataIn1 = 32'd1111
; 
32'd173506: dataIn1 = 32'd6347
; 
32'd173507: dataIn1 = 32'd7948
; 
32'd173508: dataIn1 = 32'd7951
; 
32'd173509: dataIn1 = 32'd7952
; 
32'd173510: dataIn1 = 32'd7976
; 
32'd173511: dataIn1 = 32'd7978
; 
32'd173512: dataIn1 = 32'd1111
; 
32'd173513: dataIn1 = 32'd6346
; 
32'd173514: dataIn1 = 32'd7948
; 
32'd173515: dataIn1 = 32'd7951
; 
32'd173516: dataIn1 = 32'd7952
; 
32'd173517: dataIn1 = 32'd7998
; 
32'd173518: dataIn1 = 32'd8000
; 
32'd173519: dataIn1 = 32'd6349
; 
32'd173520: dataIn1 = 32'd6350
; 
32'd173521: dataIn1 = 32'd7953
; 
32'd173522: dataIn1 = 32'd7954
; 
32'd173523: dataIn1 = 32'd7955
; 
32'd173524: dataIn1 = 32'd7956
; 
32'd173525: dataIn1 = 32'd7957
; 
32'd173526: dataIn1 = 32'd6348
; 
32'd173527: dataIn1 = 32'd6350
; 
32'd173528: dataIn1 = 32'd7953
; 
32'd173529: dataIn1 = 32'd7954
; 
32'd173530: dataIn1 = 32'd7955
; 
32'd173531: dataIn1 = 32'd7958
; 
32'd173532: dataIn1 = 32'd7959
; 
32'd173533: dataIn1 = 32'd6348
; 
32'd173534: dataIn1 = 32'd6349
; 
32'd173535: dataIn1 = 32'd7953
; 
32'd173536: dataIn1 = 32'd7954
; 
32'd173537: dataIn1 = 32'd7955
; 
32'd173538: dataIn1 = 32'd7960
; 
32'd173539: dataIn1 = 32'd7961
; 
32'd173540: dataIn1 = 32'd5197
; 
32'd173541: dataIn1 = 32'd6350
; 
32'd173542: dataIn1 = 32'd7949
; 
32'd173543: dataIn1 = 32'd7953
; 
32'd173544: dataIn1 = 32'd7956
; 
32'd173545: dataIn1 = 32'd7957
; 
32'd173546: dataIn1 = 32'd7974
; 
32'd173547: dataIn1 = 32'd5197
; 
32'd173548: dataIn1 = 32'd6349
; 
32'd173549: dataIn1 = 32'd7942
; 
32'd173550: dataIn1 = 32'd7953
; 
32'd173551: dataIn1 = 32'd7956
; 
32'd173552: dataIn1 = 32'd7957
; 
32'd173553: dataIn1 = 32'd7969
; 
32'd173554: dataIn1 = 32'd2656
; 
32'd173555: dataIn1 = 32'd6350
; 
32'd173556: dataIn1 = 32'd7954
; 
32'd173557: dataIn1 = 32'd7958
; 
32'd173558: dataIn1 = 32'd7959
; 
32'd173559: dataIn1 = 32'd7975
; 
32'd173560: dataIn1 = 32'd7977
; 
32'd173561: dataIn1 = 32'd2656
; 
32'd173562: dataIn1 = 32'd6348
; 
32'd173563: dataIn1 = 32'd7954
; 
32'd173564: dataIn1 = 32'd7958
; 
32'd173565: dataIn1 = 32'd7959
; 
32'd173566: dataIn1 = 32'd7963
; 
32'd173567: dataIn1 = 32'd7967
; 
32'd173568: dataIn1 = 32'd5200
; 
32'd173569: dataIn1 = 32'd6349
; 
32'd173570: dataIn1 = 32'd7955
; 
32'd173571: dataIn1 = 32'd7960
; 
32'd173572: dataIn1 = 32'd7961
; 
32'd173573: dataIn1 = 32'd7971
; 
32'd173574: dataIn1 = 32'd7973
; 
32'd173575: dataIn1 = 32'd5200
; 
32'd173576: dataIn1 = 32'd6348
; 
32'd173577: dataIn1 = 32'd7955
; 
32'd173578: dataIn1 = 32'd7960
; 
32'd173579: dataIn1 = 32'd7961
; 
32'd173580: dataIn1 = 32'd7964
; 
32'd173581: dataIn1 = 32'd7968
; 
32'd173582: dataIn1 = 32'd4977
; 
32'd173583: dataIn1 = 32'd6351
; 
32'd173584: dataIn1 = 32'd7962
; 
32'd173585: dataIn1 = 32'd7963
; 
32'd173586: dataIn1 = 32'd7964
; 
32'd173587: dataIn1 = 32'd7965
; 
32'd173588: dataIn1 = 32'd7966
; 
32'd173589: dataIn1 = 32'd4977
; 
32'd173590: dataIn1 = 32'd6348
; 
32'd173591: dataIn1 = 32'd7959
; 
32'd173592: dataIn1 = 32'd7962
; 
32'd173593: dataIn1 = 32'd7963
; 
32'd173594: dataIn1 = 32'd7964
; 
32'd173595: dataIn1 = 32'd7967
; 
32'd173596: dataIn1 = 32'd6348
; 
32'd173597: dataIn1 = 32'd6351
; 
32'd173598: dataIn1 = 32'd7961
; 
32'd173599: dataIn1 = 32'd7962
; 
32'd173600: dataIn1 = 32'd7963
; 
32'd173601: dataIn1 = 32'd7964
; 
32'd173602: dataIn1 = 32'd7968
; 
32'd173603: dataIn1 = 32'd8
; 
32'd173604: dataIn1 = 32'd4717
; 
32'd173605: dataIn1 = 32'd4977
; 
32'd173606: dataIn1 = 32'd7962
; 
32'd173607: dataIn1 = 32'd7965
; 
32'd173608: dataIn1 = 32'd7966
; 
32'd173609: dataIn1 = 32'd8
; 
32'd173610: dataIn1 = 32'd6351
; 
32'd173611: dataIn1 = 32'd7858
; 
32'd173612: dataIn1 = 32'd7962
; 
32'd173613: dataIn1 = 32'd7965
; 
32'd173614: dataIn1 = 32'd7966
; 
32'd173615: dataIn1 = 32'd9060
; 
32'd173616: dataIn1 = 32'd2656
; 
32'd173617: dataIn1 = 32'd4975
; 
32'd173618: dataIn1 = 32'd4977
; 
32'd173619: dataIn1 = 32'd7959
; 
32'd173620: dataIn1 = 32'd7963
; 
32'd173621: dataIn1 = 32'd7967
; 
32'd173622: dataIn1 = 32'd5200
; 
32'd173623: dataIn1 = 32'd6351
; 
32'd173624: dataIn1 = 32'd7961
; 
32'd173625: dataIn1 = 32'd7964
; 
32'd173626: dataIn1 = 32'd7968
; 
32'd173627: dataIn1 = 32'd9057
; 
32'd173628: dataIn1 = 32'd9061
; 
32'd173629: dataIn1 = 32'd6345
; 
32'd173630: dataIn1 = 32'd6349
; 
32'd173631: dataIn1 = 32'd7942
; 
32'd173632: dataIn1 = 32'd7957
; 
32'd173633: dataIn1 = 32'd7969
; 
32'd173634: dataIn1 = 32'd7970
; 
32'd173635: dataIn1 = 32'd7971
; 
32'd173636: dataIn1 = 32'd6345
; 
32'd173637: dataIn1 = 32'd6352
; 
32'd173638: dataIn1 = 32'd7943
; 
32'd173639: dataIn1 = 32'd7969
; 
32'd173640: dataIn1 = 32'd7970
; 
32'd173641: dataIn1 = 32'd7971
; 
32'd173642: dataIn1 = 32'd7972
; 
32'd173643: dataIn1 = 32'd6349
; 
32'd173644: dataIn1 = 32'd6352
; 
32'd173645: dataIn1 = 32'd7960
; 
32'd173646: dataIn1 = 32'd7969
; 
32'd173647: dataIn1 = 32'd7970
; 
32'd173648: dataIn1 = 32'd7971
; 
32'd173649: dataIn1 = 32'd7973
; 
32'd173650: dataIn1 = 32'd2717
; 
32'd173651: dataIn1 = 32'd6352
; 
32'd173652: dataIn1 = 32'd7943
; 
32'd173653: dataIn1 = 32'd7970
; 
32'd173654: dataIn1 = 32'd7972
; 
32'd173655: dataIn1 = 32'd9049
; 
32'd173656: dataIn1 = 32'd9068
; 
32'd173657: dataIn1 = 32'd5200
; 
32'd173658: dataIn1 = 32'd6352
; 
32'd173659: dataIn1 = 32'd7960
; 
32'd173660: dataIn1 = 32'd7971
; 
32'd173661: dataIn1 = 32'd7973
; 
32'd173662: dataIn1 = 32'd9056
; 
32'd173663: dataIn1 = 32'd9067
; 
32'd173664: dataIn1 = 32'd6347
; 
32'd173665: dataIn1 = 32'd6350
; 
32'd173666: dataIn1 = 32'd7949
; 
32'd173667: dataIn1 = 32'd7956
; 
32'd173668: dataIn1 = 32'd7974
; 
32'd173669: dataIn1 = 32'd7975
; 
32'd173670: dataIn1 = 32'd7976
; 
32'd173671: dataIn1 = 32'd4978
; 
32'd173672: dataIn1 = 32'd6350
; 
32'd173673: dataIn1 = 32'd7958
; 
32'd173674: dataIn1 = 32'd7974
; 
32'd173675: dataIn1 = 32'd7975
; 
32'd173676: dataIn1 = 32'd7976
; 
32'd173677: dataIn1 = 32'd7977
; 
32'd173678: dataIn1 = 32'd4978
; 
32'd173679: dataIn1 = 32'd6347
; 
32'd173680: dataIn1 = 32'd7951
; 
32'd173681: dataIn1 = 32'd7974
; 
32'd173682: dataIn1 = 32'd7975
; 
32'd173683: dataIn1 = 32'd7976
; 
32'd173684: dataIn1 = 32'd7978
; 
32'd173685: dataIn1 = 32'd2656
; 
32'd173686: dataIn1 = 32'd4976
; 
32'd173687: dataIn1 = 32'd4978
; 
32'd173688: dataIn1 = 32'd7958
; 
32'd173689: dataIn1 = 32'd7975
; 
32'd173690: dataIn1 = 32'd7977
; 
32'd173691: dataIn1 = 32'd1111
; 
32'd173692: dataIn1 = 32'd4967
; 
32'd173693: dataIn1 = 32'd4978
; 
32'd173694: dataIn1 = 32'd7951
; 
32'd173695: dataIn1 = 32'd7976
; 
32'd173696: dataIn1 = 32'd7978
; 
32'd173697: dataIn1 = 32'd6354
; 
32'd173698: dataIn1 = 32'd6355
; 
32'd173699: dataIn1 = 32'd7979
; 
32'd173700: dataIn1 = 32'd7980
; 
32'd173701: dataIn1 = 32'd7981
; 
32'd173702: dataIn1 = 32'd7982
; 
32'd173703: dataIn1 = 32'd7983
; 
32'd173704: dataIn1 = 32'd6353
; 
32'd173705: dataIn1 = 32'd6355
; 
32'd173706: dataIn1 = 32'd7979
; 
32'd173707: dataIn1 = 32'd7980
; 
32'd173708: dataIn1 = 32'd7981
; 
32'd173709: dataIn1 = 32'd7984
; 
32'd173710: dataIn1 = 32'd7985
; 
32'd173711: dataIn1 = 32'd6353
; 
32'd173712: dataIn1 = 32'd6354
; 
32'd173713: dataIn1 = 32'd7979
; 
32'd173714: dataIn1 = 32'd7980
; 
32'd173715: dataIn1 = 32'd7981
; 
32'd173716: dataIn1 = 32'd7986
; 
32'd173717: dataIn1 = 32'd7987
; 
32'd173718: dataIn1 = 32'd2655
; 
32'd173719: dataIn1 = 32'd6355
; 
32'd173720: dataIn1 = 32'd7979
; 
32'd173721: dataIn1 = 32'd7982
; 
32'd173722: dataIn1 = 32'd7983
; 
32'd173723: dataIn1 = 32'd7996
; 
32'd173724: dataIn1 = 32'd7999
; 
32'd173725: dataIn1 = 32'd2655
; 
32'd173726: dataIn1 = 32'd6354
; 
32'd173727: dataIn1 = 32'd7979
; 
32'd173728: dataIn1 = 32'd7982
; 
32'd173729: dataIn1 = 32'd7983
; 
32'd173730: dataIn1 = 32'd7991
; 
32'd173731: dataIn1 = 32'd7994
; 
32'd173732: dataIn1 = 32'd5198
; 
32'd173733: dataIn1 = 32'd6355
; 
32'd173734: dataIn1 = 32'd7950
; 
32'd173735: dataIn1 = 32'd7980
; 
32'd173736: dataIn1 = 32'd7984
; 
32'd173737: dataIn1 = 32'd7985
; 
32'd173738: dataIn1 = 32'd7997
; 
32'd173739: dataIn1 = 32'd5198
; 
32'd173740: dataIn1 = 32'd6353
; 
32'd173741: dataIn1 = 32'd7937
; 
32'd173742: dataIn1 = 32'd7980
; 
32'd173743: dataIn1 = 32'd7984
; 
32'd173744: dataIn1 = 32'd7985
; 
32'd173745: dataIn1 = 32'd7989
; 
32'd173746: dataIn1 = 32'd5194
; 
32'd173747: dataIn1 = 32'd6354
; 
32'd173748: dataIn1 = 32'd7910
; 
32'd173749: dataIn1 = 32'd7981
; 
32'd173750: dataIn1 = 32'd7986
; 
32'd173751: dataIn1 = 32'd7987
; 
32'd173752: dataIn1 = 32'd7993
; 
32'd173753: dataIn1 = 32'd5194
; 
32'd173754: dataIn1 = 32'd6353
; 
32'd173755: dataIn1 = 32'd7903
; 
32'd173756: dataIn1 = 32'd7981
; 
32'd173757: dataIn1 = 32'd7986
; 
32'd173758: dataIn1 = 32'd7987
; 
32'd173759: dataIn1 = 32'd7990
; 
32'd173760: dataIn1 = 32'd6328
; 
32'd173761: dataIn1 = 32'd6343
; 
32'd173762: dataIn1 = 32'd7902
; 
32'd173763: dataIn1 = 32'd7935
; 
32'd173764: dataIn1 = 32'd7988
; 
32'd173765: dataIn1 = 32'd7989
; 
32'd173766: dataIn1 = 32'd7990
; 
32'd173767: dataIn1 = 32'd6343
; 
32'd173768: dataIn1 = 32'd6353
; 
32'd173769: dataIn1 = 32'd7937
; 
32'd173770: dataIn1 = 32'd7985
; 
32'd173771: dataIn1 = 32'd7988
; 
32'd173772: dataIn1 = 32'd7989
; 
32'd173773: dataIn1 = 32'd7990
; 
32'd173774: dataIn1 = 32'd6328
; 
32'd173775: dataIn1 = 32'd6353
; 
32'd173776: dataIn1 = 32'd7903
; 
32'd173777: dataIn1 = 32'd7987
; 
32'd173778: dataIn1 = 32'd7988
; 
32'd173779: dataIn1 = 32'd7989
; 
32'd173780: dataIn1 = 32'd7990
; 
32'd173781: dataIn1 = 32'd4972
; 
32'd173782: dataIn1 = 32'd6354
; 
32'd173783: dataIn1 = 32'd7983
; 
32'd173784: dataIn1 = 32'd7991
; 
32'd173785: dataIn1 = 32'd7992
; 
32'd173786: dataIn1 = 32'd7993
; 
32'd173787: dataIn1 = 32'd7994
; 
32'd173788: dataIn1 = 32'd4972
; 
32'd173789: dataIn1 = 32'd6329
; 
32'd173790: dataIn1 = 32'd7909
; 
32'd173791: dataIn1 = 32'd7991
; 
32'd173792: dataIn1 = 32'd7992
; 
32'd173793: dataIn1 = 32'd7993
; 
32'd173794: dataIn1 = 32'd7995
; 
32'd173795: dataIn1 = 32'd6329
; 
32'd173796: dataIn1 = 32'd6354
; 
32'd173797: dataIn1 = 32'd7910
; 
32'd173798: dataIn1 = 32'd7986
; 
32'd173799: dataIn1 = 32'd7991
; 
32'd173800: dataIn1 = 32'd7992
; 
32'd173801: dataIn1 = 32'd7993
; 
32'd173802: dataIn1 = 32'd2655
; 
32'd173803: dataIn1 = 32'd4969
; 
32'd173804: dataIn1 = 32'd4972
; 
32'd173805: dataIn1 = 32'd7983
; 
32'd173806: dataIn1 = 32'd7991
; 
32'd173807: dataIn1 = 32'd7994
; 
32'd173808: dataIn1 = 32'd139
; 
32'd173809: dataIn1 = 32'd4723
; 
32'd173810: dataIn1 = 32'd4972
; 
32'd173811: dataIn1 = 32'd7909
; 
32'd173812: dataIn1 = 32'd7992
; 
32'd173813: dataIn1 = 32'd7995
; 
32'd173814: dataIn1 = 32'd4973
; 
32'd173815: dataIn1 = 32'd6355
; 
32'd173816: dataIn1 = 32'd7982
; 
32'd173817: dataIn1 = 32'd7996
; 
32'd173818: dataIn1 = 32'd7997
; 
32'd173819: dataIn1 = 32'd7998
; 
32'd173820: dataIn1 = 32'd7999
; 
32'd173821: dataIn1 = 32'd6346
; 
32'd173822: dataIn1 = 32'd6355
; 
32'd173823: dataIn1 = 32'd7950
; 
32'd173824: dataIn1 = 32'd7984
; 
32'd173825: dataIn1 = 32'd7996
; 
32'd173826: dataIn1 = 32'd7997
; 
32'd173827: dataIn1 = 32'd7998
; 
32'd173828: dataIn1 = 32'd4973
; 
32'd173829: dataIn1 = 32'd6346
; 
32'd173830: dataIn1 = 32'd7952
; 
32'd173831: dataIn1 = 32'd7996
; 
32'd173832: dataIn1 = 32'd7997
; 
32'd173833: dataIn1 = 32'd7998
; 
32'd173834: dataIn1 = 32'd8000
; 
32'd173835: dataIn1 = 32'd2655
; 
32'd173836: dataIn1 = 32'd4971
; 
32'd173837: dataIn1 = 32'd4973
; 
32'd173838: dataIn1 = 32'd7982
; 
32'd173839: dataIn1 = 32'd7996
; 
32'd173840: dataIn1 = 32'd7999
; 
32'd173841: dataIn1 = 32'd1111
; 
32'd173842: dataIn1 = 32'd4968
; 
32'd173843: dataIn1 = 32'd4973
; 
32'd173844: dataIn1 = 32'd7952
; 
32'd173845: dataIn1 = 32'd7998
; 
32'd173846: dataIn1 = 32'd8000
; 
32'd173847: dataIn1 = 32'd6357
; 
32'd173848: dataIn1 = 32'd6358
; 
32'd173849: dataIn1 = 32'd8001
; 
32'd173850: dataIn1 = 32'd8002
; 
32'd173851: dataIn1 = 32'd8003
; 
32'd173852: dataIn1 = 32'd8004
; 
32'd173853: dataIn1 = 32'd8005
; 
32'd173854: dataIn1 = 32'd6356
; 
32'd173855: dataIn1 = 32'd6358
; 
32'd173856: dataIn1 = 32'd8001
; 
32'd173857: dataIn1 = 32'd8002
; 
32'd173858: dataIn1 = 32'd8003
; 
32'd173859: dataIn1 = 32'd8006
; 
32'd173860: dataIn1 = 32'd8007
; 
32'd173861: dataIn1 = 32'd6356
; 
32'd173862: dataIn1 = 32'd6357
; 
32'd173863: dataIn1 = 32'd8001
; 
32'd173864: dataIn1 = 32'd8002
; 
32'd173865: dataIn1 = 32'd8003
; 
32'd173866: dataIn1 = 32'd8008
; 
32'd173867: dataIn1 = 32'd8009
; 
32'd173868: dataIn1 = 32'd5201
; 
32'd173869: dataIn1 = 32'd6358
; 
32'd173870: dataIn1 = 32'd6360
; 
32'd173871: dataIn1 = 32'd8001
; 
32'd173872: dataIn1 = 32'd8004
; 
32'd173873: dataIn1 = 32'd8005
; 
32'd173874: dataIn1 = 32'd5201
; 
32'd173875: dataIn1 = 32'd6357
; 
32'd173876: dataIn1 = 32'd8001
; 
32'd173877: dataIn1 = 32'd8004
; 
32'd173878: dataIn1 = 32'd8005
; 
32'd173879: dataIn1 = 32'd8013
; 
32'd173880: dataIn1 = 32'd8016
; 
32'd173881: dataIn1 = 32'd5196
; 
32'd173882: dataIn1 = 32'd6336
; 
32'd173883: dataIn1 = 32'd6358
; 
32'd173884: dataIn1 = 32'd8002
; 
32'd173885: dataIn1 = 32'd8006
; 
32'd173886: dataIn1 = 32'd8007
; 
32'd173887: dataIn1 = 32'd5196
; 
32'd173888: dataIn1 = 32'd6356
; 
32'd173889: dataIn1 = 32'd7920
; 
32'd173890: dataIn1 = 32'd8002
; 
32'd173891: dataIn1 = 32'd8006
; 
32'd173892: dataIn1 = 32'd8007
; 
32'd173893: dataIn1 = 32'd8011
; 
32'd173894: dataIn1 = 32'd5199
; 
32'd173895: dataIn1 = 32'd6357
; 
32'd173896: dataIn1 = 32'd7945
; 
32'd173897: dataIn1 = 32'd8003
; 
32'd173898: dataIn1 = 32'd8008
; 
32'd173899: dataIn1 = 32'd8009
; 
32'd173900: dataIn1 = 32'd8015
; 
32'd173901: dataIn1 = 32'd5199
; 
32'd173902: dataIn1 = 32'd6356
; 
32'd173903: dataIn1 = 32'd7938
; 
32'd173904: dataIn1 = 32'd8003
; 
32'd173905: dataIn1 = 32'd8008
; 
32'd173906: dataIn1 = 32'd8009
; 
32'd173907: dataIn1 = 32'd8012
; 
32'd173908: dataIn1 = 32'd6333
; 
32'd173909: dataIn1 = 32'd6342
; 
32'd173910: dataIn1 = 32'd7919
; 
32'd173911: dataIn1 = 32'd7936
; 
32'd173912: dataIn1 = 32'd8010
; 
32'd173913: dataIn1 = 32'd8011
; 
32'd173914: dataIn1 = 32'd8012
; 
32'd173915: dataIn1 = 32'd6333
; 
32'd173916: dataIn1 = 32'd6356
; 
32'd173917: dataIn1 = 32'd7920
; 
32'd173918: dataIn1 = 32'd8007
; 
32'd173919: dataIn1 = 32'd8010
; 
32'd173920: dataIn1 = 32'd8011
; 
32'd173921: dataIn1 = 32'd8012
; 
32'd173922: dataIn1 = 32'd6342
; 
32'd173923: dataIn1 = 32'd6356
; 
32'd173924: dataIn1 = 32'd7938
; 
32'd173925: dataIn1 = 32'd8009
; 
32'd173926: dataIn1 = 32'd8010
; 
32'd173927: dataIn1 = 32'd8011
; 
32'd173928: dataIn1 = 32'd8012
; 
32'd173929: dataIn1 = 32'd6357
; 
32'd173930: dataIn1 = 32'd6359
; 
32'd173931: dataIn1 = 32'd8005
; 
32'd173932: dataIn1 = 32'd8013
; 
32'd173933: dataIn1 = 32'd8014
; 
32'd173934: dataIn1 = 32'd8015
; 
32'd173935: dataIn1 = 32'd8016
; 
32'd173936: dataIn1 = 32'd6344
; 
32'd173937: dataIn1 = 32'd6359
; 
32'd173938: dataIn1 = 32'd7944
; 
32'd173939: dataIn1 = 32'd8013
; 
32'd173940: dataIn1 = 32'd8014
; 
32'd173941: dataIn1 = 32'd8015
; 
32'd173942: dataIn1 = 32'd8017
; 
32'd173943: dataIn1 = 32'd6344
; 
32'd173944: dataIn1 = 32'd6357
; 
32'd173945: dataIn1 = 32'd7945
; 
32'd173946: dataIn1 = 32'd8008
; 
32'd173947: dataIn1 = 32'd8013
; 
32'd173948: dataIn1 = 32'd8014
; 
32'd173949: dataIn1 = 32'd8015
; 
32'd173950: dataIn1 = 32'd5201
; 
32'd173951: dataIn1 = 32'd6359
; 
32'd173952: dataIn1 = 32'd8005
; 
32'd173953: dataIn1 = 32'd8013
; 
32'd173954: dataIn1 = 32'd8016
; 
32'd173955: dataIn1 = 32'd9069
; 
32'd173956: dataIn1 = 32'd9072
; 
32'd173957: dataIn1 = 32'd2717
; 
32'd173958: dataIn1 = 32'd6359
; 
32'd173959: dataIn1 = 32'd7944
; 
32'd173960: dataIn1 = 32'd8014
; 
32'd173961: dataIn1 = 32'd8017
; 
32'd173962: dataIn1 = 32'd9050
; 
32'd173963: dataIn1 = 32'd9071
; 
32'd173964: dataIn1 = 32'd6362
; 
32'd173965: dataIn1 = 32'd6363
; 
32'd173966: dataIn1 = 32'd8018
; 
32'd173967: dataIn1 = 32'd8019
; 
32'd173968: dataIn1 = 32'd8020
; 
32'd173969: dataIn1 = 32'd8021
; 
32'd173970: dataIn1 = 32'd8022
; 
32'd173971: dataIn1 = 32'd6361
; 
32'd173972: dataIn1 = 32'd6363
; 
32'd173973: dataIn1 = 32'd8018
; 
32'd173974: dataIn1 = 32'd8019
; 
32'd173975: dataIn1 = 32'd8020
; 
32'd173976: dataIn1 = 32'd8023
; 
32'd173977: dataIn1 = 32'd8024
; 
32'd173978: dataIn1 = 32'd6361
; 
32'd173979: dataIn1 = 32'd6362
; 
32'd173980: dataIn1 = 32'd8018
; 
32'd173981: dataIn1 = 32'd8019
; 
32'd173982: dataIn1 = 32'd8020
; 
32'd173983: dataIn1 = 32'd8025
; 
32'd173984: dataIn1 = 32'd8026
; 
32'd173985: dataIn1 = 32'd5202
; 
32'd173986: dataIn1 = 32'd6363
; 
32'd173987: dataIn1 = 32'd8018
; 
32'd173988: dataIn1 = 32'd8021
; 
32'd173989: dataIn1 = 32'd8022
; 
32'd173990: dataIn1 = 32'd8041
; 
32'd173991: dataIn1 = 32'd8044
; 
32'd173992: dataIn1 = 32'd5202
; 
32'd173993: dataIn1 = 32'd6362
; 
32'd173994: dataIn1 = 32'd8018
; 
32'd173995: dataIn1 = 32'd8021
; 
32'd173996: dataIn1 = 32'd8022
; 
32'd173997: dataIn1 = 32'd8034
; 
32'd173998: dataIn1 = 32'd8037
; 
32'd173999: dataIn1 = 32'd5203
; 
32'd174000: dataIn1 = 32'd6363
; 
32'd174001: dataIn1 = 32'd8019
; 
32'd174002: dataIn1 = 32'd8023
; 
32'd174003: dataIn1 = 32'd8024
; 
32'd174004: dataIn1 = 32'd8042
; 
32'd174005: dataIn1 = 32'd8045
; 
32'd174006: dataIn1 = 32'd5203
; 
32'd174007: dataIn1 = 32'd6361
; 
32'd174008: dataIn1 = 32'd8019
; 
32'd174009: dataIn1 = 32'd8023
; 
32'd174010: dataIn1 = 32'd8024
; 
32'd174011: dataIn1 = 32'd8028
; 
32'd174012: dataIn1 = 32'd8032
; 
32'd174013: dataIn1 = 32'd5204
; 
32'd174014: dataIn1 = 32'd6362
; 
32'd174015: dataIn1 = 32'd8020
; 
32'd174016: dataIn1 = 32'd8025
; 
32'd174017: dataIn1 = 32'd8026
; 
32'd174018: dataIn1 = 32'd8036
; 
32'd174019: dataIn1 = 32'd8040
; 
32'd174020: dataIn1 = 32'd5204
; 
32'd174021: dataIn1 = 32'd6361
; 
32'd174022: dataIn1 = 32'd8020
; 
32'd174023: dataIn1 = 32'd8025
; 
32'd174024: dataIn1 = 32'd8026
; 
32'd174025: dataIn1 = 32'd8029
; 
32'd174026: dataIn1 = 32'd8033
; 
32'd174027: dataIn1 = 32'd6364
; 
32'd174028: dataIn1 = 32'd6365
; 
32'd174029: dataIn1 = 32'd8027
; 
32'd174030: dataIn1 = 32'd8028
; 
32'd174031: dataIn1 = 32'd8029
; 
32'd174032: dataIn1 = 32'd8030
; 
32'd174033: dataIn1 = 32'd8031
; 
32'd174034: dataIn1 = 32'd6361
; 
32'd174035: dataIn1 = 32'd6365
; 
32'd174036: dataIn1 = 32'd8024
; 
32'd174037: dataIn1 = 32'd8027
; 
32'd174038: dataIn1 = 32'd8028
; 
32'd174039: dataIn1 = 32'd8029
; 
32'd174040: dataIn1 = 32'd8032
; 
32'd174041: dataIn1 = 32'd6361
; 
32'd174042: dataIn1 = 32'd6364
; 
32'd174043: dataIn1 = 32'd8026
; 
32'd174044: dataIn1 = 32'd8027
; 
32'd174045: dataIn1 = 32'd8028
; 
32'd174046: dataIn1 = 32'd8029
; 
32'd174047: dataIn1 = 32'd8033
; 
32'd174048: dataIn1 = 32'd1112
; 
32'd174049: dataIn1 = 32'd6365
; 
32'd174050: dataIn1 = 32'd8027
; 
32'd174051: dataIn1 = 32'd8030
; 
32'd174052: dataIn1 = 32'd8031
; 
32'd174053: dataIn1 = 32'd8074
; 
32'd174054: dataIn1 = 32'd8077
; 
32'd174055: dataIn1 = 32'd1112
; 
32'd174056: dataIn1 = 32'd6364
; 
32'd174057: dataIn1 = 32'd8027
; 
32'd174058: dataIn1 = 32'd8030
; 
32'd174059: dataIn1 = 32'd8031
; 
32'd174060: dataIn1 = 32'd8096
; 
32'd174061: dataIn1 = 32'd8099
; 
32'd174062: dataIn1 = 32'd5203
; 
32'd174063: dataIn1 = 32'd6365
; 
32'd174064: dataIn1 = 32'd8024
; 
32'd174065: dataIn1 = 32'd8028
; 
32'd174066: dataIn1 = 32'd8032
; 
32'd174067: dataIn1 = 32'd8071
; 
32'd174068: dataIn1 = 32'd8075
; 
32'd174069: dataIn1 = 32'd5204
; 
32'd174070: dataIn1 = 32'd6364
; 
32'd174071: dataIn1 = 32'd8026
; 
32'd174072: dataIn1 = 32'd8029
; 
32'd174073: dataIn1 = 32'd8033
; 
32'd174074: dataIn1 = 32'd8095
; 
32'd174075: dataIn1 = 32'd8098
; 
32'd174076: dataIn1 = 32'd6362
; 
32'd174077: dataIn1 = 32'd6367
; 
32'd174078: dataIn1 = 32'd8022
; 
32'd174079: dataIn1 = 32'd8034
; 
32'd174080: dataIn1 = 32'd8035
; 
32'd174081: dataIn1 = 32'd8036
; 
32'd174082: dataIn1 = 32'd8037
; 
32'd174083: dataIn1 = 32'd6366
; 
32'd174084: dataIn1 = 32'd6367
; 
32'd174085: dataIn1 = 32'd8034
; 
32'd174086: dataIn1 = 32'd8035
; 
32'd174087: dataIn1 = 32'd8036
; 
32'd174088: dataIn1 = 32'd8038
; 
32'd174089: dataIn1 = 32'd8039
; 
32'd174090: dataIn1 = 32'd6362
; 
32'd174091: dataIn1 = 32'd6366
; 
32'd174092: dataIn1 = 32'd8025
; 
32'd174093: dataIn1 = 32'd8034
; 
32'd174094: dataIn1 = 32'd8035
; 
32'd174095: dataIn1 = 32'd8036
; 
32'd174096: dataIn1 = 32'd8040
; 
32'd174097: dataIn1 = 32'd5202
; 
32'd174098: dataIn1 = 32'd6367
; 
32'd174099: dataIn1 = 32'd8022
; 
32'd174100: dataIn1 = 32'd8034
; 
32'd174101: dataIn1 = 32'd8037
; 
32'd174102: dataIn1 = 32'd8052
; 
32'd174103: dataIn1 = 32'd8057
; 
32'd174104: dataIn1 = 32'd2718
; 
32'd174105: dataIn1 = 32'd6367
; 
32'd174106: dataIn1 = 32'd8035
; 
32'd174107: dataIn1 = 32'd8038
; 
32'd174108: dataIn1 = 32'd8039
; 
32'd174109: dataIn1 = 32'd8058
; 
32'd174110: dataIn1 = 32'd8060
; 
32'd174111: dataIn1 = 32'd2718
; 
32'd174112: dataIn1 = 32'd6366
; 
32'd174113: dataIn1 = 32'd8035
; 
32'd174114: dataIn1 = 32'd8038
; 
32'd174115: dataIn1 = 32'd8039
; 
32'd174116: dataIn1 = 32'd8102
; 
32'd174117: dataIn1 = 32'd8105
; 
32'd174118: dataIn1 = 32'd5204
; 
32'd174119: dataIn1 = 32'd6366
; 
32'd174120: dataIn1 = 32'd8025
; 
32'd174121: dataIn1 = 32'd8036
; 
32'd174122: dataIn1 = 32'd8040
; 
32'd174123: dataIn1 = 32'd8094
; 
32'd174124: dataIn1 = 32'd8103
; 
32'd174125: dataIn1 = 32'd6363
; 
32'd174126: dataIn1 = 32'd6369
; 
32'd174127: dataIn1 = 32'd8021
; 
32'd174128: dataIn1 = 32'd8041
; 
32'd174129: dataIn1 = 32'd8042
; 
32'd174130: dataIn1 = 32'd8043
; 
32'd174131: dataIn1 = 32'd8044
; 
32'd174132: dataIn1 = 32'd6363
; 
32'd174133: dataIn1 = 32'd6368
; 
32'd174134: dataIn1 = 32'd8023
; 
32'd174135: dataIn1 = 32'd8041
; 
32'd174136: dataIn1 = 32'd8042
; 
32'd174137: dataIn1 = 32'd8043
; 
32'd174138: dataIn1 = 32'd8045
; 
32'd174139: dataIn1 = 32'd6368
; 
32'd174140: dataIn1 = 32'd6369
; 
32'd174141: dataIn1 = 32'd8041
; 
32'd174142: dataIn1 = 32'd8042
; 
32'd174143: dataIn1 = 32'd8043
; 
32'd174144: dataIn1 = 32'd8046
; 
32'd174145: dataIn1 = 32'd8047
; 
32'd174146: dataIn1 = 32'd5202
; 
32'd174147: dataIn1 = 32'd6369
; 
32'd174148: dataIn1 = 32'd8021
; 
32'd174149: dataIn1 = 32'd8041
; 
32'd174150: dataIn1 = 32'd8044
; 
32'd174151: dataIn1 = 32'd8051
; 
32'd174152: dataIn1 = 32'd8062
; 
32'd174153: dataIn1 = 32'd5203
; 
32'd174154: dataIn1 = 32'd6368
; 
32'd174155: dataIn1 = 32'd8023
; 
32'd174156: dataIn1 = 32'd8042
; 
32'd174157: dataIn1 = 32'd8045
; 
32'd174158: dataIn1 = 32'd8070
; 
32'd174159: dataIn1 = 32'd8085
; 
32'd174160: dataIn1 = 32'd2716
; 
32'd174161: dataIn1 = 32'd6369
; 
32'd174162: dataIn1 = 32'd7889
; 
32'd174163: dataIn1 = 32'd8043
; 
32'd174164: dataIn1 = 32'd8046
; 
32'd174165: dataIn1 = 32'd8047
; 
32'd174166: dataIn1 = 32'd8064
; 
32'd174167: dataIn1 = 32'd2716
; 
32'd174168: dataIn1 = 32'd6368
; 
32'd174169: dataIn1 = 32'd7915
; 
32'd174170: dataIn1 = 32'd8043
; 
32'd174171: dataIn1 = 32'd8046
; 
32'd174172: dataIn1 = 32'd8047
; 
32'd174173: dataIn1 = 32'd8086
; 
32'd174174: dataIn1 = 32'd6371
; 
32'd174175: dataIn1 = 32'd6372
; 
32'd174176: dataIn1 = 32'd8048
; 
32'd174177: dataIn1 = 32'd8049
; 
32'd174178: dataIn1 = 32'd8050
; 
32'd174179: dataIn1 = 32'd8051
; 
32'd174180: dataIn1 = 32'd8052
; 
32'd174181: dataIn1 = 32'd6370
; 
32'd174182: dataIn1 = 32'd6372
; 
32'd174183: dataIn1 = 32'd8048
; 
32'd174184: dataIn1 = 32'd8049
; 
32'd174185: dataIn1 = 32'd8050
; 
32'd174186: dataIn1 = 32'd8053
; 
32'd174187: dataIn1 = 32'd8054
; 
32'd174188: dataIn1 = 32'd6370
; 
32'd174189: dataIn1 = 32'd6371
; 
32'd174190: dataIn1 = 32'd8048
; 
32'd174191: dataIn1 = 32'd8049
; 
32'd174192: dataIn1 = 32'd8050
; 
32'd174193: dataIn1 = 32'd8055
; 
32'd174194: dataIn1 = 32'd8056
; 
32'd174195: dataIn1 = 32'd5202
; 
32'd174196: dataIn1 = 32'd6372
; 
32'd174197: dataIn1 = 32'd8044
; 
32'd174198: dataIn1 = 32'd8048
; 
32'd174199: dataIn1 = 32'd8051
; 
32'd174200: dataIn1 = 32'd8052
; 
32'd174201: dataIn1 = 32'd8062
; 
32'd174202: dataIn1 = 32'd5202
; 
32'd174203: dataIn1 = 32'd6371
; 
32'd174204: dataIn1 = 32'd8037
; 
32'd174205: dataIn1 = 32'd8048
; 
32'd174206: dataIn1 = 32'd8051
; 
32'd174207: dataIn1 = 32'd8052
; 
32'd174208: dataIn1 = 32'd8057
; 
32'd174209: dataIn1 = 32'd5191
; 
32'd174210: dataIn1 = 32'd6372
; 
32'd174211: dataIn1 = 32'd7888
; 
32'd174212: dataIn1 = 32'd8049
; 
32'd174213: dataIn1 = 32'd8053
; 
32'd174214: dataIn1 = 32'd8054
; 
32'd174215: dataIn1 = 32'd8063
; 
32'd174216: dataIn1 = 32'd5191
; 
32'd174217: dataIn1 = 32'd6320
; 
32'd174218: dataIn1 = 32'd6370
; 
32'd174219: dataIn1 = 32'd8049
; 
32'd174220: dataIn1 = 32'd8053
; 
32'd174221: dataIn1 = 32'd8054
; 
32'd174222: dataIn1 = 32'd5205
; 
32'd174223: dataIn1 = 32'd6371
; 
32'd174224: dataIn1 = 32'd8050
; 
32'd174225: dataIn1 = 32'd8055
; 
32'd174226: dataIn1 = 32'd8056
; 
32'd174227: dataIn1 = 32'd8059
; 
32'd174228: dataIn1 = 32'd8061
; 
32'd174229: dataIn1 = 32'd5205
; 
32'd174230: dataIn1 = 32'd6370
; 
32'd174231: dataIn1 = 32'd6373
; 
32'd174232: dataIn1 = 32'd8050
; 
32'd174233: dataIn1 = 32'd8055
; 
32'd174234: dataIn1 = 32'd8056
; 
32'd174235: dataIn1 = 32'd6367
; 
32'd174236: dataIn1 = 32'd6371
; 
32'd174237: dataIn1 = 32'd8037
; 
32'd174238: dataIn1 = 32'd8052
; 
32'd174239: dataIn1 = 32'd8057
; 
32'd174240: dataIn1 = 32'd8058
; 
32'd174241: dataIn1 = 32'd8059
; 
32'd174242: dataIn1 = 32'd6367
; 
32'd174243: dataIn1 = 32'd6374
; 
32'd174244: dataIn1 = 32'd8038
; 
32'd174245: dataIn1 = 32'd8057
; 
32'd174246: dataIn1 = 32'd8058
; 
32'd174247: dataIn1 = 32'd8059
; 
32'd174248: dataIn1 = 32'd8060
; 
32'd174249: dataIn1 = 32'd6371
; 
32'd174250: dataIn1 = 32'd6374
; 
32'd174251: dataIn1 = 32'd8055
; 
32'd174252: dataIn1 = 32'd8057
; 
32'd174253: dataIn1 = 32'd8058
; 
32'd174254: dataIn1 = 32'd8059
; 
32'd174255: dataIn1 = 32'd8061
; 
32'd174256: dataIn1 = 32'd2718
; 
32'd174257: dataIn1 = 32'd6374
; 
32'd174258: dataIn1 = 32'd8038
; 
32'd174259: dataIn1 = 32'd8058
; 
32'd174260: dataIn1 = 32'd8060
; 
32'd174261: dataIn1 = 32'd9093
; 
32'd174262: dataIn1 = 32'd9126
; 
32'd174263: dataIn1 = 32'd5205
; 
32'd174264: dataIn1 = 32'd6374
; 
32'd174265: dataIn1 = 32'd8055
; 
32'd174266: dataIn1 = 32'd8059
; 
32'd174267: dataIn1 = 32'd8061
; 
32'd174268: dataIn1 = 32'd9125
; 
32'd174269: dataIn1 = 32'd9128
; 
32'd174270: dataIn1 = 32'd6369
; 
32'd174271: dataIn1 = 32'd6372
; 
32'd174272: dataIn1 = 32'd8044
; 
32'd174273: dataIn1 = 32'd8051
; 
32'd174274: dataIn1 = 32'd8062
; 
32'd174275: dataIn1 = 32'd8063
; 
32'd174276: dataIn1 = 32'd8064
; 
32'd174277: dataIn1 = 32'd6323
; 
32'd174278: dataIn1 = 32'd6372
; 
32'd174279: dataIn1 = 32'd7888
; 
32'd174280: dataIn1 = 32'd8053
; 
32'd174281: dataIn1 = 32'd8062
; 
32'd174282: dataIn1 = 32'd8063
; 
32'd174283: dataIn1 = 32'd8064
; 
32'd174284: dataIn1 = 32'd6323
; 
32'd174285: dataIn1 = 32'd6369
; 
32'd174286: dataIn1 = 32'd7889
; 
32'd174287: dataIn1 = 32'd8046
; 
32'd174288: dataIn1 = 32'd8062
; 
32'd174289: dataIn1 = 32'd8063
; 
32'd174290: dataIn1 = 32'd8064
; 
32'd174291: dataIn1 = 32'd6376
; 
32'd174292: dataIn1 = 32'd6377
; 
32'd174293: dataIn1 = 32'd8065
; 
32'd174294: dataIn1 = 32'd8066
; 
32'd174295: dataIn1 = 32'd8067
; 
32'd174296: dataIn1 = 32'd8068
; 
32'd174297: dataIn1 = 32'd8069
; 
32'd174298: dataIn1 = 32'd6375
; 
32'd174299: dataIn1 = 32'd6377
; 
32'd174300: dataIn1 = 32'd8065
; 
32'd174301: dataIn1 = 32'd8066
; 
32'd174302: dataIn1 = 32'd8067
; 
32'd174303: dataIn1 = 32'd8070
; 
32'd174304: dataIn1 = 32'd8071
; 
32'd174305: dataIn1 = 32'd6375
; 
32'd174306: dataIn1 = 32'd6376
; 
32'd174307: dataIn1 = 32'd8065
; 
32'd174308: dataIn1 = 32'd8066
; 
32'd174309: dataIn1 = 32'd8067
; 
32'd174310: dataIn1 = 32'd8072
; 
32'd174311: dataIn1 = 32'd8073
; 
32'd174312: dataIn1 = 32'd5193
; 
32'd174313: dataIn1 = 32'd6377
; 
32'd174314: dataIn1 = 32'd7914
; 
32'd174315: dataIn1 = 32'd8065
; 
32'd174316: dataIn1 = 32'd8068
; 
32'd174317: dataIn1 = 32'd8069
; 
32'd174318: dataIn1 = 32'd8084
; 
32'd174319: dataIn1 = 32'd5193
; 
32'd174320: dataIn1 = 32'd6376
; 
32'd174321: dataIn1 = 32'd7907
; 
32'd174322: dataIn1 = 32'd8065
; 
32'd174323: dataIn1 = 32'd8068
; 
32'd174324: dataIn1 = 32'd8069
; 
32'd174325: dataIn1 = 32'd8079
; 
32'd174326: dataIn1 = 32'd5203
; 
32'd174327: dataIn1 = 32'd6377
; 
32'd174328: dataIn1 = 32'd8045
; 
32'd174329: dataIn1 = 32'd8066
; 
32'd174330: dataIn1 = 32'd8070
; 
32'd174331: dataIn1 = 32'd8071
; 
32'd174332: dataIn1 = 32'd8085
; 
32'd174333: dataIn1 = 32'd5203
; 
32'd174334: dataIn1 = 32'd6375
; 
32'd174335: dataIn1 = 32'd8032
; 
32'd174336: dataIn1 = 32'd8066
; 
32'd174337: dataIn1 = 32'd8070
; 
32'd174338: dataIn1 = 32'd8071
; 
32'd174339: dataIn1 = 32'd8075
; 
32'd174340: dataIn1 = 32'd2660
; 
32'd174341: dataIn1 = 32'd6376
; 
32'd174342: dataIn1 = 32'd8067
; 
32'd174343: dataIn1 = 32'd8072
; 
32'd174344: dataIn1 = 32'd8073
; 
32'd174345: dataIn1 = 32'd8081
; 
32'd174346: dataIn1 = 32'd8083
; 
32'd174347: dataIn1 = 32'd2660
; 
32'd174348: dataIn1 = 32'd6375
; 
32'd174349: dataIn1 = 32'd8067
; 
32'd174350: dataIn1 = 32'd8072
; 
32'd174351: dataIn1 = 32'd8073
; 
32'd174352: dataIn1 = 32'd8076
; 
32'd174353: dataIn1 = 32'd8078
; 
32'd174354: dataIn1 = 32'd4992
; 
32'd174355: dataIn1 = 32'd6365
; 
32'd174356: dataIn1 = 32'd8030
; 
32'd174357: dataIn1 = 32'd8074
; 
32'd174358: dataIn1 = 32'd8075
; 
32'd174359: dataIn1 = 32'd8076
; 
32'd174360: dataIn1 = 32'd8077
; 
32'd174361: dataIn1 = 32'd6365
; 
32'd174362: dataIn1 = 32'd6375
; 
32'd174363: dataIn1 = 32'd8032
; 
32'd174364: dataIn1 = 32'd8071
; 
32'd174365: dataIn1 = 32'd8074
; 
32'd174366: dataIn1 = 32'd8075
; 
32'd174367: dataIn1 = 32'd8076
; 
32'd174368: dataIn1 = 32'd4992
; 
32'd174369: dataIn1 = 32'd6375
; 
32'd174370: dataIn1 = 32'd8073
; 
32'd174371: dataIn1 = 32'd8074
; 
32'd174372: dataIn1 = 32'd8075
; 
32'd174373: dataIn1 = 32'd8076
; 
32'd174374: dataIn1 = 32'd8078
; 
32'd174375: dataIn1 = 32'd1112
; 
32'd174376: dataIn1 = 32'd4985
; 
32'd174377: dataIn1 = 32'd4992
; 
32'd174378: dataIn1 = 32'd8030
; 
32'd174379: dataIn1 = 32'd8074
; 
32'd174380: dataIn1 = 32'd8077
; 
32'd174381: dataIn1 = 32'd2660
; 
32'd174382: dataIn1 = 32'd4989
; 
32'd174383: dataIn1 = 32'd4992
; 
32'd174384: dataIn1 = 32'd8073
; 
32'd174385: dataIn1 = 32'd8076
; 
32'd174386: dataIn1 = 32'd8078
; 
32'd174387: dataIn1 = 32'd6330
; 
32'd174388: dataIn1 = 32'd6376
; 
32'd174389: dataIn1 = 32'd7907
; 
32'd174390: dataIn1 = 32'd8069
; 
32'd174391: dataIn1 = 32'd8079
; 
32'd174392: dataIn1 = 32'd8080
; 
32'd174393: dataIn1 = 32'd8081
; 
32'd174394: dataIn1 = 32'd4991
; 
32'd174395: dataIn1 = 32'd6330
; 
32'd174396: dataIn1 = 32'd7908
; 
32'd174397: dataIn1 = 32'd8079
; 
32'd174398: dataIn1 = 32'd8080
; 
32'd174399: dataIn1 = 32'd8081
; 
32'd174400: dataIn1 = 32'd8082
; 
32'd174401: dataIn1 = 32'd4991
; 
32'd174402: dataIn1 = 32'd6376
; 
32'd174403: dataIn1 = 32'd8072
; 
32'd174404: dataIn1 = 32'd8079
; 
32'd174405: dataIn1 = 32'd8080
; 
32'd174406: dataIn1 = 32'd8081
; 
32'd174407: dataIn1 = 32'd8083
; 
32'd174408: dataIn1 = 32'd139
; 
32'd174409: dataIn1 = 32'd4724
; 
32'd174410: dataIn1 = 32'd4991
; 
32'd174411: dataIn1 = 32'd7908
; 
32'd174412: dataIn1 = 32'd8080
; 
32'd174413: dataIn1 = 32'd8082
; 
32'd174414: dataIn1 = 32'd2660
; 
32'd174415: dataIn1 = 32'd4988
; 
32'd174416: dataIn1 = 32'd4991
; 
32'd174417: dataIn1 = 32'd8072
; 
32'd174418: dataIn1 = 32'd8081
; 
32'd174419: dataIn1 = 32'd8083
; 
32'd174420: dataIn1 = 32'd6331
; 
32'd174421: dataIn1 = 32'd6377
; 
32'd174422: dataIn1 = 32'd7914
; 
32'd174423: dataIn1 = 32'd8068
; 
32'd174424: dataIn1 = 32'd8084
; 
32'd174425: dataIn1 = 32'd8085
; 
32'd174426: dataIn1 = 32'd8086
; 
32'd174427: dataIn1 = 32'd6368
; 
32'd174428: dataIn1 = 32'd6377
; 
32'd174429: dataIn1 = 32'd8045
; 
32'd174430: dataIn1 = 32'd8070
; 
32'd174431: dataIn1 = 32'd8084
; 
32'd174432: dataIn1 = 32'd8085
; 
32'd174433: dataIn1 = 32'd8086
; 
32'd174434: dataIn1 = 32'd6331
; 
32'd174435: dataIn1 = 32'd6368
; 
32'd174436: dataIn1 = 32'd7915
; 
32'd174437: dataIn1 = 32'd8047
; 
32'd174438: dataIn1 = 32'd8084
; 
32'd174439: dataIn1 = 32'd8085
; 
32'd174440: dataIn1 = 32'd8086
; 
32'd174441: dataIn1 = 32'd6379
; 
32'd174442: dataIn1 = 32'd6380
; 
32'd174443: dataIn1 = 32'd8087
; 
32'd174444: dataIn1 = 32'd8088
; 
32'd174445: dataIn1 = 32'd8089
; 
32'd174446: dataIn1 = 32'd8090
; 
32'd174447: dataIn1 = 32'd8091
; 
32'd174448: dataIn1 = 32'd6378
; 
32'd174449: dataIn1 = 32'd6380
; 
32'd174450: dataIn1 = 32'd8087
; 
32'd174451: dataIn1 = 32'd8088
; 
32'd174452: dataIn1 = 32'd8089
; 
32'd174453: dataIn1 = 32'd8092
; 
32'd174454: dataIn1 = 32'd8093
; 
32'd174455: dataIn1 = 32'd6378
; 
32'd174456: dataIn1 = 32'd6379
; 
32'd174457: dataIn1 = 32'd8087
; 
32'd174458: dataIn1 = 32'd8088
; 
32'd174459: dataIn1 = 32'd8089
; 
32'd174460: dataIn1 = 32'd8094
; 
32'd174461: dataIn1 = 32'd8095
; 
32'd174462: dataIn1 = 32'd5206
; 
32'd174463: dataIn1 = 32'd6380
; 
32'd174464: dataIn1 = 32'd8087
; 
32'd174465: dataIn1 = 32'd8090
; 
32'd174466: dataIn1 = 32'd8091
; 
32'd174467: dataIn1 = 32'd8106
; 
32'd174468: dataIn1 = 32'd8109
; 
32'd174469: dataIn1 = 32'd5206
; 
32'd174470: dataIn1 = 32'd6379
; 
32'd174471: dataIn1 = 32'd8087
; 
32'd174472: dataIn1 = 32'd8090
; 
32'd174473: dataIn1 = 32'd8091
; 
32'd174474: dataIn1 = 32'd8101
; 
32'd174475: dataIn1 = 32'd8104
; 
32'd174476: dataIn1 = 32'd2661
; 
32'd174477: dataIn1 = 32'd6380
; 
32'd174478: dataIn1 = 32'd8088
; 
32'd174479: dataIn1 = 32'd8092
; 
32'd174480: dataIn1 = 32'd8093
; 
32'd174481: dataIn1 = 32'd8107
; 
32'd174482: dataIn1 = 32'd8110
; 
32'd174483: dataIn1 = 32'd2661
; 
32'd174484: dataIn1 = 32'd6378
; 
32'd174485: dataIn1 = 32'd8088
; 
32'd174486: dataIn1 = 32'd8092
; 
32'd174487: dataIn1 = 32'd8093
; 
32'd174488: dataIn1 = 32'd8097
; 
32'd174489: dataIn1 = 32'd8100
; 
32'd174490: dataIn1 = 32'd5204
; 
32'd174491: dataIn1 = 32'd6379
; 
32'd174492: dataIn1 = 32'd8040
; 
32'd174493: dataIn1 = 32'd8089
; 
32'd174494: dataIn1 = 32'd8094
; 
32'd174495: dataIn1 = 32'd8095
; 
32'd174496: dataIn1 = 32'd8103
; 
32'd174497: dataIn1 = 32'd5204
; 
32'd174498: dataIn1 = 32'd6378
; 
32'd174499: dataIn1 = 32'd8033
; 
32'd174500: dataIn1 = 32'd8089
; 
32'd174501: dataIn1 = 32'd8094
; 
32'd174502: dataIn1 = 32'd8095
; 
32'd174503: dataIn1 = 32'd8098
; 
32'd174504: dataIn1 = 32'd4996
; 
32'd174505: dataIn1 = 32'd6364
; 
32'd174506: dataIn1 = 32'd8031
; 
32'd174507: dataIn1 = 32'd8096
; 
32'd174508: dataIn1 = 32'd8097
; 
32'd174509: dataIn1 = 32'd8098
; 
32'd174510: dataIn1 = 32'd8099
; 
32'd174511: dataIn1 = 32'd4996
; 
32'd174512: dataIn1 = 32'd6378
; 
32'd174513: dataIn1 = 32'd8093
; 
32'd174514: dataIn1 = 32'd8096
; 
32'd174515: dataIn1 = 32'd8097
; 
32'd174516: dataIn1 = 32'd8098
; 
32'd174517: dataIn1 = 32'd8100
; 
32'd174518: dataIn1 = 32'd6364
; 
32'd174519: dataIn1 = 32'd6378
; 
32'd174520: dataIn1 = 32'd8033
; 
32'd174521: dataIn1 = 32'd8095
; 
32'd174522: dataIn1 = 32'd8096
; 
32'd174523: dataIn1 = 32'd8097
; 
32'd174524: dataIn1 = 32'd8098
; 
32'd174525: dataIn1 = 32'd1112
; 
32'd174526: dataIn1 = 32'd4984
; 
32'd174527: dataIn1 = 32'd4996
; 
32'd174528: dataIn1 = 32'd8031
; 
32'd174529: dataIn1 = 32'd8096
; 
32'd174530: dataIn1 = 32'd8099
; 
32'd174531: dataIn1 = 32'd2661
; 
32'd174532: dataIn1 = 32'd4994
; 
32'd174533: dataIn1 = 32'd4996
; 
32'd174534: dataIn1 = 32'd8093
; 
32'd174535: dataIn1 = 32'd8097
; 
32'd174536: dataIn1 = 32'd8100
; 
32'd174537: dataIn1 = 32'd6379
; 
32'd174538: dataIn1 = 32'd6381
; 
32'd174539: dataIn1 = 32'd8091
; 
32'd174540: dataIn1 = 32'd8101
; 
32'd174541: dataIn1 = 32'd8102
; 
32'd174542: dataIn1 = 32'd8103
; 
32'd174543: dataIn1 = 32'd8104
; 
32'd174544: dataIn1 = 32'd6366
; 
32'd174545: dataIn1 = 32'd6381
; 
32'd174546: dataIn1 = 32'd8039
; 
32'd174547: dataIn1 = 32'd8101
; 
32'd174548: dataIn1 = 32'd8102
; 
32'd174549: dataIn1 = 32'd8103
; 
32'd174550: dataIn1 = 32'd8105
; 
32'd174551: dataIn1 = 32'd6366
; 
32'd174552: dataIn1 = 32'd6379
; 
32'd174553: dataIn1 = 32'd8040
; 
32'd174554: dataIn1 = 32'd8094
; 
32'd174555: dataIn1 = 32'd8101
; 
32'd174556: dataIn1 = 32'd8102
; 
32'd174557: dataIn1 = 32'd8103
; 
32'd174558: dataIn1 = 32'd5206
; 
32'd174559: dataIn1 = 32'd6381
; 
32'd174560: dataIn1 = 32'd8091
; 
32'd174561: dataIn1 = 32'd8101
; 
32'd174562: dataIn1 = 32'd8104
; 
32'd174563: dataIn1 = 32'd9109
; 
32'd174564: dataIn1 = 32'd9116
; 
32'd174565: dataIn1 = 32'd2718
; 
32'd174566: dataIn1 = 32'd6381
; 
32'd174567: dataIn1 = 32'd8039
; 
32'd174568: dataIn1 = 32'd8102
; 
32'd174569: dataIn1 = 32'd8105
; 
32'd174570: dataIn1 = 32'd9092
; 
32'd174571: dataIn1 = 32'd9115
; 
32'd174572: dataIn1 = 32'd6380
; 
32'd174573: dataIn1 = 32'd6382
; 
32'd174574: dataIn1 = 32'd8090
; 
32'd174575: dataIn1 = 32'd8106
; 
32'd174576: dataIn1 = 32'd8107
; 
32'd174577: dataIn1 = 32'd8108
; 
32'd174578: dataIn1 = 32'd8109
; 
32'd174579: dataIn1 = 32'd4997
; 
32'd174580: dataIn1 = 32'd6380
; 
32'd174581: dataIn1 = 32'd8092
; 
32'd174582: dataIn1 = 32'd8106
; 
32'd174583: dataIn1 = 32'd8107
; 
32'd174584: dataIn1 = 32'd8108
; 
32'd174585: dataIn1 = 32'd8110
; 
32'd174586: dataIn1 = 32'd4997
; 
32'd174587: dataIn1 = 32'd6382
; 
32'd174588: dataIn1 = 32'd8106
; 
32'd174589: dataIn1 = 32'd8107
; 
32'd174590: dataIn1 = 32'd8108
; 
32'd174591: dataIn1 = 32'd8111
; 
32'd174592: dataIn1 = 32'd8112
; 
32'd174593: dataIn1 = 32'd5206
; 
32'd174594: dataIn1 = 32'd6382
; 
32'd174595: dataIn1 = 32'd8090
; 
32'd174596: dataIn1 = 32'd8106
; 
32'd174597: dataIn1 = 32'd8109
; 
32'd174598: dataIn1 = 32'd9110
; 
32'd174599: dataIn1 = 32'd9113
; 
32'd174600: dataIn1 = 32'd2661
; 
32'd174601: dataIn1 = 32'd4995
; 
32'd174602: dataIn1 = 32'd4997
; 
32'd174603: dataIn1 = 32'd8092
; 
32'd174604: dataIn1 = 32'd8107
; 
32'd174605: dataIn1 = 32'd8110
; 
32'd174606: dataIn1 = 32'd9
; 
32'd174607: dataIn1 = 32'd6382
; 
32'd174608: dataIn1 = 32'd8108
; 
32'd174609: dataIn1 = 32'd8111
; 
32'd174610: dataIn1 = 32'd8112
; 
32'd174611: dataIn1 = 32'd8219
; 
32'd174612: dataIn1 = 32'd9111
; 
32'd174613: dataIn1 = 32'd9
; 
32'd174614: dataIn1 = 32'd4734
; 
32'd174615: dataIn1 = 32'd4997
; 
32'd174616: dataIn1 = 32'd8108
; 
32'd174617: dataIn1 = 32'd8111
; 
32'd174618: dataIn1 = 32'd8112
; 
32'd174619: dataIn1 = 32'd6384
; 
32'd174620: dataIn1 = 32'd6385
; 
32'd174621: dataIn1 = 32'd8113
; 
32'd174622: dataIn1 = 32'd8114
; 
32'd174623: dataIn1 = 32'd8115
; 
32'd174624: dataIn1 = 32'd8116
; 
32'd174625: dataIn1 = 32'd8117
; 
32'd174626: dataIn1 = 32'd6383
; 
32'd174627: dataIn1 = 32'd6385
; 
32'd174628: dataIn1 = 32'd8113
; 
32'd174629: dataIn1 = 32'd8114
; 
32'd174630: dataIn1 = 32'd8115
; 
32'd174631: dataIn1 = 32'd8118
; 
32'd174632: dataIn1 = 32'd8119
; 
32'd174633: dataIn1 = 32'd6383
; 
32'd174634: dataIn1 = 32'd6384
; 
32'd174635: dataIn1 = 32'd8113
; 
32'd174636: dataIn1 = 32'd8114
; 
32'd174637: dataIn1 = 32'd8115
; 
32'd174638: dataIn1 = 32'd8120
; 
32'd174639: dataIn1 = 32'd8121
; 
32'd174640: dataIn1 = 32'd5207
; 
32'd174641: dataIn1 = 32'd6385
; 
32'd174642: dataIn1 = 32'd8113
; 
32'd174643: dataIn1 = 32'd8116
; 
32'd174644: dataIn1 = 32'd8117
; 
32'd174645: dataIn1 = 32'd8129
; 
32'd174646: dataIn1 = 32'd8132
; 
32'd174647: dataIn1 = 32'd5207
; 
32'd174648: dataIn1 = 32'd6384
; 
32'd174649: dataIn1 = 32'd6389
; 
32'd174650: dataIn1 = 32'd8113
; 
32'd174651: dataIn1 = 32'd8116
; 
32'd174652: dataIn1 = 32'd8117
; 
32'd174653: dataIn1 = 32'd5208
; 
32'd174654: dataIn1 = 32'd6385
; 
32'd174655: dataIn1 = 32'd8114
; 
32'd174656: dataIn1 = 32'd8118
; 
32'd174657: dataIn1 = 32'd8119
; 
32'd174658: dataIn1 = 32'd8130
; 
32'd174659: dataIn1 = 32'd8133
; 
32'd174660: dataIn1 = 32'd5208
; 
32'd174661: dataIn1 = 32'd6383
; 
32'd174662: dataIn1 = 32'd8114
; 
32'd174663: dataIn1 = 32'd8118
; 
32'd174664: dataIn1 = 32'd8119
; 
32'd174665: dataIn1 = 32'd8123
; 
32'd174666: dataIn1 = 32'd8127
; 
32'd174667: dataIn1 = 32'd5209
; 
32'd174668: dataIn1 = 32'd6384
; 
32'd174669: dataIn1 = 32'd6388
; 
32'd174670: dataIn1 = 32'd8115
; 
32'd174671: dataIn1 = 32'd8120
; 
32'd174672: dataIn1 = 32'd8121
; 
32'd174673: dataIn1 = 32'd5209
; 
32'd174674: dataIn1 = 32'd6383
; 
32'd174675: dataIn1 = 32'd8115
; 
32'd174676: dataIn1 = 32'd8120
; 
32'd174677: dataIn1 = 32'd8121
; 
32'd174678: dataIn1 = 32'd8124
; 
32'd174679: dataIn1 = 32'd8128
; 
32'd174680: dataIn1 = 32'd6386
; 
32'd174681: dataIn1 = 32'd6387
; 
32'd174682: dataIn1 = 32'd8122
; 
32'd174683: dataIn1 = 32'd8123
; 
32'd174684: dataIn1 = 32'd8124
; 
32'd174685: dataIn1 = 32'd8125
; 
32'd174686: dataIn1 = 32'd8126
; 
32'd174687: dataIn1 = 32'd6383
; 
32'd174688: dataIn1 = 32'd6387
; 
32'd174689: dataIn1 = 32'd8119
; 
32'd174690: dataIn1 = 32'd8122
; 
32'd174691: dataIn1 = 32'd8123
; 
32'd174692: dataIn1 = 32'd8124
; 
32'd174693: dataIn1 = 32'd8127
; 
32'd174694: dataIn1 = 32'd6383
; 
32'd174695: dataIn1 = 32'd6386
; 
32'd174696: dataIn1 = 32'd8121
; 
32'd174697: dataIn1 = 32'd8122
; 
32'd174698: dataIn1 = 32'd8123
; 
32'd174699: dataIn1 = 32'd8124
; 
32'd174700: dataIn1 = 32'd8128
; 
32'd174701: dataIn1 = 32'd2719
; 
32'd174702: dataIn1 = 32'd6387
; 
32'd174703: dataIn1 = 32'd8122
; 
32'd174704: dataIn1 = 32'd8125
; 
32'd174705: dataIn1 = 32'd8126
; 
32'd174706: dataIn1 = 32'd8152
; 
32'd174707: dataIn1 = 32'd8155
; 
32'd174708: dataIn1 = 32'd2719
; 
32'd174709: dataIn1 = 32'd6386
; 
32'd174710: dataIn1 = 32'd8122
; 
32'd174711: dataIn1 = 32'd8125
; 
32'd174712: dataIn1 = 32'd8126
; 
32'd174713: dataIn1 = 32'd8169
; 
32'd174714: dataIn1 = 32'd8172
; 
32'd174715: dataIn1 = 32'd5208
; 
32'd174716: dataIn1 = 32'd6387
; 
32'd174717: dataIn1 = 32'd8119
; 
32'd174718: dataIn1 = 32'd8123
; 
32'd174719: dataIn1 = 32'd8127
; 
32'd174720: dataIn1 = 32'd8149
; 
32'd174721: dataIn1 = 32'd8153
; 
32'd174722: dataIn1 = 32'd5209
; 
32'd174723: dataIn1 = 32'd6386
; 
32'd174724: dataIn1 = 32'd8121
; 
32'd174725: dataIn1 = 32'd8124
; 
32'd174726: dataIn1 = 32'd8128
; 
32'd174727: dataIn1 = 32'd8171
; 
32'd174728: dataIn1 = 32'd8175
; 
32'd174729: dataIn1 = 32'd6385
; 
32'd174730: dataIn1 = 32'd6391
; 
32'd174731: dataIn1 = 32'd8116
; 
32'd174732: dataIn1 = 32'd8129
; 
32'd174733: dataIn1 = 32'd8130
; 
32'd174734: dataIn1 = 32'd8131
; 
32'd174735: dataIn1 = 32'd8132
; 
32'd174736: dataIn1 = 32'd6385
; 
32'd174737: dataIn1 = 32'd6390
; 
32'd174738: dataIn1 = 32'd8118
; 
32'd174739: dataIn1 = 32'd8129
; 
32'd174740: dataIn1 = 32'd8130
; 
32'd174741: dataIn1 = 32'd8131
; 
32'd174742: dataIn1 = 32'd8133
; 
32'd174743: dataIn1 = 32'd6390
; 
32'd174744: dataIn1 = 32'd6391
; 
32'd174745: dataIn1 = 32'd8129
; 
32'd174746: dataIn1 = 32'd8130
; 
32'd174747: dataIn1 = 32'd8131
; 
32'd174748: dataIn1 = 32'd8134
; 
32'd174749: dataIn1 = 32'd8135
; 
32'd174750: dataIn1 = 32'd5207
; 
32'd174751: dataIn1 = 32'd6391
; 
32'd174752: dataIn1 = 32'd8116
; 
32'd174753: dataIn1 = 32'd8129
; 
32'd174754: dataIn1 = 32'd8132
; 
32'd174755: dataIn1 = 32'd8136
; 
32'd174756: dataIn1 = 32'd8139
; 
32'd174757: dataIn1 = 32'd5208
; 
32'd174758: dataIn1 = 32'd6390
; 
32'd174759: dataIn1 = 32'd8118
; 
32'd174760: dataIn1 = 32'd8130
; 
32'd174761: dataIn1 = 32'd8133
; 
32'd174762: dataIn1 = 32'd8148
; 
32'd174763: dataIn1 = 32'd8165
; 
32'd174764: dataIn1 = 32'd2721
; 
32'd174765: dataIn1 = 32'd6391
; 
32'd174766: dataIn1 = 32'd8131
; 
32'd174767: dataIn1 = 32'd8134
; 
32'd174768: dataIn1 = 32'd8135
; 
32'd174769: dataIn1 = 32'd8138
; 
32'd174770: dataIn1 = 32'd8142
; 
32'd174771: dataIn1 = 32'd2721
; 
32'd174772: dataIn1 = 32'd6390
; 
32'd174773: dataIn1 = 32'd8131
; 
32'd174774: dataIn1 = 32'd8134
; 
32'd174775: dataIn1 = 32'd8135
; 
32'd174776: dataIn1 = 32'd8166
; 
32'd174777: dataIn1 = 32'd8168
; 
32'd174778: dataIn1 = 32'd6391
; 
32'd174779: dataIn1 = 32'd6394
; 
32'd174780: dataIn1 = 32'd8132
; 
32'd174781: dataIn1 = 32'd8136
; 
32'd174782: dataIn1 = 32'd8137
; 
32'd174783: dataIn1 = 32'd8138
; 
32'd174784: dataIn1 = 32'd8139
; 
32'd174785: dataIn1 = 32'd6394
; 
32'd174786: dataIn1 = 32'd6398
; 
32'd174787: dataIn1 = 32'd8136
; 
32'd174788: dataIn1 = 32'd8137
; 
32'd174789: dataIn1 = 32'd8138
; 
32'd174790: dataIn1 = 32'd8140
; 
32'd174791: dataIn1 = 32'd8141
; 
32'd174792: dataIn1 = 32'd6391
; 
32'd174793: dataIn1 = 32'd6398
; 
32'd174794: dataIn1 = 32'd8134
; 
32'd174795: dataIn1 = 32'd8136
; 
32'd174796: dataIn1 = 32'd8137
; 
32'd174797: dataIn1 = 32'd8138
; 
32'd174798: dataIn1 = 32'd8142
; 
32'd174799: dataIn1 = 32'd5207
; 
32'd174800: dataIn1 = 32'd6394
; 
32'd174801: dataIn1 = 32'd8132
; 
32'd174802: dataIn1 = 32'd8136
; 
32'd174803: dataIn1 = 32'd8139
; 
32'd174804: dataIn1 = 32'd9735
; 
32'd174805: dataIn1 = 32'd9765
; 
32'd174806: dataIn1 = 32'd5210
; 
32'd174807: dataIn1 = 32'd6394
; 
32'd174808: dataIn1 = 32'd8137
; 
32'd174809: dataIn1 = 32'd8140
; 
32'd174810: dataIn1 = 32'd8141
; 
32'd174811: dataIn1 = 32'd9736
; 
32'd174812: dataIn1 = 32'd9766
; 
32'd174813: dataIn1 = 32'd5210
; 
32'd174814: dataIn1 = 32'd6398
; 
32'd174815: dataIn1 = 32'd8137
; 
32'd174816: dataIn1 = 32'd8140
; 
32'd174817: dataIn1 = 32'd8141
; 
32'd174818: dataIn1 = 32'd8306
; 
32'd174819: dataIn1 = 32'd8315
; 
32'd174820: dataIn1 = 32'd2721
; 
32'd174821: dataIn1 = 32'd6398
; 
32'd174822: dataIn1 = 32'd8134
; 
32'd174823: dataIn1 = 32'd8138
; 
32'd174824: dataIn1 = 32'd8142
; 
32'd174825: dataIn1 = 32'd8299
; 
32'd174826: dataIn1 = 32'd8316
; 
32'd174827: dataIn1 = 32'd6400
; 
32'd174828: dataIn1 = 32'd6401
; 
32'd174829: dataIn1 = 32'd8143
; 
32'd174830: dataIn1 = 32'd8144
; 
32'd174831: dataIn1 = 32'd8145
; 
32'd174832: dataIn1 = 32'd8146
; 
32'd174833: dataIn1 = 32'd8147
; 
32'd174834: dataIn1 = 32'd6399
; 
32'd174835: dataIn1 = 32'd6401
; 
32'd174836: dataIn1 = 32'd8143
; 
32'd174837: dataIn1 = 32'd8144
; 
32'd174838: dataIn1 = 32'd8145
; 
32'd174839: dataIn1 = 32'd8148
; 
32'd174840: dataIn1 = 32'd8149
; 
32'd174841: dataIn1 = 32'd6399
; 
32'd174842: dataIn1 = 32'd6400
; 
32'd174843: dataIn1 = 32'd8143
; 
32'd174844: dataIn1 = 32'd8144
; 
32'd174845: dataIn1 = 32'd8145
; 
32'd174846: dataIn1 = 32'd8150
; 
32'd174847: dataIn1 = 32'd8151
; 
32'd174848: dataIn1 = 32'd5212
; 
32'd174849: dataIn1 = 32'd6401
; 
32'd174850: dataIn1 = 32'd8143
; 
32'd174851: dataIn1 = 32'd8146
; 
32'd174852: dataIn1 = 32'd8147
; 
32'd174853: dataIn1 = 32'd8164
; 
32'd174854: dataIn1 = 32'd8167
; 
32'd174855: dataIn1 = 32'd5212
; 
32'd174856: dataIn1 = 32'd6400
; 
32'd174857: dataIn1 = 32'd8143
; 
32'd174858: dataIn1 = 32'd8146
; 
32'd174859: dataIn1 = 32'd8147
; 
32'd174860: dataIn1 = 32'd8157
; 
32'd174861: dataIn1 = 32'd8160
; 
32'd174862: dataIn1 = 32'd5208
; 
32'd174863: dataIn1 = 32'd6401
; 
32'd174864: dataIn1 = 32'd8133
; 
32'd174865: dataIn1 = 32'd8144
; 
32'd174866: dataIn1 = 32'd8148
; 
32'd174867: dataIn1 = 32'd8149
; 
32'd174868: dataIn1 = 32'd8165
; 
32'd174869: dataIn1 = 32'd5208
; 
32'd174870: dataIn1 = 32'd6399
; 
32'd174871: dataIn1 = 32'd8127
; 
32'd174872: dataIn1 = 32'd8144
; 
32'd174873: dataIn1 = 32'd8148
; 
32'd174874: dataIn1 = 32'd8149
; 
32'd174875: dataIn1 = 32'd8153
; 
32'd174876: dataIn1 = 32'd5213
; 
32'd174877: dataIn1 = 32'd6400
; 
32'd174878: dataIn1 = 32'd8145
; 
32'd174879: dataIn1 = 32'd8150
; 
32'd174880: dataIn1 = 32'd8151
; 
32'd174881: dataIn1 = 32'd8159
; 
32'd174882: dataIn1 = 32'd8163
; 
32'd174883: dataIn1 = 32'd5213
; 
32'd174884: dataIn1 = 32'd6399
; 
32'd174885: dataIn1 = 32'd8145
; 
32'd174886: dataIn1 = 32'd8150
; 
32'd174887: dataIn1 = 32'd8151
; 
32'd174888: dataIn1 = 32'd8154
; 
32'd174889: dataIn1 = 32'd8156
; 
32'd174890: dataIn1 = 32'd6387
; 
32'd174891: dataIn1 = 32'd6402
; 
32'd174892: dataIn1 = 32'd8125
; 
32'd174893: dataIn1 = 32'd8152
; 
32'd174894: dataIn1 = 32'd8153
; 
32'd174895: dataIn1 = 32'd8154
; 
32'd174896: dataIn1 = 32'd8155
; 
32'd174897: dataIn1 = 32'd6387
; 
32'd174898: dataIn1 = 32'd6399
; 
32'd174899: dataIn1 = 32'd8127
; 
32'd174900: dataIn1 = 32'd8149
; 
32'd174901: dataIn1 = 32'd8152
; 
32'd174902: dataIn1 = 32'd8153
; 
32'd174903: dataIn1 = 32'd8154
; 
32'd174904: dataIn1 = 32'd6399
; 
32'd174905: dataIn1 = 32'd6402
; 
32'd174906: dataIn1 = 32'd8151
; 
32'd174907: dataIn1 = 32'd8152
; 
32'd174908: dataIn1 = 32'd8153
; 
32'd174909: dataIn1 = 32'd8154
; 
32'd174910: dataIn1 = 32'd8156
; 
32'd174911: dataIn1 = 32'd2719
; 
32'd174912: dataIn1 = 32'd6402
; 
32'd174913: dataIn1 = 32'd8125
; 
32'd174914: dataIn1 = 32'd8152
; 
32'd174915: dataIn1 = 32'd8155
; 
32'd174916: dataIn1 = 32'd8188
; 
32'd174917: dataIn1 = 32'd8241
; 
32'd174918: dataIn1 = 32'd5213
; 
32'd174919: dataIn1 = 32'd6402
; 
32'd174920: dataIn1 = 32'd8151
; 
32'd174921: dataIn1 = 32'd8154
; 
32'd174922: dataIn1 = 32'd8156
; 
32'd174923: dataIn1 = 32'd8240
; 
32'd174924: dataIn1 = 32'd8243
; 
32'd174925: dataIn1 = 32'd6400
; 
32'd174926: dataIn1 = 32'd6404
; 
32'd174927: dataIn1 = 32'd8147
; 
32'd174928: dataIn1 = 32'd8157
; 
32'd174929: dataIn1 = 32'd8158
; 
32'd174930: dataIn1 = 32'd8159
; 
32'd174931: dataIn1 = 32'd8160
; 
32'd174932: dataIn1 = 32'd6403
; 
32'd174933: dataIn1 = 32'd6404
; 
32'd174934: dataIn1 = 32'd8157
; 
32'd174935: dataIn1 = 32'd8158
; 
32'd174936: dataIn1 = 32'd8159
; 
32'd174937: dataIn1 = 32'd8161
; 
32'd174938: dataIn1 = 32'd8162
; 
32'd174939: dataIn1 = 32'd6400
; 
32'd174940: dataIn1 = 32'd6403
; 
32'd174941: dataIn1 = 32'd8150
; 
32'd174942: dataIn1 = 32'd8157
; 
32'd174943: dataIn1 = 32'd8158
; 
32'd174944: dataIn1 = 32'd8159
; 
32'd174945: dataIn1 = 32'd8163
; 
32'd174946: dataIn1 = 32'd5212
; 
32'd174947: dataIn1 = 32'd6404
; 
32'd174948: dataIn1 = 32'd8147
; 
32'd174949: dataIn1 = 32'd8157
; 
32'd174950: dataIn1 = 32'd8160
; 
32'd174951: dataIn1 = 32'd8321
; 
32'd174952: dataIn1 = 32'd8331
; 
32'd174953: dataIn1 = 32'd142
; 
32'd174954: dataIn1 = 32'd6404
; 
32'd174955: dataIn1 = 32'd8158
; 
32'd174956: dataIn1 = 32'd8161
; 
32'd174957: dataIn1 = 32'd8162
; 
32'd174958: dataIn1 = 32'd8332
; 
32'd174959: dataIn1 = 32'd8334
; 
32'd174960: dataIn1 = 32'd142
; 
32'd174961: dataIn1 = 32'd6403
; 
32'd174962: dataIn1 = 32'd8158
; 
32'd174963: dataIn1 = 32'd8161
; 
32'd174964: dataIn1 = 32'd8162
; 
32'd174965: dataIn1 = 32'd8245
; 
32'd174966: dataIn1 = 32'd8248
; 
32'd174967: dataIn1 = 32'd5213
; 
32'd174968: dataIn1 = 32'd6403
; 
32'd174969: dataIn1 = 32'd8150
; 
32'd174970: dataIn1 = 32'd8159
; 
32'd174971: dataIn1 = 32'd8163
; 
32'd174972: dataIn1 = 32'd8239
; 
32'd174973: dataIn1 = 32'd8246
; 
32'd174974: dataIn1 = 32'd6401
; 
32'd174975: dataIn1 = 32'd6405
; 
32'd174976: dataIn1 = 32'd8146
; 
32'd174977: dataIn1 = 32'd8164
; 
32'd174978: dataIn1 = 32'd8165
; 
32'd174979: dataIn1 = 32'd8166
; 
32'd174980: dataIn1 = 32'd8167
; 
32'd174981: dataIn1 = 32'd6390
; 
32'd174982: dataIn1 = 32'd6401
; 
32'd174983: dataIn1 = 32'd8133
; 
32'd174984: dataIn1 = 32'd8148
; 
32'd174985: dataIn1 = 32'd8164
; 
32'd174986: dataIn1 = 32'd8165
; 
32'd174987: dataIn1 = 32'd8166
; 
32'd174988: dataIn1 = 32'd6390
; 
32'd174989: dataIn1 = 32'd6405
; 
32'd174990: dataIn1 = 32'd8135
; 
32'd174991: dataIn1 = 32'd8164
; 
32'd174992: dataIn1 = 32'd8165
; 
32'd174993: dataIn1 = 32'd8166
; 
32'd174994: dataIn1 = 32'd8168
; 
32'd174995: dataIn1 = 32'd5212
; 
32'd174996: dataIn1 = 32'd6405
; 
32'd174997: dataIn1 = 32'd8146
; 
32'd174998: dataIn1 = 32'd8164
; 
32'd174999: dataIn1 = 32'd8167
; 
32'd175000: dataIn1 = 32'd8320
; 
32'd175001: dataIn1 = 32'd8336
; 
32'd175002: dataIn1 = 32'd2721
; 
32'd175003: dataIn1 = 32'd6405
; 
32'd175004: dataIn1 = 32'd8135
; 
32'd175005: dataIn1 = 32'd8166
; 
32'd175006: dataIn1 = 32'd8168
; 
32'd175007: dataIn1 = 32'd8300
; 
32'd175008: dataIn1 = 32'd8338
; 
32'd175009: dataIn1 = 32'd6386
; 
32'd175010: dataIn1 = 32'd6407
; 
32'd175011: dataIn1 = 32'd8126
; 
32'd175012: dataIn1 = 32'd8169
; 
32'd175013: dataIn1 = 32'd8170
; 
32'd175014: dataIn1 = 32'd8171
; 
32'd175015: dataIn1 = 32'd8172
; 
32'd175016: dataIn1 = 32'd6406
; 
32'd175017: dataIn1 = 32'd6407
; 
32'd175018: dataIn1 = 32'd8169
; 
32'd175019: dataIn1 = 32'd8170
; 
32'd175020: dataIn1 = 32'd8171
; 
32'd175021: dataIn1 = 32'd8173
; 
32'd175022: dataIn1 = 32'd8174
; 
32'd175023: dataIn1 = 32'd6386
; 
32'd175024: dataIn1 = 32'd6406
; 
32'd175025: dataIn1 = 32'd8128
; 
32'd175026: dataIn1 = 32'd8169
; 
32'd175027: dataIn1 = 32'd8170
; 
32'd175028: dataIn1 = 32'd8171
; 
32'd175029: dataIn1 = 32'd8175
; 
32'd175030: dataIn1 = 32'd2719
; 
32'd175031: dataIn1 = 32'd6407
; 
32'd175032: dataIn1 = 32'd8126
; 
32'd175033: dataIn1 = 32'd8169
; 
32'd175034: dataIn1 = 32'd8172
; 
32'd175035: dataIn1 = 32'd8189
; 
32'd175036: dataIn1 = 32'd8263
; 
32'd175037: dataIn1 = 32'd5215
; 
32'd175038: dataIn1 = 32'd6407
; 
32'd175039: dataIn1 = 32'd8170
; 
32'd175040: dataIn1 = 32'd8173
; 
32'd175041: dataIn1 = 32'd8174
; 
32'd175042: dataIn1 = 32'd8260
; 
32'd175043: dataIn1 = 32'd8264
; 
32'd175044: dataIn1 = 32'd5215
; 
32'd175045: dataIn1 = 32'd6406
; 
32'd175046: dataIn1 = 32'd6714
; 
32'd175047: dataIn1 = 32'd8170
; 
32'd175048: dataIn1 = 32'd8173
; 
32'd175049: dataIn1 = 32'd8174
; 
32'd175050: dataIn1 = 32'd5209
; 
32'd175051: dataIn1 = 32'd6406
; 
32'd175052: dataIn1 = 32'd6408
; 
32'd175053: dataIn1 = 32'd8128
; 
32'd175054: dataIn1 = 32'd8171
; 
32'd175055: dataIn1 = 32'd8175
; 
32'd175056: dataIn1 = 32'd6411
; 
32'd175057: dataIn1 = 32'd6412
; 
32'd175058: dataIn1 = 32'd8176
; 
32'd175059: dataIn1 = 32'd8177
; 
32'd175060: dataIn1 = 32'd8178
; 
32'd175061: dataIn1 = 32'd8179
; 
32'd175062: dataIn1 = 32'd8180
; 
32'd175063: dataIn1 = 32'd6410
; 
32'd175064: dataIn1 = 32'd6412
; 
32'd175065: dataIn1 = 32'd8176
; 
32'd175066: dataIn1 = 32'd8177
; 
32'd175067: dataIn1 = 32'd8178
; 
32'd175068: dataIn1 = 32'd8181
; 
32'd175069: dataIn1 = 32'd8182
; 
32'd175070: dataIn1 = 32'd6410
; 
32'd175071: dataIn1 = 32'd6411
; 
32'd175072: dataIn1 = 32'd8176
; 
32'd175073: dataIn1 = 32'd8177
; 
32'd175074: dataIn1 = 32'd8178
; 
32'd175075: dataIn1 = 32'd8183
; 
32'd175076: dataIn1 = 32'd8184
; 
32'd175077: dataIn1 = 32'd5216
; 
32'd175078: dataIn1 = 32'd6412
; 
32'd175079: dataIn1 = 32'd8176
; 
32'd175080: dataIn1 = 32'd8179
; 
32'd175081: dataIn1 = 32'd8180
; 
32'd175082: dataIn1 = 32'd8199
; 
32'd175083: dataIn1 = 32'd8202
; 
32'd175084: dataIn1 = 32'd5216
; 
32'd175085: dataIn1 = 32'd6411
; 
32'd175086: dataIn1 = 32'd8176
; 
32'd175087: dataIn1 = 32'd8179
; 
32'd175088: dataIn1 = 32'd8180
; 
32'd175089: dataIn1 = 32'd8192
; 
32'd175090: dataIn1 = 32'd8195
; 
32'd175091: dataIn1 = 32'd5217
; 
32'd175092: dataIn1 = 32'd6412
; 
32'd175093: dataIn1 = 32'd8177
; 
32'd175094: dataIn1 = 32'd8181
; 
32'd175095: dataIn1 = 32'd8182
; 
32'd175096: dataIn1 = 32'd8200
; 
32'd175097: dataIn1 = 32'd8203
; 
32'd175098: dataIn1 = 32'd5217
; 
32'd175099: dataIn1 = 32'd6410
; 
32'd175100: dataIn1 = 32'd8177
; 
32'd175101: dataIn1 = 32'd8181
; 
32'd175102: dataIn1 = 32'd8182
; 
32'd175103: dataIn1 = 32'd8186
; 
32'd175104: dataIn1 = 32'd8190
; 
32'd175105: dataIn1 = 32'd5218
; 
32'd175106: dataIn1 = 32'd6411
; 
32'd175107: dataIn1 = 32'd8178
; 
32'd175108: dataIn1 = 32'd8183
; 
32'd175109: dataIn1 = 32'd8184
; 
32'd175110: dataIn1 = 32'd8194
; 
32'd175111: dataIn1 = 32'd8198
; 
32'd175112: dataIn1 = 32'd5218
; 
32'd175113: dataIn1 = 32'd6410
; 
32'd175114: dataIn1 = 32'd8178
; 
32'd175115: dataIn1 = 32'd8183
; 
32'd175116: dataIn1 = 32'd8184
; 
32'd175117: dataIn1 = 32'd8187
; 
32'd175118: dataIn1 = 32'd8191
; 
32'd175119: dataIn1 = 32'd6413
; 
32'd175120: dataIn1 = 32'd6414
; 
32'd175121: dataIn1 = 32'd8185
; 
32'd175122: dataIn1 = 32'd8186
; 
32'd175123: dataIn1 = 32'd8187
; 
32'd175124: dataIn1 = 32'd8188
; 
32'd175125: dataIn1 = 32'd8189
; 
32'd175126: dataIn1 = 32'd6410
; 
32'd175127: dataIn1 = 32'd6414
; 
32'd175128: dataIn1 = 32'd8182
; 
32'd175129: dataIn1 = 32'd8185
; 
32'd175130: dataIn1 = 32'd8186
; 
32'd175131: dataIn1 = 32'd8187
; 
32'd175132: dataIn1 = 32'd8190
; 
32'd175133: dataIn1 = 32'd6410
; 
32'd175134: dataIn1 = 32'd6413
; 
32'd175135: dataIn1 = 32'd8184
; 
32'd175136: dataIn1 = 32'd8185
; 
32'd175137: dataIn1 = 32'd8186
; 
32'd175138: dataIn1 = 32'd8187
; 
32'd175139: dataIn1 = 32'd8191
; 
32'd175140: dataIn1 = 32'd2719
; 
32'd175141: dataIn1 = 32'd6414
; 
32'd175142: dataIn1 = 32'd8155
; 
32'd175143: dataIn1 = 32'd8185
; 
32'd175144: dataIn1 = 32'd8188
; 
32'd175145: dataIn1 = 32'd8189
; 
32'd175146: dataIn1 = 32'd8241
; 
32'd175147: dataIn1 = 32'd2719
; 
32'd175148: dataIn1 = 32'd6413
; 
32'd175149: dataIn1 = 32'd8172
; 
32'd175150: dataIn1 = 32'd8185
; 
32'd175151: dataIn1 = 32'd8188
; 
32'd175152: dataIn1 = 32'd8189
; 
32'd175153: dataIn1 = 32'd8263
; 
32'd175154: dataIn1 = 32'd5217
; 
32'd175155: dataIn1 = 32'd6414
; 
32'd175156: dataIn1 = 32'd8182
; 
32'd175157: dataIn1 = 32'd8186
; 
32'd175158: dataIn1 = 32'd8190
; 
32'd175159: dataIn1 = 32'd8238
; 
32'd175160: dataIn1 = 32'd8242
; 
32'd175161: dataIn1 = 32'd5218
; 
32'd175162: dataIn1 = 32'd6413
; 
32'd175163: dataIn1 = 32'd8184
; 
32'd175164: dataIn1 = 32'd8187
; 
32'd175165: dataIn1 = 32'd8191
; 
32'd175166: dataIn1 = 32'd8262
; 
32'd175167: dataIn1 = 32'd8265
; 
32'd175168: dataIn1 = 32'd6411
; 
32'd175169: dataIn1 = 32'd6416
; 
32'd175170: dataIn1 = 32'd8180
; 
32'd175171: dataIn1 = 32'd8192
; 
32'd175172: dataIn1 = 32'd8193
; 
32'd175173: dataIn1 = 32'd8194
; 
32'd175174: dataIn1 = 32'd8195
; 
32'd175175: dataIn1 = 32'd6415
; 
32'd175176: dataIn1 = 32'd6416
; 
32'd175177: dataIn1 = 32'd8192
; 
32'd175178: dataIn1 = 32'd8193
; 
32'd175179: dataIn1 = 32'd8194
; 
32'd175180: dataIn1 = 32'd8196
; 
32'd175181: dataIn1 = 32'd8197
; 
32'd175182: dataIn1 = 32'd6411
; 
32'd175183: dataIn1 = 32'd6415
; 
32'd175184: dataIn1 = 32'd8183
; 
32'd175185: dataIn1 = 32'd8192
; 
32'd175186: dataIn1 = 32'd8193
; 
32'd175187: dataIn1 = 32'd8194
; 
32'd175188: dataIn1 = 32'd8198
; 
32'd175189: dataIn1 = 32'd5216
; 
32'd175190: dataIn1 = 32'd6416
; 
32'd175191: dataIn1 = 32'd8180
; 
32'd175192: dataIn1 = 32'd8192
; 
32'd175193: dataIn1 = 32'd8195
; 
32'd175194: dataIn1 = 32'd8210
; 
32'd175195: dataIn1 = 32'd8222
; 
32'd175196: dataIn1 = 32'd2722
; 
32'd175197: dataIn1 = 32'd6416
; 
32'd175198: dataIn1 = 32'd8193
; 
32'd175199: dataIn1 = 32'd8196
; 
32'd175200: dataIn1 = 32'd8197
; 
32'd175201: dataIn1 = 32'd8223
; 
32'd175202: dataIn1 = 32'd8225
; 
32'd175203: dataIn1 = 32'd2722
; 
32'd175204: dataIn1 = 32'd6415
; 
32'd175205: dataIn1 = 32'd8193
; 
32'd175206: dataIn1 = 32'd8196
; 
32'd175207: dataIn1 = 32'd8197
; 
32'd175208: dataIn1 = 32'd8267
; 
32'd175209: dataIn1 = 32'd8270
; 
32'd175210: dataIn1 = 32'd5218
; 
32'd175211: dataIn1 = 32'd6415
; 
32'd175212: dataIn1 = 32'd8183
; 
32'd175213: dataIn1 = 32'd8194
; 
32'd175214: dataIn1 = 32'd8198
; 
32'd175215: dataIn1 = 32'd8261
; 
32'd175216: dataIn1 = 32'd8268
; 
32'd175217: dataIn1 = 32'd6412
; 
32'd175218: dataIn1 = 32'd6418
; 
32'd175219: dataIn1 = 32'd8179
; 
32'd175220: dataIn1 = 32'd8199
; 
32'd175221: dataIn1 = 32'd8200
; 
32'd175222: dataIn1 = 32'd8201
; 
32'd175223: dataIn1 = 32'd8202
; 
32'd175224: dataIn1 = 32'd6412
; 
32'd175225: dataIn1 = 32'd6417
; 
32'd175226: dataIn1 = 32'd8181
; 
32'd175227: dataIn1 = 32'd8199
; 
32'd175228: dataIn1 = 32'd8200
; 
32'd175229: dataIn1 = 32'd8201
; 
32'd175230: dataIn1 = 32'd8203
; 
32'd175231: dataIn1 = 32'd6417
; 
32'd175232: dataIn1 = 32'd6418
; 
32'd175233: dataIn1 = 32'd8199
; 
32'd175234: dataIn1 = 32'd8200
; 
32'd175235: dataIn1 = 32'd8201
; 
32'd175236: dataIn1 = 32'd8204
; 
32'd175237: dataIn1 = 32'd8205
; 
32'd175238: dataIn1 = 32'd5216
; 
32'd175239: dataIn1 = 32'd6418
; 
32'd175240: dataIn1 = 32'd8179
; 
32'd175241: dataIn1 = 32'd8199
; 
32'd175242: dataIn1 = 32'd8202
; 
32'd175243: dataIn1 = 32'd8209
; 
32'd175244: dataIn1 = 32'd8227
; 
32'd175245: dataIn1 = 32'd5217
; 
32'd175246: dataIn1 = 32'd6417
; 
32'd175247: dataIn1 = 32'd8181
; 
32'd175248: dataIn1 = 32'd8200
; 
32'd175249: dataIn1 = 32'd8203
; 
32'd175250: dataIn1 = 32'd8237
; 
32'd175251: dataIn1 = 32'd8250
; 
32'd175252: dataIn1 = 32'd1113
; 
32'd175253: dataIn1 = 32'd6418
; 
32'd175254: dataIn1 = 32'd8201
; 
32'd175255: dataIn1 = 32'd8204
; 
32'd175256: dataIn1 = 32'd8205
; 
32'd175257: dataIn1 = 32'd8229
; 
32'd175258: dataIn1 = 32'd8231
; 
32'd175259: dataIn1 = 32'd1113
; 
32'd175260: dataIn1 = 32'd6417
; 
32'd175261: dataIn1 = 32'd8201
; 
32'd175262: dataIn1 = 32'd8204
; 
32'd175263: dataIn1 = 32'd8205
; 
32'd175264: dataIn1 = 32'd8251
; 
32'd175265: dataIn1 = 32'd8253
; 
32'd175266: dataIn1 = 32'd6420
; 
32'd175267: dataIn1 = 32'd6421
; 
32'd175268: dataIn1 = 32'd8206
; 
32'd175269: dataIn1 = 32'd8207
; 
32'd175270: dataIn1 = 32'd8208
; 
32'd175271: dataIn1 = 32'd8209
; 
32'd175272: dataIn1 = 32'd8210
; 
32'd175273: dataIn1 = 32'd6419
; 
32'd175274: dataIn1 = 32'd6421
; 
32'd175275: dataIn1 = 32'd8206
; 
32'd175276: dataIn1 = 32'd8207
; 
32'd175277: dataIn1 = 32'd8208
; 
32'd175278: dataIn1 = 32'd8211
; 
32'd175279: dataIn1 = 32'd8212
; 
32'd175280: dataIn1 = 32'd6419
; 
32'd175281: dataIn1 = 32'd6420
; 
32'd175282: dataIn1 = 32'd8206
; 
32'd175283: dataIn1 = 32'd8207
; 
32'd175284: dataIn1 = 32'd8208
; 
32'd175285: dataIn1 = 32'd8213
; 
32'd175286: dataIn1 = 32'd8214
; 
32'd175287: dataIn1 = 32'd5216
; 
32'd175288: dataIn1 = 32'd6421
; 
32'd175289: dataIn1 = 32'd8202
; 
32'd175290: dataIn1 = 32'd8206
; 
32'd175291: dataIn1 = 32'd8209
; 
32'd175292: dataIn1 = 32'd8210
; 
32'd175293: dataIn1 = 32'd8227
; 
32'd175294: dataIn1 = 32'd5216
; 
32'd175295: dataIn1 = 32'd6420
; 
32'd175296: dataIn1 = 32'd8195
; 
32'd175297: dataIn1 = 32'd8206
; 
32'd175298: dataIn1 = 32'd8209
; 
32'd175299: dataIn1 = 32'd8210
; 
32'd175300: dataIn1 = 32'd8222
; 
32'd175301: dataIn1 = 32'd2666
; 
32'd175302: dataIn1 = 32'd6421
; 
32'd175303: dataIn1 = 32'd8207
; 
32'd175304: dataIn1 = 32'd8211
; 
32'd175305: dataIn1 = 32'd8212
; 
32'd175306: dataIn1 = 32'd8228
; 
32'd175307: dataIn1 = 32'd8230
; 
32'd175308: dataIn1 = 32'd2666
; 
32'd175309: dataIn1 = 32'd6419
; 
32'd175310: dataIn1 = 32'd8207
; 
32'd175311: dataIn1 = 32'd8211
; 
32'd175312: dataIn1 = 32'd8212
; 
32'd175313: dataIn1 = 32'd8216
; 
32'd175314: dataIn1 = 32'd8220
; 
32'd175315: dataIn1 = 32'd5219
; 
32'd175316: dataIn1 = 32'd6420
; 
32'd175317: dataIn1 = 32'd8208
; 
32'd175318: dataIn1 = 32'd8213
; 
32'd175319: dataIn1 = 32'd8214
; 
32'd175320: dataIn1 = 32'd8224
; 
32'd175321: dataIn1 = 32'd8226
; 
32'd175322: dataIn1 = 32'd5219
; 
32'd175323: dataIn1 = 32'd6419
; 
32'd175324: dataIn1 = 32'd8208
; 
32'd175325: dataIn1 = 32'd8213
; 
32'd175326: dataIn1 = 32'd8214
; 
32'd175327: dataIn1 = 32'd8217
; 
32'd175328: dataIn1 = 32'd8221
; 
32'd175329: dataIn1 = 32'd5015
; 
32'd175330: dataIn1 = 32'd6422
; 
32'd175331: dataIn1 = 32'd8215
; 
32'd175332: dataIn1 = 32'd8216
; 
32'd175333: dataIn1 = 32'd8217
; 
32'd175334: dataIn1 = 32'd8218
; 
32'd175335: dataIn1 = 32'd8219
; 
32'd175336: dataIn1 = 32'd5015
; 
32'd175337: dataIn1 = 32'd6419
; 
32'd175338: dataIn1 = 32'd8212
; 
32'd175339: dataIn1 = 32'd8215
; 
32'd175340: dataIn1 = 32'd8216
; 
32'd175341: dataIn1 = 32'd8217
; 
32'd175342: dataIn1 = 32'd8220
; 
32'd175343: dataIn1 = 32'd6419
; 
32'd175344: dataIn1 = 32'd6422
; 
32'd175345: dataIn1 = 32'd8214
; 
32'd175346: dataIn1 = 32'd8215
; 
32'd175347: dataIn1 = 32'd8216
; 
32'd175348: dataIn1 = 32'd8217
; 
32'd175349: dataIn1 = 32'd8221
; 
32'd175350: dataIn1 = 32'd9
; 
32'd175351: dataIn1 = 32'd4735
; 
32'd175352: dataIn1 = 32'd5015
; 
32'd175353: dataIn1 = 32'd8215
; 
32'd175354: dataIn1 = 32'd8218
; 
32'd175355: dataIn1 = 32'd8219
; 
32'd175356: dataIn1 = 32'd9
; 
32'd175357: dataIn1 = 32'd6422
; 
32'd175358: dataIn1 = 32'd8111
; 
32'd175359: dataIn1 = 32'd8215
; 
32'd175360: dataIn1 = 32'd8218
; 
32'd175361: dataIn1 = 32'd8219
; 
32'd175362: dataIn1 = 32'd9111
; 
32'd175363: dataIn1 = 32'd2666
; 
32'd175364: dataIn1 = 32'd5013
; 
32'd175365: dataIn1 = 32'd5015
; 
32'd175366: dataIn1 = 32'd8212
; 
32'd175367: dataIn1 = 32'd8216
; 
32'd175368: dataIn1 = 32'd8220
; 
32'd175369: dataIn1 = 32'd5219
; 
32'd175370: dataIn1 = 32'd6422
; 
32'd175371: dataIn1 = 32'd8214
; 
32'd175372: dataIn1 = 32'd8217
; 
32'd175373: dataIn1 = 32'd8221
; 
32'd175374: dataIn1 = 32'd9108
; 
32'd175375: dataIn1 = 32'd9112
; 
32'd175376: dataIn1 = 32'd6416
; 
32'd175377: dataIn1 = 32'd6420
; 
32'd175378: dataIn1 = 32'd8195
; 
32'd175379: dataIn1 = 32'd8210
; 
32'd175380: dataIn1 = 32'd8222
; 
32'd175381: dataIn1 = 32'd8223
; 
32'd175382: dataIn1 = 32'd8224
; 
32'd175383: dataIn1 = 32'd6416
; 
32'd175384: dataIn1 = 32'd6423
; 
32'd175385: dataIn1 = 32'd8196
; 
32'd175386: dataIn1 = 32'd8222
; 
32'd175387: dataIn1 = 32'd8223
; 
32'd175388: dataIn1 = 32'd8224
; 
32'd175389: dataIn1 = 32'd8225
; 
32'd175390: dataIn1 = 32'd6420
; 
32'd175391: dataIn1 = 32'd6423
; 
32'd175392: dataIn1 = 32'd8213
; 
32'd175393: dataIn1 = 32'd8222
; 
32'd175394: dataIn1 = 32'd8223
; 
32'd175395: dataIn1 = 32'd8224
; 
32'd175396: dataIn1 = 32'd8226
; 
32'd175397: dataIn1 = 32'd2722
; 
32'd175398: dataIn1 = 32'd6423
; 
32'd175399: dataIn1 = 32'd8196
; 
32'd175400: dataIn1 = 32'd8223
; 
32'd175401: dataIn1 = 32'd8225
; 
32'd175402: dataIn1 = 32'd9100
; 
32'd175403: dataIn1 = 32'd9119
; 
32'd175404: dataIn1 = 32'd5219
; 
32'd175405: dataIn1 = 32'd6423
; 
32'd175406: dataIn1 = 32'd8213
; 
32'd175407: dataIn1 = 32'd8224
; 
32'd175408: dataIn1 = 32'd8226
; 
32'd175409: dataIn1 = 32'd9107
; 
32'd175410: dataIn1 = 32'd9118
; 
32'd175411: dataIn1 = 32'd6418
; 
32'd175412: dataIn1 = 32'd6421
; 
32'd175413: dataIn1 = 32'd8202
; 
32'd175414: dataIn1 = 32'd8209
; 
32'd175415: dataIn1 = 32'd8227
; 
32'd175416: dataIn1 = 32'd8228
; 
32'd175417: dataIn1 = 32'd8229
; 
32'd175418: dataIn1 = 32'd5016
; 
32'd175419: dataIn1 = 32'd6421
; 
32'd175420: dataIn1 = 32'd8211
; 
32'd175421: dataIn1 = 32'd8227
; 
32'd175422: dataIn1 = 32'd8228
; 
32'd175423: dataIn1 = 32'd8229
; 
32'd175424: dataIn1 = 32'd8230
; 
32'd175425: dataIn1 = 32'd5016
; 
32'd175426: dataIn1 = 32'd6418
; 
32'd175427: dataIn1 = 32'd8204
; 
32'd175428: dataIn1 = 32'd8227
; 
32'd175429: dataIn1 = 32'd8228
; 
32'd175430: dataIn1 = 32'd8229
; 
32'd175431: dataIn1 = 32'd8231
; 
32'd175432: dataIn1 = 32'd2666
; 
32'd175433: dataIn1 = 32'd5014
; 
32'd175434: dataIn1 = 32'd5016
; 
32'd175435: dataIn1 = 32'd8211
; 
32'd175436: dataIn1 = 32'd8228
; 
32'd175437: dataIn1 = 32'd8230
; 
32'd175438: dataIn1 = 32'd1113
; 
32'd175439: dataIn1 = 32'd5005
; 
32'd175440: dataIn1 = 32'd5016
; 
32'd175441: dataIn1 = 32'd8204
; 
32'd175442: dataIn1 = 32'd8229
; 
32'd175443: dataIn1 = 32'd8231
; 
32'd175444: dataIn1 = 32'd6425
; 
32'd175445: dataIn1 = 32'd6426
; 
32'd175446: dataIn1 = 32'd8232
; 
32'd175447: dataIn1 = 32'd8233
; 
32'd175448: dataIn1 = 32'd8234
; 
32'd175449: dataIn1 = 32'd8235
; 
32'd175450: dataIn1 = 32'd8236
; 
32'd175451: dataIn1 = 32'd6424
; 
32'd175452: dataIn1 = 32'd6426
; 
32'd175453: dataIn1 = 32'd8232
; 
32'd175454: dataIn1 = 32'd8233
; 
32'd175455: dataIn1 = 32'd8234
; 
32'd175456: dataIn1 = 32'd8237
; 
32'd175457: dataIn1 = 32'd8238
; 
32'd175458: dataIn1 = 32'd6424
; 
32'd175459: dataIn1 = 32'd6425
; 
32'd175460: dataIn1 = 32'd8232
; 
32'd175461: dataIn1 = 32'd8233
; 
32'd175462: dataIn1 = 32'd8234
; 
32'd175463: dataIn1 = 32'd8239
; 
32'd175464: dataIn1 = 32'd8240
; 
32'd175465: dataIn1 = 32'd2665
; 
32'd175466: dataIn1 = 32'd6426
; 
32'd175467: dataIn1 = 32'd8232
; 
32'd175468: dataIn1 = 32'd8235
; 
32'd175469: dataIn1 = 32'd8236
; 
32'd175470: dataIn1 = 32'd8249
; 
32'd175471: dataIn1 = 32'd8252
; 
32'd175472: dataIn1 = 32'd2665
; 
32'd175473: dataIn1 = 32'd6425
; 
32'd175474: dataIn1 = 32'd8232
; 
32'd175475: dataIn1 = 32'd8235
; 
32'd175476: dataIn1 = 32'd8236
; 
32'd175477: dataIn1 = 32'd8244
; 
32'd175478: dataIn1 = 32'd8247
; 
32'd175479: dataIn1 = 32'd5217
; 
32'd175480: dataIn1 = 32'd6426
; 
32'd175481: dataIn1 = 32'd8203
; 
32'd175482: dataIn1 = 32'd8233
; 
32'd175483: dataIn1 = 32'd8237
; 
32'd175484: dataIn1 = 32'd8238
; 
32'd175485: dataIn1 = 32'd8250
; 
32'd175486: dataIn1 = 32'd5217
; 
32'd175487: dataIn1 = 32'd6424
; 
32'd175488: dataIn1 = 32'd8190
; 
32'd175489: dataIn1 = 32'd8233
; 
32'd175490: dataIn1 = 32'd8237
; 
32'd175491: dataIn1 = 32'd8238
; 
32'd175492: dataIn1 = 32'd8242
; 
32'd175493: dataIn1 = 32'd5213
; 
32'd175494: dataIn1 = 32'd6425
; 
32'd175495: dataIn1 = 32'd8163
; 
32'd175496: dataIn1 = 32'd8234
; 
32'd175497: dataIn1 = 32'd8239
; 
32'd175498: dataIn1 = 32'd8240
; 
32'd175499: dataIn1 = 32'd8246
; 
32'd175500: dataIn1 = 32'd5213
; 
32'd175501: dataIn1 = 32'd6424
; 
32'd175502: dataIn1 = 32'd8156
; 
32'd175503: dataIn1 = 32'd8234
; 
32'd175504: dataIn1 = 32'd8239
; 
32'd175505: dataIn1 = 32'd8240
; 
32'd175506: dataIn1 = 32'd8243
; 
32'd175507: dataIn1 = 32'd6402
; 
32'd175508: dataIn1 = 32'd6414
; 
32'd175509: dataIn1 = 32'd8155
; 
32'd175510: dataIn1 = 32'd8188
; 
32'd175511: dataIn1 = 32'd8241
; 
32'd175512: dataIn1 = 32'd8242
; 
32'd175513: dataIn1 = 32'd8243
; 
32'd175514: dataIn1 = 32'd6414
; 
32'd175515: dataIn1 = 32'd6424
; 
32'd175516: dataIn1 = 32'd8190
; 
32'd175517: dataIn1 = 32'd8238
; 
32'd175518: dataIn1 = 32'd8241
; 
32'd175519: dataIn1 = 32'd8242
; 
32'd175520: dataIn1 = 32'd8243
; 
32'd175521: dataIn1 = 32'd6402
; 
32'd175522: dataIn1 = 32'd6424
; 
32'd175523: dataIn1 = 32'd8156
; 
32'd175524: dataIn1 = 32'd8240
; 
32'd175525: dataIn1 = 32'd8241
; 
32'd175526: dataIn1 = 32'd8242
; 
32'd175527: dataIn1 = 32'd8243
; 
32'd175528: dataIn1 = 32'd5010
; 
32'd175529: dataIn1 = 32'd6425
; 
32'd175530: dataIn1 = 32'd8236
; 
32'd175531: dataIn1 = 32'd8244
; 
32'd175532: dataIn1 = 32'd8245
; 
32'd175533: dataIn1 = 32'd8246
; 
32'd175534: dataIn1 = 32'd8247
; 
32'd175535: dataIn1 = 32'd5010
; 
32'd175536: dataIn1 = 32'd6403
; 
32'd175537: dataIn1 = 32'd8162
; 
32'd175538: dataIn1 = 32'd8244
; 
32'd175539: dataIn1 = 32'd8245
; 
32'd175540: dataIn1 = 32'd8246
; 
32'd175541: dataIn1 = 32'd8248
; 
32'd175542: dataIn1 = 32'd6403
; 
32'd175543: dataIn1 = 32'd6425
; 
32'd175544: dataIn1 = 32'd8163
; 
32'd175545: dataIn1 = 32'd8239
; 
32'd175546: dataIn1 = 32'd8244
; 
32'd175547: dataIn1 = 32'd8245
; 
32'd175548: dataIn1 = 32'd8246
; 
32'd175549: dataIn1 = 32'd2665
; 
32'd175550: dataIn1 = 32'd5007
; 
32'd175551: dataIn1 = 32'd5010
; 
32'd175552: dataIn1 = 32'd8236
; 
32'd175553: dataIn1 = 32'd8244
; 
32'd175554: dataIn1 = 32'd8247
; 
32'd175555: dataIn1 = 32'd142
; 
32'd175556: dataIn1 = 32'd4741
; 
32'd175557: dataIn1 = 32'd5010
; 
32'd175558: dataIn1 = 32'd8162
; 
32'd175559: dataIn1 = 32'd8245
; 
32'd175560: dataIn1 = 32'd8248
; 
32'd175561: dataIn1 = 32'd5011
; 
32'd175562: dataIn1 = 32'd6426
; 
32'd175563: dataIn1 = 32'd8235
; 
32'd175564: dataIn1 = 32'd8249
; 
32'd175565: dataIn1 = 32'd8250
; 
32'd175566: dataIn1 = 32'd8251
; 
32'd175567: dataIn1 = 32'd8252
; 
32'd175568: dataIn1 = 32'd6417
; 
32'd175569: dataIn1 = 32'd6426
; 
32'd175570: dataIn1 = 32'd8203
; 
32'd175571: dataIn1 = 32'd8237
; 
32'd175572: dataIn1 = 32'd8249
; 
32'd175573: dataIn1 = 32'd8250
; 
32'd175574: dataIn1 = 32'd8251
; 
32'd175575: dataIn1 = 32'd5011
; 
32'd175576: dataIn1 = 32'd6417
; 
32'd175577: dataIn1 = 32'd8205
; 
32'd175578: dataIn1 = 32'd8249
; 
32'd175579: dataIn1 = 32'd8250
; 
32'd175580: dataIn1 = 32'd8251
; 
32'd175581: dataIn1 = 32'd8253
; 
32'd175582: dataIn1 = 32'd2665
; 
32'd175583: dataIn1 = 32'd5009
; 
32'd175584: dataIn1 = 32'd5011
; 
32'd175585: dataIn1 = 32'd8235
; 
32'd175586: dataIn1 = 32'd8249
; 
32'd175587: dataIn1 = 32'd8252
; 
32'd175588: dataIn1 = 32'd1113
; 
32'd175589: dataIn1 = 32'd5006
; 
32'd175590: dataIn1 = 32'd5011
; 
32'd175591: dataIn1 = 32'd8205
; 
32'd175592: dataIn1 = 32'd8251
; 
32'd175593: dataIn1 = 32'd8253
; 
32'd175594: dataIn1 = 32'd6428
; 
32'd175595: dataIn1 = 32'd6429
; 
32'd175596: dataIn1 = 32'd8254
; 
32'd175597: dataIn1 = 32'd8255
; 
32'd175598: dataIn1 = 32'd8256
; 
32'd175599: dataIn1 = 32'd8257
; 
32'd175600: dataIn1 = 32'd8258
; 
32'd175601: dataIn1 = 32'd6427
; 
32'd175602: dataIn1 = 32'd6429
; 
32'd175603: dataIn1 = 32'd8254
; 
32'd175604: dataIn1 = 32'd8255
; 
32'd175605: dataIn1 = 32'd8256
; 
32'd175606: dataIn1 = 32'd8259
; 
32'd175607: dataIn1 = 32'd8260
; 
32'd175608: dataIn1 = 32'd6427
; 
32'd175609: dataIn1 = 32'd6428
; 
32'd175610: dataIn1 = 32'd8254
; 
32'd175611: dataIn1 = 32'd8255
; 
32'd175612: dataIn1 = 32'd8256
; 
32'd175613: dataIn1 = 32'd8261
; 
32'd175614: dataIn1 = 32'd8262
; 
32'd175615: dataIn1 = 32'd5220
; 
32'd175616: dataIn1 = 32'd6429
; 
32'd175617: dataIn1 = 32'd6765
; 
32'd175618: dataIn1 = 32'd8254
; 
32'd175619: dataIn1 = 32'd8257
; 
32'd175620: dataIn1 = 32'd8258
; 
32'd175621: dataIn1 = 32'd5220
; 
32'd175622: dataIn1 = 32'd6428
; 
32'd175623: dataIn1 = 32'd8254
; 
32'd175624: dataIn1 = 32'd8257
; 
32'd175625: dataIn1 = 32'd8258
; 
32'd175626: dataIn1 = 32'd8266
; 
32'd175627: dataIn1 = 32'd8269
; 
32'd175628: dataIn1 = 32'd5215
; 
32'd175629: dataIn1 = 32'd6429
; 
32'd175630: dataIn1 = 32'd6764
; 
32'd175631: dataIn1 = 32'd8255
; 
32'd175632: dataIn1 = 32'd8259
; 
32'd175633: dataIn1 = 32'd8260
; 
32'd175634: dataIn1 = 32'd5215
; 
32'd175635: dataIn1 = 32'd6427
; 
32'd175636: dataIn1 = 32'd8173
; 
32'd175637: dataIn1 = 32'd8255
; 
32'd175638: dataIn1 = 32'd8259
; 
32'd175639: dataIn1 = 32'd8260
; 
32'd175640: dataIn1 = 32'd8264
; 
32'd175641: dataIn1 = 32'd5218
; 
32'd175642: dataIn1 = 32'd6428
; 
32'd175643: dataIn1 = 32'd8198
; 
32'd175644: dataIn1 = 32'd8256
; 
32'd175645: dataIn1 = 32'd8261
; 
32'd175646: dataIn1 = 32'd8262
; 
32'd175647: dataIn1 = 32'd8268
; 
32'd175648: dataIn1 = 32'd5218
; 
32'd175649: dataIn1 = 32'd6427
; 
32'd175650: dataIn1 = 32'd8191
; 
32'd175651: dataIn1 = 32'd8256
; 
32'd175652: dataIn1 = 32'd8261
; 
32'd175653: dataIn1 = 32'd8262
; 
32'd175654: dataIn1 = 32'd8265
; 
32'd175655: dataIn1 = 32'd6407
; 
32'd175656: dataIn1 = 32'd6413
; 
32'd175657: dataIn1 = 32'd8172
; 
32'd175658: dataIn1 = 32'd8189
; 
32'd175659: dataIn1 = 32'd8263
; 
32'd175660: dataIn1 = 32'd8264
; 
32'd175661: dataIn1 = 32'd8265
; 
32'd175662: dataIn1 = 32'd6407
; 
32'd175663: dataIn1 = 32'd6427
; 
32'd175664: dataIn1 = 32'd8173
; 
32'd175665: dataIn1 = 32'd8260
; 
32'd175666: dataIn1 = 32'd8263
; 
32'd175667: dataIn1 = 32'd8264
; 
32'd175668: dataIn1 = 32'd8265
; 
32'd175669: dataIn1 = 32'd6413
; 
32'd175670: dataIn1 = 32'd6427
; 
32'd175671: dataIn1 = 32'd8191
; 
32'd175672: dataIn1 = 32'd8262
; 
32'd175673: dataIn1 = 32'd8263
; 
32'd175674: dataIn1 = 32'd8264
; 
32'd175675: dataIn1 = 32'd8265
; 
32'd175676: dataIn1 = 32'd6428
; 
32'd175677: dataIn1 = 32'd6430
; 
32'd175678: dataIn1 = 32'd8258
; 
32'd175679: dataIn1 = 32'd8266
; 
32'd175680: dataIn1 = 32'd8267
; 
32'd175681: dataIn1 = 32'd8268
; 
32'd175682: dataIn1 = 32'd8269
; 
32'd175683: dataIn1 = 32'd6415
; 
32'd175684: dataIn1 = 32'd6430
; 
32'd175685: dataIn1 = 32'd8197
; 
32'd175686: dataIn1 = 32'd8266
; 
32'd175687: dataIn1 = 32'd8267
; 
32'd175688: dataIn1 = 32'd8268
; 
32'd175689: dataIn1 = 32'd8270
; 
32'd175690: dataIn1 = 32'd6415
; 
32'd175691: dataIn1 = 32'd6428
; 
32'd175692: dataIn1 = 32'd8198
; 
32'd175693: dataIn1 = 32'd8261
; 
32'd175694: dataIn1 = 32'd8266
; 
32'd175695: dataIn1 = 32'd8267
; 
32'd175696: dataIn1 = 32'd8268
; 
32'd175697: dataIn1 = 32'd5220
; 
32'd175698: dataIn1 = 32'd6430
; 
32'd175699: dataIn1 = 32'd8258
; 
32'd175700: dataIn1 = 32'd8266
; 
32'd175701: dataIn1 = 32'd8269
; 
32'd175702: dataIn1 = 32'd9120
; 
32'd175703: dataIn1 = 32'd9123
; 
32'd175704: dataIn1 = 32'd2722
; 
32'd175705: dataIn1 = 32'd6430
; 
32'd175706: dataIn1 = 32'd8197
; 
32'd175707: dataIn1 = 32'd8267
; 
32'd175708: dataIn1 = 32'd8270
; 
32'd175709: dataIn1 = 32'd9101
; 
32'd175710: dataIn1 = 32'd9122
; 
32'd175711: dataIn1 = 32'd6432
; 
32'd175712: dataIn1 = 32'd6433
; 
32'd175713: dataIn1 = 32'd8271
; 
32'd175714: dataIn1 = 32'd8272
; 
32'd175715: dataIn1 = 32'd8273
; 
32'd175716: dataIn1 = 32'd8274
; 
32'd175717: dataIn1 = 32'd8275
; 
32'd175718: dataIn1 = 32'd6431
; 
32'd175719: dataIn1 = 32'd6433
; 
32'd175720: dataIn1 = 32'd8271
; 
32'd175721: dataIn1 = 32'd8272
; 
32'd175722: dataIn1 = 32'd8273
; 
32'd175723: dataIn1 = 32'd8276
; 
32'd175724: dataIn1 = 32'd8277
; 
32'd175725: dataIn1 = 32'd6431
; 
32'd175726: dataIn1 = 32'd6432
; 
32'd175727: dataIn1 = 32'd8271
; 
32'd175728: dataIn1 = 32'd8272
; 
32'd175729: dataIn1 = 32'd8273
; 
32'd175730: dataIn1 = 32'd8278
; 
32'd175731: dataIn1 = 32'd8279
; 
32'd175732: dataIn1 = 32'd5221
; 
32'd175733: dataIn1 = 32'd6433
; 
32'd175734: dataIn1 = 32'd8271
; 
32'd175735: dataIn1 = 32'd8274
; 
32'd175736: dataIn1 = 32'd8275
; 
32'd175737: dataIn1 = 32'd8294
; 
32'd175738: dataIn1 = 32'd8297
; 
32'd175739: dataIn1 = 32'd5221
; 
32'd175740: dataIn1 = 32'd6432
; 
32'd175741: dataIn1 = 32'd8271
; 
32'd175742: dataIn1 = 32'd8274
; 
32'd175743: dataIn1 = 32'd8275
; 
32'd175744: dataIn1 = 32'd8287
; 
32'd175745: dataIn1 = 32'd8290
; 
32'd175746: dataIn1 = 32'd5222
; 
32'd175747: dataIn1 = 32'd6433
; 
32'd175748: dataIn1 = 32'd8272
; 
32'd175749: dataIn1 = 32'd8276
; 
32'd175750: dataIn1 = 32'd8277
; 
32'd175751: dataIn1 = 32'd8295
; 
32'd175752: dataIn1 = 32'd8298
; 
32'd175753: dataIn1 = 32'd5222
; 
32'd175754: dataIn1 = 32'd6431
; 
32'd175755: dataIn1 = 32'd8272
; 
32'd175756: dataIn1 = 32'd8276
; 
32'd175757: dataIn1 = 32'd8277
; 
32'd175758: dataIn1 = 32'd8281
; 
32'd175759: dataIn1 = 32'd8285
; 
32'd175760: dataIn1 = 32'd5223
; 
32'd175761: dataIn1 = 32'd6432
; 
32'd175762: dataIn1 = 32'd8273
; 
32'd175763: dataIn1 = 32'd8278
; 
32'd175764: dataIn1 = 32'd8279
; 
32'd175765: dataIn1 = 32'd8289
; 
32'd175766: dataIn1 = 32'd8293
; 
32'd175767: dataIn1 = 32'd5223
; 
32'd175768: dataIn1 = 32'd6431
; 
32'd175769: dataIn1 = 32'd8273
; 
32'd175770: dataIn1 = 32'd8278
; 
32'd175771: dataIn1 = 32'd8279
; 
32'd175772: dataIn1 = 32'd8282
; 
32'd175773: dataIn1 = 32'd8286
; 
32'd175774: dataIn1 = 32'd6434
; 
32'd175775: dataIn1 = 32'd6435
; 
32'd175776: dataIn1 = 32'd8280
; 
32'd175777: dataIn1 = 32'd8281
; 
32'd175778: dataIn1 = 32'd8282
; 
32'd175779: dataIn1 = 32'd8283
; 
32'd175780: dataIn1 = 32'd8284
; 
32'd175781: dataIn1 = 32'd6431
; 
32'd175782: dataIn1 = 32'd6435
; 
32'd175783: dataIn1 = 32'd8277
; 
32'd175784: dataIn1 = 32'd8280
; 
32'd175785: dataIn1 = 32'd8281
; 
32'd175786: dataIn1 = 32'd8282
; 
32'd175787: dataIn1 = 32'd8285
; 
32'd175788: dataIn1 = 32'd6431
; 
32'd175789: dataIn1 = 32'd6434
; 
32'd175790: dataIn1 = 32'd8279
; 
32'd175791: dataIn1 = 32'd8280
; 
32'd175792: dataIn1 = 32'd8281
; 
32'd175793: dataIn1 = 32'd8282
; 
32'd175794: dataIn1 = 32'd8286
; 
32'd175795: dataIn1 = 32'd1114
; 
32'd175796: dataIn1 = 32'd6435
; 
32'd175797: dataIn1 = 32'd8280
; 
32'd175798: dataIn1 = 32'd8283
; 
32'd175799: dataIn1 = 32'd8284
; 
32'd175800: dataIn1 = 32'd8326
; 
32'd175801: dataIn1 = 32'd8329
; 
32'd175802: dataIn1 = 32'd1114
; 
32'd175803: dataIn1 = 32'd6434
; 
32'd175804: dataIn1 = 32'd8280
; 
32'd175805: dataIn1 = 32'd8283
; 
32'd175806: dataIn1 = 32'd8284
; 
32'd175807: dataIn1 = 32'd8348
; 
32'd175808: dataIn1 = 32'd8351
; 
32'd175809: dataIn1 = 32'd5222
; 
32'd175810: dataIn1 = 32'd6435
; 
32'd175811: dataIn1 = 32'd8277
; 
32'd175812: dataIn1 = 32'd8281
; 
32'd175813: dataIn1 = 32'd8285
; 
32'd175814: dataIn1 = 32'd8323
; 
32'd175815: dataIn1 = 32'd8327
; 
32'd175816: dataIn1 = 32'd5223
; 
32'd175817: dataIn1 = 32'd6434
; 
32'd175818: dataIn1 = 32'd8279
; 
32'd175819: dataIn1 = 32'd8282
; 
32'd175820: dataIn1 = 32'd8286
; 
32'd175821: dataIn1 = 32'd8347
; 
32'd175822: dataIn1 = 32'd8350
; 
32'd175823: dataIn1 = 32'd6432
; 
32'd175824: dataIn1 = 32'd6437
; 
32'd175825: dataIn1 = 32'd8275
; 
32'd175826: dataIn1 = 32'd8287
; 
32'd175827: dataIn1 = 32'd8288
; 
32'd175828: dataIn1 = 32'd8289
; 
32'd175829: dataIn1 = 32'd8290
; 
32'd175830: dataIn1 = 32'd6436
; 
32'd175831: dataIn1 = 32'd6437
; 
32'd175832: dataIn1 = 32'd8287
; 
32'd175833: dataIn1 = 32'd8288
; 
32'd175834: dataIn1 = 32'd8289
; 
32'd175835: dataIn1 = 32'd8291
; 
32'd175836: dataIn1 = 32'd8292
; 
32'd175837: dataIn1 = 32'd6432
; 
32'd175838: dataIn1 = 32'd6436
; 
32'd175839: dataIn1 = 32'd8278
; 
32'd175840: dataIn1 = 32'd8287
; 
32'd175841: dataIn1 = 32'd8288
; 
32'd175842: dataIn1 = 32'd8289
; 
32'd175843: dataIn1 = 32'd8293
; 
32'd175844: dataIn1 = 32'd5221
; 
32'd175845: dataIn1 = 32'd6437
; 
32'd175846: dataIn1 = 32'd8275
; 
32'd175847: dataIn1 = 32'd8287
; 
32'd175848: dataIn1 = 32'd8290
; 
32'd175849: dataIn1 = 32'd8305
; 
32'd175850: dataIn1 = 32'd8310
; 
32'd175851: dataIn1 = 32'd2723
; 
32'd175852: dataIn1 = 32'd6437
; 
32'd175853: dataIn1 = 32'd8288
; 
32'd175854: dataIn1 = 32'd8291
; 
32'd175855: dataIn1 = 32'd8292
; 
32'd175856: dataIn1 = 32'd8311
; 
32'd175857: dataIn1 = 32'd8313
; 
32'd175858: dataIn1 = 32'd2723
; 
32'd175859: dataIn1 = 32'd6436
; 
32'd175860: dataIn1 = 32'd8288
; 
32'd175861: dataIn1 = 32'd8291
; 
32'd175862: dataIn1 = 32'd8292
; 
32'd175863: dataIn1 = 32'd8354
; 
32'd175864: dataIn1 = 32'd8357
; 
32'd175865: dataIn1 = 32'd5223
; 
32'd175866: dataIn1 = 32'd6436
; 
32'd175867: dataIn1 = 32'd8278
; 
32'd175868: dataIn1 = 32'd8289
; 
32'd175869: dataIn1 = 32'd8293
; 
32'd175870: dataIn1 = 32'd8346
; 
32'd175871: dataIn1 = 32'd8355
; 
32'd175872: dataIn1 = 32'd6433
; 
32'd175873: dataIn1 = 32'd6439
; 
32'd175874: dataIn1 = 32'd8274
; 
32'd175875: dataIn1 = 32'd8294
; 
32'd175876: dataIn1 = 32'd8295
; 
32'd175877: dataIn1 = 32'd8296
; 
32'd175878: dataIn1 = 32'd8297
; 
32'd175879: dataIn1 = 32'd6433
; 
32'd175880: dataIn1 = 32'd6438
; 
32'd175881: dataIn1 = 32'd8276
; 
32'd175882: dataIn1 = 32'd8294
; 
32'd175883: dataIn1 = 32'd8295
; 
32'd175884: dataIn1 = 32'd8296
; 
32'd175885: dataIn1 = 32'd8298
; 
32'd175886: dataIn1 = 32'd6438
; 
32'd175887: dataIn1 = 32'd6439
; 
32'd175888: dataIn1 = 32'd8294
; 
32'd175889: dataIn1 = 32'd8295
; 
32'd175890: dataIn1 = 32'd8296
; 
32'd175891: dataIn1 = 32'd8299
; 
32'd175892: dataIn1 = 32'd8300
; 
32'd175893: dataIn1 = 32'd5221
; 
32'd175894: dataIn1 = 32'd6439
; 
32'd175895: dataIn1 = 32'd8274
; 
32'd175896: dataIn1 = 32'd8294
; 
32'd175897: dataIn1 = 32'd8297
; 
32'd175898: dataIn1 = 32'd8304
; 
32'd175899: dataIn1 = 32'd8314
; 
32'd175900: dataIn1 = 32'd5222
; 
32'd175901: dataIn1 = 32'd6438
; 
32'd175902: dataIn1 = 32'd8276
; 
32'd175903: dataIn1 = 32'd8295
; 
32'd175904: dataIn1 = 32'd8298
; 
32'd175905: dataIn1 = 32'd8322
; 
32'd175906: dataIn1 = 32'd8337
; 
32'd175907: dataIn1 = 32'd2721
; 
32'd175908: dataIn1 = 32'd6439
; 
32'd175909: dataIn1 = 32'd8142
; 
32'd175910: dataIn1 = 32'd8296
; 
32'd175911: dataIn1 = 32'd8299
; 
32'd175912: dataIn1 = 32'd8300
; 
32'd175913: dataIn1 = 32'd8316
; 
32'd175914: dataIn1 = 32'd2721
; 
32'd175915: dataIn1 = 32'd6438
; 
32'd175916: dataIn1 = 32'd8168
; 
32'd175917: dataIn1 = 32'd8296
; 
32'd175918: dataIn1 = 32'd8299
; 
32'd175919: dataIn1 = 32'd8300
; 
32'd175920: dataIn1 = 32'd8338
; 
32'd175921: dataIn1 = 32'd6441
; 
32'd175922: dataIn1 = 32'd6442
; 
32'd175923: dataIn1 = 32'd8301
; 
32'd175924: dataIn1 = 32'd8302
; 
32'd175925: dataIn1 = 32'd8303
; 
32'd175926: dataIn1 = 32'd8304
; 
32'd175927: dataIn1 = 32'd8305
; 
32'd175928: dataIn1 = 32'd6440
; 
32'd175929: dataIn1 = 32'd6442
; 
32'd175930: dataIn1 = 32'd8301
; 
32'd175931: dataIn1 = 32'd8302
; 
32'd175932: dataIn1 = 32'd8303
; 
32'd175933: dataIn1 = 32'd8306
; 
32'd175934: dataIn1 = 32'd8307
; 
32'd175935: dataIn1 = 32'd6440
; 
32'd175936: dataIn1 = 32'd6441
; 
32'd175937: dataIn1 = 32'd8301
; 
32'd175938: dataIn1 = 32'd8302
; 
32'd175939: dataIn1 = 32'd8303
; 
32'd175940: dataIn1 = 32'd8308
; 
32'd175941: dataIn1 = 32'd8309
; 
32'd175942: dataIn1 = 32'd5221
; 
32'd175943: dataIn1 = 32'd6442
; 
32'd175944: dataIn1 = 32'd8297
; 
32'd175945: dataIn1 = 32'd8301
; 
32'd175946: dataIn1 = 32'd8304
; 
32'd175947: dataIn1 = 32'd8305
; 
32'd175948: dataIn1 = 32'd8314
; 
32'd175949: dataIn1 = 32'd5221
; 
32'd175950: dataIn1 = 32'd6441
; 
32'd175951: dataIn1 = 32'd8290
; 
32'd175952: dataIn1 = 32'd8301
; 
32'd175953: dataIn1 = 32'd8304
; 
32'd175954: dataIn1 = 32'd8305
; 
32'd175955: dataIn1 = 32'd8310
; 
32'd175956: dataIn1 = 32'd5210
; 
32'd175957: dataIn1 = 32'd6442
; 
32'd175958: dataIn1 = 32'd8141
; 
32'd175959: dataIn1 = 32'd8302
; 
32'd175960: dataIn1 = 32'd8306
; 
32'd175961: dataIn1 = 32'd8307
; 
32'd175962: dataIn1 = 32'd8315
; 
32'd175963: dataIn1 = 32'd5210
; 
32'd175964: dataIn1 = 32'd6440
; 
32'd175965: dataIn1 = 32'd8302
; 
32'd175966: dataIn1 = 32'd8306
; 
32'd175967: dataIn1 = 32'd8307
; 
32'd175968: dataIn1 = 32'd10278
; 
32'd175969: dataIn1 = 32'd10280
; 
32'd175970: dataIn1 = 32'd5224
; 
32'd175971: dataIn1 = 32'd6441
; 
32'd175972: dataIn1 = 32'd8303
; 
32'd175973: dataIn1 = 32'd8308
; 
32'd175974: dataIn1 = 32'd8309
; 
32'd175975: dataIn1 = 32'd8312
; 
32'd175976: dataIn1 = 32'd9275
; 
32'd175977: dataIn1 = 32'd5224
; 
32'd175978: dataIn1 = 32'd6440
; 
32'd175979: dataIn1 = 32'd6443
; 
32'd175980: dataIn1 = 32'd8303
; 
32'd175981: dataIn1 = 32'd8308
; 
32'd175982: dataIn1 = 32'd8309
; 
32'd175983: dataIn1 = 32'd6437
; 
32'd175984: dataIn1 = 32'd6441
; 
32'd175985: dataIn1 = 32'd8290
; 
32'd175986: dataIn1 = 32'd8305
; 
32'd175987: dataIn1 = 32'd8310
; 
32'd175988: dataIn1 = 32'd8311
; 
32'd175989: dataIn1 = 32'd8312
; 
32'd175990: dataIn1 = 32'd6437
; 
32'd175991: dataIn1 = 32'd6444
; 
32'd175992: dataIn1 = 32'd8291
; 
32'd175993: dataIn1 = 32'd8310
; 
32'd175994: dataIn1 = 32'd8311
; 
32'd175995: dataIn1 = 32'd8312
; 
32'd175996: dataIn1 = 32'd8313
; 
32'd175997: dataIn1 = 32'd6441
; 
32'd175998: dataIn1 = 32'd6444
; 
32'd175999: dataIn1 = 32'd8308
; 
32'd176000: dataIn1 = 32'd8310
; 
32'd176001: dataIn1 = 32'd8311
; 
32'd176002: dataIn1 = 32'd8312
; 
32'd176003: dataIn1 = 32'd9275
; 
32'd176004: dataIn1 = 32'd2723
; 
32'd176005: dataIn1 = 32'd6444
; 
32'd176006: dataIn1 = 32'd8291
; 
32'd176007: dataIn1 = 32'd8311
; 
32'd176008: dataIn1 = 32'd8313
; 
32'd176009: dataIn1 = 32'd9145
; 
32'd176010: dataIn1 = 32'd9178
; 
32'd176011: dataIn1 = 32'd6439
; 
32'd176012: dataIn1 = 32'd6442
; 
32'd176013: dataIn1 = 32'd8297
; 
32'd176014: dataIn1 = 32'd8304
; 
32'd176015: dataIn1 = 32'd8314
; 
32'd176016: dataIn1 = 32'd8315
; 
32'd176017: dataIn1 = 32'd8316
; 
32'd176018: dataIn1 = 32'd6398
; 
32'd176019: dataIn1 = 32'd6442
; 
32'd176020: dataIn1 = 32'd8141
; 
32'd176021: dataIn1 = 32'd8306
; 
32'd176022: dataIn1 = 32'd8314
; 
32'd176023: dataIn1 = 32'd8315
; 
32'd176024: dataIn1 = 32'd8316
; 
32'd176025: dataIn1 = 32'd6398
; 
32'd176026: dataIn1 = 32'd6439
; 
32'd176027: dataIn1 = 32'd8142
; 
32'd176028: dataIn1 = 32'd8299
; 
32'd176029: dataIn1 = 32'd8314
; 
32'd176030: dataIn1 = 32'd8315
; 
32'd176031: dataIn1 = 32'd8316
; 
32'd176032: dataIn1 = 32'd6446
; 
32'd176033: dataIn1 = 32'd6447
; 
32'd176034: dataIn1 = 32'd8317
; 
32'd176035: dataIn1 = 32'd8318
; 
32'd176036: dataIn1 = 32'd8319
; 
32'd176037: dataIn1 = 32'd8320
; 
32'd176038: dataIn1 = 32'd8321
; 
32'd176039: dataIn1 = 32'd6445
; 
32'd176040: dataIn1 = 32'd6447
; 
32'd176041: dataIn1 = 32'd8317
; 
32'd176042: dataIn1 = 32'd8318
; 
32'd176043: dataIn1 = 32'd8319
; 
32'd176044: dataIn1 = 32'd8322
; 
32'd176045: dataIn1 = 32'd8323
; 
32'd176046: dataIn1 = 32'd6445
; 
32'd176047: dataIn1 = 32'd6446
; 
32'd176048: dataIn1 = 32'd8317
; 
32'd176049: dataIn1 = 32'd8318
; 
32'd176050: dataIn1 = 32'd8319
; 
32'd176051: dataIn1 = 32'd8324
; 
32'd176052: dataIn1 = 32'd8325
; 
32'd176053: dataIn1 = 32'd5212
; 
32'd176054: dataIn1 = 32'd6447
; 
32'd176055: dataIn1 = 32'd8167
; 
32'd176056: dataIn1 = 32'd8317
; 
32'd176057: dataIn1 = 32'd8320
; 
32'd176058: dataIn1 = 32'd8321
; 
32'd176059: dataIn1 = 32'd8336
; 
32'd176060: dataIn1 = 32'd5212
; 
32'd176061: dataIn1 = 32'd6446
; 
32'd176062: dataIn1 = 32'd8160
; 
32'd176063: dataIn1 = 32'd8317
; 
32'd176064: dataIn1 = 32'd8320
; 
32'd176065: dataIn1 = 32'd8321
; 
32'd176066: dataIn1 = 32'd8331
; 
32'd176067: dataIn1 = 32'd5222
; 
32'd176068: dataIn1 = 32'd6447
; 
32'd176069: dataIn1 = 32'd8298
; 
32'd176070: dataIn1 = 32'd8318
; 
32'd176071: dataIn1 = 32'd8322
; 
32'd176072: dataIn1 = 32'd8323
; 
32'd176073: dataIn1 = 32'd8337
; 
32'd176074: dataIn1 = 32'd5222
; 
32'd176075: dataIn1 = 32'd6445
; 
32'd176076: dataIn1 = 32'd8285
; 
32'd176077: dataIn1 = 32'd8318
; 
32'd176078: dataIn1 = 32'd8322
; 
32'd176079: dataIn1 = 32'd8323
; 
32'd176080: dataIn1 = 32'd8327
; 
32'd176081: dataIn1 = 32'd2670
; 
32'd176082: dataIn1 = 32'd6446
; 
32'd176083: dataIn1 = 32'd8319
; 
32'd176084: dataIn1 = 32'd8324
; 
32'd176085: dataIn1 = 32'd8325
; 
32'd176086: dataIn1 = 32'd8333
; 
32'd176087: dataIn1 = 32'd8335
; 
32'd176088: dataIn1 = 32'd2670
; 
32'd176089: dataIn1 = 32'd6445
; 
32'd176090: dataIn1 = 32'd8319
; 
32'd176091: dataIn1 = 32'd8324
; 
32'd176092: dataIn1 = 32'd8325
; 
32'd176093: dataIn1 = 32'd8328
; 
32'd176094: dataIn1 = 32'd8330
; 
32'd176095: dataIn1 = 32'd5030
; 
32'd176096: dataIn1 = 32'd6435
; 
32'd176097: dataIn1 = 32'd8283
; 
32'd176098: dataIn1 = 32'd8326
; 
32'd176099: dataIn1 = 32'd8327
; 
32'd176100: dataIn1 = 32'd8328
; 
32'd176101: dataIn1 = 32'd8329
; 
32'd176102: dataIn1 = 32'd6435
; 
32'd176103: dataIn1 = 32'd6445
; 
32'd176104: dataIn1 = 32'd8285
; 
32'd176105: dataIn1 = 32'd8323
; 
32'd176106: dataIn1 = 32'd8326
; 
32'd176107: dataIn1 = 32'd8327
; 
32'd176108: dataIn1 = 32'd8328
; 
32'd176109: dataIn1 = 32'd5030
; 
32'd176110: dataIn1 = 32'd6445
; 
32'd176111: dataIn1 = 32'd8325
; 
32'd176112: dataIn1 = 32'd8326
; 
32'd176113: dataIn1 = 32'd8327
; 
32'd176114: dataIn1 = 32'd8328
; 
32'd176115: dataIn1 = 32'd8330
; 
32'd176116: dataIn1 = 32'd1114
; 
32'd176117: dataIn1 = 32'd5023
; 
32'd176118: dataIn1 = 32'd5030
; 
32'd176119: dataIn1 = 32'd8283
; 
32'd176120: dataIn1 = 32'd8326
; 
32'd176121: dataIn1 = 32'd8329
; 
32'd176122: dataIn1 = 32'd2670
; 
32'd176123: dataIn1 = 32'd5027
; 
32'd176124: dataIn1 = 32'd5030
; 
32'd176125: dataIn1 = 32'd8325
; 
32'd176126: dataIn1 = 32'd8328
; 
32'd176127: dataIn1 = 32'd8330
; 
32'd176128: dataIn1 = 32'd6404
; 
32'd176129: dataIn1 = 32'd6446
; 
32'd176130: dataIn1 = 32'd8160
; 
32'd176131: dataIn1 = 32'd8321
; 
32'd176132: dataIn1 = 32'd8331
; 
32'd176133: dataIn1 = 32'd8332
; 
32'd176134: dataIn1 = 32'd8333
; 
32'd176135: dataIn1 = 32'd5029
; 
32'd176136: dataIn1 = 32'd6404
; 
32'd176137: dataIn1 = 32'd8161
; 
32'd176138: dataIn1 = 32'd8331
; 
32'd176139: dataIn1 = 32'd8332
; 
32'd176140: dataIn1 = 32'd8333
; 
32'd176141: dataIn1 = 32'd8334
; 
32'd176142: dataIn1 = 32'd5029
; 
32'd176143: dataIn1 = 32'd6446
; 
32'd176144: dataIn1 = 32'd8324
; 
32'd176145: dataIn1 = 32'd8331
; 
32'd176146: dataIn1 = 32'd8332
; 
32'd176147: dataIn1 = 32'd8333
; 
32'd176148: dataIn1 = 32'd8335
; 
32'd176149: dataIn1 = 32'd142
; 
32'd176150: dataIn1 = 32'd4742
; 
32'd176151: dataIn1 = 32'd5029
; 
32'd176152: dataIn1 = 32'd8161
; 
32'd176153: dataIn1 = 32'd8332
; 
32'd176154: dataIn1 = 32'd8334
; 
32'd176155: dataIn1 = 32'd2670
; 
32'd176156: dataIn1 = 32'd5026
; 
32'd176157: dataIn1 = 32'd5029
; 
32'd176158: dataIn1 = 32'd8324
; 
32'd176159: dataIn1 = 32'd8333
; 
32'd176160: dataIn1 = 32'd8335
; 
32'd176161: dataIn1 = 32'd6405
; 
32'd176162: dataIn1 = 32'd6447
; 
32'd176163: dataIn1 = 32'd8167
; 
32'd176164: dataIn1 = 32'd8320
; 
32'd176165: dataIn1 = 32'd8336
; 
32'd176166: dataIn1 = 32'd8337
; 
32'd176167: dataIn1 = 32'd8338
; 
32'd176168: dataIn1 = 32'd6438
; 
32'd176169: dataIn1 = 32'd6447
; 
32'd176170: dataIn1 = 32'd8298
; 
32'd176171: dataIn1 = 32'd8322
; 
32'd176172: dataIn1 = 32'd8336
; 
32'd176173: dataIn1 = 32'd8337
; 
32'd176174: dataIn1 = 32'd8338
; 
32'd176175: dataIn1 = 32'd6405
; 
32'd176176: dataIn1 = 32'd6438
; 
32'd176177: dataIn1 = 32'd8168
; 
32'd176178: dataIn1 = 32'd8300
; 
32'd176179: dataIn1 = 32'd8336
; 
32'd176180: dataIn1 = 32'd8337
; 
32'd176181: dataIn1 = 32'd8338
; 
32'd176182: dataIn1 = 32'd6449
; 
32'd176183: dataIn1 = 32'd6450
; 
32'd176184: dataIn1 = 32'd8339
; 
32'd176185: dataIn1 = 32'd8340
; 
32'd176186: dataIn1 = 32'd8341
; 
32'd176187: dataIn1 = 32'd8342
; 
32'd176188: dataIn1 = 32'd8343
; 
32'd176189: dataIn1 = 32'd6448
; 
32'd176190: dataIn1 = 32'd6450
; 
32'd176191: dataIn1 = 32'd8339
; 
32'd176192: dataIn1 = 32'd8340
; 
32'd176193: dataIn1 = 32'd8341
; 
32'd176194: dataIn1 = 32'd8344
; 
32'd176195: dataIn1 = 32'd8345
; 
32'd176196: dataIn1 = 32'd6448
; 
32'd176197: dataIn1 = 32'd6449
; 
32'd176198: dataIn1 = 32'd8339
; 
32'd176199: dataIn1 = 32'd8340
; 
32'd176200: dataIn1 = 32'd8341
; 
32'd176201: dataIn1 = 32'd8346
; 
32'd176202: dataIn1 = 32'd8347
; 
32'd176203: dataIn1 = 32'd5225
; 
32'd176204: dataIn1 = 32'd6450
; 
32'd176205: dataIn1 = 32'd8339
; 
32'd176206: dataIn1 = 32'd8342
; 
32'd176207: dataIn1 = 32'd8343
; 
32'd176208: dataIn1 = 32'd8358
; 
32'd176209: dataIn1 = 32'd8361
; 
32'd176210: dataIn1 = 32'd5225
; 
32'd176211: dataIn1 = 32'd6449
; 
32'd176212: dataIn1 = 32'd8339
; 
32'd176213: dataIn1 = 32'd8342
; 
32'd176214: dataIn1 = 32'd8343
; 
32'd176215: dataIn1 = 32'd8353
; 
32'd176216: dataIn1 = 32'd8356
; 
32'd176217: dataIn1 = 32'd2671
; 
32'd176218: dataIn1 = 32'd6450
; 
32'd176219: dataIn1 = 32'd8340
; 
32'd176220: dataIn1 = 32'd8344
; 
32'd176221: dataIn1 = 32'd8345
; 
32'd176222: dataIn1 = 32'd8359
; 
32'd176223: dataIn1 = 32'd8362
; 
32'd176224: dataIn1 = 32'd2671
; 
32'd176225: dataIn1 = 32'd6448
; 
32'd176226: dataIn1 = 32'd8340
; 
32'd176227: dataIn1 = 32'd8344
; 
32'd176228: dataIn1 = 32'd8345
; 
32'd176229: dataIn1 = 32'd8349
; 
32'd176230: dataIn1 = 32'd8352
; 
32'd176231: dataIn1 = 32'd5223
; 
32'd176232: dataIn1 = 32'd6449
; 
32'd176233: dataIn1 = 32'd8293
; 
32'd176234: dataIn1 = 32'd8341
; 
32'd176235: dataIn1 = 32'd8346
; 
32'd176236: dataIn1 = 32'd8347
; 
32'd176237: dataIn1 = 32'd8355
; 
32'd176238: dataIn1 = 32'd5223
; 
32'd176239: dataIn1 = 32'd6448
; 
32'd176240: dataIn1 = 32'd8286
; 
32'd176241: dataIn1 = 32'd8341
; 
32'd176242: dataIn1 = 32'd8346
; 
32'd176243: dataIn1 = 32'd8347
; 
32'd176244: dataIn1 = 32'd8350
; 
32'd176245: dataIn1 = 32'd5034
; 
32'd176246: dataIn1 = 32'd6434
; 
32'd176247: dataIn1 = 32'd8284
; 
32'd176248: dataIn1 = 32'd8348
; 
32'd176249: dataIn1 = 32'd8349
; 
32'd176250: dataIn1 = 32'd8350
; 
32'd176251: dataIn1 = 32'd8351
; 
32'd176252: dataIn1 = 32'd5034
; 
32'd176253: dataIn1 = 32'd6448
; 
32'd176254: dataIn1 = 32'd8345
; 
32'd176255: dataIn1 = 32'd8348
; 
32'd176256: dataIn1 = 32'd8349
; 
32'd176257: dataIn1 = 32'd8350
; 
32'd176258: dataIn1 = 32'd8352
; 
32'd176259: dataIn1 = 32'd6434
; 
32'd176260: dataIn1 = 32'd6448
; 
32'd176261: dataIn1 = 32'd8286
; 
32'd176262: dataIn1 = 32'd8347
; 
32'd176263: dataIn1 = 32'd8348
; 
32'd176264: dataIn1 = 32'd8349
; 
32'd176265: dataIn1 = 32'd8350
; 
32'd176266: dataIn1 = 32'd1114
; 
32'd176267: dataIn1 = 32'd5022
; 
32'd176268: dataIn1 = 32'd5034
; 
32'd176269: dataIn1 = 32'd8284
; 
32'd176270: dataIn1 = 32'd8348
; 
32'd176271: dataIn1 = 32'd8351
; 
32'd176272: dataIn1 = 32'd2671
; 
32'd176273: dataIn1 = 32'd5032
; 
32'd176274: dataIn1 = 32'd5034
; 
32'd176275: dataIn1 = 32'd8345
; 
32'd176276: dataIn1 = 32'd8349
; 
32'd176277: dataIn1 = 32'd8352
; 
32'd176278: dataIn1 = 32'd6449
; 
32'd176279: dataIn1 = 32'd6451
; 
32'd176280: dataIn1 = 32'd8343
; 
32'd176281: dataIn1 = 32'd8353
; 
32'd176282: dataIn1 = 32'd8354
; 
32'd176283: dataIn1 = 32'd8355
; 
32'd176284: dataIn1 = 32'd8356
; 
32'd176285: dataIn1 = 32'd6436
; 
32'd176286: dataIn1 = 32'd6451
; 
32'd176287: dataIn1 = 32'd8292
; 
32'd176288: dataIn1 = 32'd8353
; 
32'd176289: dataIn1 = 32'd8354
; 
32'd176290: dataIn1 = 32'd8355
; 
32'd176291: dataIn1 = 32'd8357
; 
32'd176292: dataIn1 = 32'd6436
; 
32'd176293: dataIn1 = 32'd6449
; 
32'd176294: dataIn1 = 32'd8293
; 
32'd176295: dataIn1 = 32'd8346
; 
32'd176296: dataIn1 = 32'd8353
; 
32'd176297: dataIn1 = 32'd8354
; 
32'd176298: dataIn1 = 32'd8355
; 
32'd176299: dataIn1 = 32'd5225
; 
32'd176300: dataIn1 = 32'd6451
; 
32'd176301: dataIn1 = 32'd8343
; 
32'd176302: dataIn1 = 32'd8353
; 
32'd176303: dataIn1 = 32'd8356
; 
32'd176304: dataIn1 = 32'd9161
; 
32'd176305: dataIn1 = 32'd9168
; 
32'd176306: dataIn1 = 32'd2723
; 
32'd176307: dataIn1 = 32'd6451
; 
32'd176308: dataIn1 = 32'd8292
; 
32'd176309: dataIn1 = 32'd8354
; 
32'd176310: dataIn1 = 32'd8357
; 
32'd176311: dataIn1 = 32'd9144
; 
32'd176312: dataIn1 = 32'd9167
; 
32'd176313: dataIn1 = 32'd6450
; 
32'd176314: dataIn1 = 32'd6452
; 
32'd176315: dataIn1 = 32'd8342
; 
32'd176316: dataIn1 = 32'd8358
; 
32'd176317: dataIn1 = 32'd8359
; 
32'd176318: dataIn1 = 32'd8360
; 
32'd176319: dataIn1 = 32'd8361
; 
32'd176320: dataIn1 = 32'd5035
; 
32'd176321: dataIn1 = 32'd6450
; 
32'd176322: dataIn1 = 32'd8344
; 
32'd176323: dataIn1 = 32'd8358
; 
32'd176324: dataIn1 = 32'd8359
; 
32'd176325: dataIn1 = 32'd8360
; 
32'd176326: dataIn1 = 32'd8362
; 
32'd176327: dataIn1 = 32'd5035
; 
32'd176328: dataIn1 = 32'd6452
; 
32'd176329: dataIn1 = 32'd8358
; 
32'd176330: dataIn1 = 32'd8359
; 
32'd176331: dataIn1 = 32'd8360
; 
32'd176332: dataIn1 = 32'd8363
; 
32'd176333: dataIn1 = 32'd8364
; 
32'd176334: dataIn1 = 32'd5225
; 
32'd176335: dataIn1 = 32'd6452
; 
32'd176336: dataIn1 = 32'd8342
; 
32'd176337: dataIn1 = 32'd8358
; 
32'd176338: dataIn1 = 32'd8361
; 
32'd176339: dataIn1 = 32'd9162
; 
32'd176340: dataIn1 = 32'd9165
; 
32'd176341: dataIn1 = 32'd2671
; 
32'd176342: dataIn1 = 32'd5033
; 
32'd176343: dataIn1 = 32'd5035
; 
32'd176344: dataIn1 = 32'd8344
; 
32'd176345: dataIn1 = 32'd8359
; 
32'd176346: dataIn1 = 32'd8362
; 
32'd176347: dataIn1 = 32'd10
; 
32'd176348: dataIn1 = 32'd6452
; 
32'd176349: dataIn1 = 32'd8360
; 
32'd176350: dataIn1 = 32'd8363
; 
32'd176351: dataIn1 = 32'd8364
; 
32'd176352: dataIn1 = 32'd8471
; 
32'd176353: dataIn1 = 32'd9163
; 
32'd176354: dataIn1 = 32'd10
; 
32'd176355: dataIn1 = 32'd4752
; 
32'd176356: dataIn1 = 32'd5035
; 
32'd176357: dataIn1 = 32'd8360
; 
32'd176358: dataIn1 = 32'd8363
; 
32'd176359: dataIn1 = 32'd8364
; 
32'd176360: dataIn1 = 32'd6454
; 
32'd176361: dataIn1 = 32'd6455
; 
32'd176362: dataIn1 = 32'd8365
; 
32'd176363: dataIn1 = 32'd8366
; 
32'd176364: dataIn1 = 32'd8367
; 
32'd176365: dataIn1 = 32'd8368
; 
32'd176366: dataIn1 = 32'd8369
; 
32'd176367: dataIn1 = 32'd6453
; 
32'd176368: dataIn1 = 32'd6455
; 
32'd176369: dataIn1 = 32'd8365
; 
32'd176370: dataIn1 = 32'd8366
; 
32'd176371: dataIn1 = 32'd8367
; 
32'd176372: dataIn1 = 32'd8370
; 
32'd176373: dataIn1 = 32'd8371
; 
32'd176374: dataIn1 = 32'd6453
; 
32'd176375: dataIn1 = 32'd6454
; 
32'd176376: dataIn1 = 32'd8365
; 
32'd176377: dataIn1 = 32'd8366
; 
32'd176378: dataIn1 = 32'd8367
; 
32'd176379: dataIn1 = 32'd8372
; 
32'd176380: dataIn1 = 32'd8373
; 
32'd176381: dataIn1 = 32'd5226
; 
32'd176382: dataIn1 = 32'd6455
; 
32'd176383: dataIn1 = 32'd8365
; 
32'd176384: dataIn1 = 32'd8368
; 
32'd176385: dataIn1 = 32'd8369
; 
32'd176386: dataIn1 = 32'd8381
; 
32'd176387: dataIn1 = 32'd8384
; 
32'd176388: dataIn1 = 32'd5226
; 
32'd176389: dataIn1 = 32'd6454
; 
32'd176390: dataIn1 = 32'd6767
; 
32'd176391: dataIn1 = 32'd8365
; 
32'd176392: dataIn1 = 32'd8368
; 
32'd176393: dataIn1 = 32'd8369
; 
32'd176394: dataIn1 = 32'd5227
; 
32'd176395: dataIn1 = 32'd6455
; 
32'd176396: dataIn1 = 32'd8366
; 
32'd176397: dataIn1 = 32'd8370
; 
32'd176398: dataIn1 = 32'd8371
; 
32'd176399: dataIn1 = 32'd8382
; 
32'd176400: dataIn1 = 32'd8385
; 
32'd176401: dataIn1 = 32'd5227
; 
32'd176402: dataIn1 = 32'd6453
; 
32'd176403: dataIn1 = 32'd8366
; 
32'd176404: dataIn1 = 32'd8370
; 
32'd176405: dataIn1 = 32'd8371
; 
32'd176406: dataIn1 = 32'd8375
; 
32'd176407: dataIn1 = 32'd8379
; 
32'd176408: dataIn1 = 32'd5228
; 
32'd176409: dataIn1 = 32'd6454
; 
32'd176410: dataIn1 = 32'd6766
; 
32'd176411: dataIn1 = 32'd8367
; 
32'd176412: dataIn1 = 32'd8372
; 
32'd176413: dataIn1 = 32'd8373
; 
32'd176414: dataIn1 = 32'd5228
; 
32'd176415: dataIn1 = 32'd6453
; 
32'd176416: dataIn1 = 32'd8367
; 
32'd176417: dataIn1 = 32'd8372
; 
32'd176418: dataIn1 = 32'd8373
; 
32'd176419: dataIn1 = 32'd8376
; 
32'd176420: dataIn1 = 32'd8380
; 
32'd176421: dataIn1 = 32'd6456
; 
32'd176422: dataIn1 = 32'd6457
; 
32'd176423: dataIn1 = 32'd8374
; 
32'd176424: dataIn1 = 32'd8375
; 
32'd176425: dataIn1 = 32'd8376
; 
32'd176426: dataIn1 = 32'd8377
; 
32'd176427: dataIn1 = 32'd8378
; 
32'd176428: dataIn1 = 32'd6453
; 
32'd176429: dataIn1 = 32'd6457
; 
32'd176430: dataIn1 = 32'd8371
; 
32'd176431: dataIn1 = 32'd8374
; 
32'd176432: dataIn1 = 32'd8375
; 
32'd176433: dataIn1 = 32'd8376
; 
32'd176434: dataIn1 = 32'd8379
; 
32'd176435: dataIn1 = 32'd6453
; 
32'd176436: dataIn1 = 32'd6456
; 
32'd176437: dataIn1 = 32'd8373
; 
32'd176438: dataIn1 = 32'd8374
; 
32'd176439: dataIn1 = 32'd8375
; 
32'd176440: dataIn1 = 32'd8376
; 
32'd176441: dataIn1 = 32'd8380
; 
32'd176442: dataIn1 = 32'd2724
; 
32'd176443: dataIn1 = 32'd6457
; 
32'd176444: dataIn1 = 32'd8374
; 
32'd176445: dataIn1 = 32'd8377
; 
32'd176446: dataIn1 = 32'd8378
; 
32'd176447: dataIn1 = 32'd8404
; 
32'd176448: dataIn1 = 32'd8407
; 
32'd176449: dataIn1 = 32'd2724
; 
32'd176450: dataIn1 = 32'd6456
; 
32'd176451: dataIn1 = 32'd8374
; 
32'd176452: dataIn1 = 32'd8377
; 
32'd176453: dataIn1 = 32'd8378
; 
32'd176454: dataIn1 = 32'd8421
; 
32'd176455: dataIn1 = 32'd8424
; 
32'd176456: dataIn1 = 32'd5227
; 
32'd176457: dataIn1 = 32'd6457
; 
32'd176458: dataIn1 = 32'd8371
; 
32'd176459: dataIn1 = 32'd8375
; 
32'd176460: dataIn1 = 32'd8379
; 
32'd176461: dataIn1 = 32'd8401
; 
32'd176462: dataIn1 = 32'd8405
; 
32'd176463: dataIn1 = 32'd5228
; 
32'd176464: dataIn1 = 32'd6456
; 
32'd176465: dataIn1 = 32'd8373
; 
32'd176466: dataIn1 = 32'd8376
; 
32'd176467: dataIn1 = 32'd8380
; 
32'd176468: dataIn1 = 32'd8423
; 
32'd176469: dataIn1 = 32'd8427
; 
32'd176470: dataIn1 = 32'd6455
; 
32'd176471: dataIn1 = 32'd6459
; 
32'd176472: dataIn1 = 32'd8368
; 
32'd176473: dataIn1 = 32'd8381
; 
32'd176474: dataIn1 = 32'd8382
; 
32'd176475: dataIn1 = 32'd8383
; 
32'd176476: dataIn1 = 32'd8384
; 
32'd176477: dataIn1 = 32'd6455
; 
32'd176478: dataIn1 = 32'd6458
; 
32'd176479: dataIn1 = 32'd8370
; 
32'd176480: dataIn1 = 32'd8381
; 
32'd176481: dataIn1 = 32'd8382
; 
32'd176482: dataIn1 = 32'd8383
; 
32'd176483: dataIn1 = 32'd8385
; 
32'd176484: dataIn1 = 32'd6458
; 
32'd176485: dataIn1 = 32'd6459
; 
32'd176486: dataIn1 = 32'd8381
; 
32'd176487: dataIn1 = 32'd8382
; 
32'd176488: dataIn1 = 32'd8383
; 
32'd176489: dataIn1 = 32'd8386
; 
32'd176490: dataIn1 = 32'd8387
; 
32'd176491: dataIn1 = 32'd5226
; 
32'd176492: dataIn1 = 32'd6459
; 
32'd176493: dataIn1 = 32'd8368
; 
32'd176494: dataIn1 = 32'd8381
; 
32'd176495: dataIn1 = 32'd8384
; 
32'd176496: dataIn1 = 32'd8388
; 
32'd176497: dataIn1 = 32'd8391
; 
32'd176498: dataIn1 = 32'd5227
; 
32'd176499: dataIn1 = 32'd6458
; 
32'd176500: dataIn1 = 32'd8370
; 
32'd176501: dataIn1 = 32'd8382
; 
32'd176502: dataIn1 = 32'd8385
; 
32'd176503: dataIn1 = 32'd8400
; 
32'd176504: dataIn1 = 32'd8417
; 
32'd176505: dataIn1 = 32'd2726
; 
32'd176506: dataIn1 = 32'd6459
; 
32'd176507: dataIn1 = 32'd8383
; 
32'd176508: dataIn1 = 32'd8386
; 
32'd176509: dataIn1 = 32'd8387
; 
32'd176510: dataIn1 = 32'd8390
; 
32'd176511: dataIn1 = 32'd8394
; 
32'd176512: dataIn1 = 32'd2726
; 
32'd176513: dataIn1 = 32'd6458
; 
32'd176514: dataIn1 = 32'd8383
; 
32'd176515: dataIn1 = 32'd8386
; 
32'd176516: dataIn1 = 32'd8387
; 
32'd176517: dataIn1 = 32'd8418
; 
32'd176518: dataIn1 = 32'd8420
; 
32'd176519: dataIn1 = 32'd6459
; 
32'd176520: dataIn1 = 32'd6461
; 
32'd176521: dataIn1 = 32'd8384
; 
32'd176522: dataIn1 = 32'd8388
; 
32'd176523: dataIn1 = 32'd8389
; 
32'd176524: dataIn1 = 32'd8390
; 
32'd176525: dataIn1 = 32'd8391
; 
32'd176526: dataIn1 = 32'd6460
; 
32'd176527: dataIn1 = 32'd6461
; 
32'd176528: dataIn1 = 32'd8388
; 
32'd176529: dataIn1 = 32'd8389
; 
32'd176530: dataIn1 = 32'd8390
; 
32'd176531: dataIn1 = 32'd8392
; 
32'd176532: dataIn1 = 32'd8393
; 
32'd176533: dataIn1 = 32'd6459
; 
32'd176534: dataIn1 = 32'd6460
; 
32'd176535: dataIn1 = 32'd8386
; 
32'd176536: dataIn1 = 32'd8388
; 
32'd176537: dataIn1 = 32'd8389
; 
32'd176538: dataIn1 = 32'd8390
; 
32'd176539: dataIn1 = 32'd8394
; 
32'd176540: dataIn1 = 32'd5226
; 
32'd176541: dataIn1 = 32'd6461
; 
32'd176542: dataIn1 = 32'd6769
; 
32'd176543: dataIn1 = 32'd8384
; 
32'd176544: dataIn1 = 32'd8388
; 
32'd176545: dataIn1 = 32'd8391
; 
32'd176546: dataIn1 = 32'd5229
; 
32'd176547: dataIn1 = 32'd6461
; 
32'd176548: dataIn1 = 32'd6768
; 
32'd176549: dataIn1 = 32'd8389
; 
32'd176550: dataIn1 = 32'd8392
; 
32'd176551: dataIn1 = 32'd8393
; 
32'd176552: dataIn1 = 32'd5229
; 
32'd176553: dataIn1 = 32'd6460
; 
32'd176554: dataIn1 = 32'd8389
; 
32'd176555: dataIn1 = 32'd8392
; 
32'd176556: dataIn1 = 32'd8393
; 
32'd176557: dataIn1 = 32'd8558
; 
32'd176558: dataIn1 = 32'd8568
; 
32'd176559: dataIn1 = 32'd2726
; 
32'd176560: dataIn1 = 32'd6460
; 
32'd176561: dataIn1 = 32'd8386
; 
32'd176562: dataIn1 = 32'd8390
; 
32'd176563: dataIn1 = 32'd8394
; 
32'd176564: dataIn1 = 32'd8551
; 
32'd176565: dataIn1 = 32'd8569
; 
32'd176566: dataIn1 = 32'd6463
; 
32'd176567: dataIn1 = 32'd6464
; 
32'd176568: dataIn1 = 32'd8395
; 
32'd176569: dataIn1 = 32'd8396
; 
32'd176570: dataIn1 = 32'd8397
; 
32'd176571: dataIn1 = 32'd8398
; 
32'd176572: dataIn1 = 32'd8399
; 
32'd176573: dataIn1 = 32'd6462
; 
32'd176574: dataIn1 = 32'd6464
; 
32'd176575: dataIn1 = 32'd8395
; 
32'd176576: dataIn1 = 32'd8396
; 
32'd176577: dataIn1 = 32'd8397
; 
32'd176578: dataIn1 = 32'd8400
; 
32'd176579: dataIn1 = 32'd8401
; 
32'd176580: dataIn1 = 32'd6462
; 
32'd176581: dataIn1 = 32'd6463
; 
32'd176582: dataIn1 = 32'd8395
; 
32'd176583: dataIn1 = 32'd8396
; 
32'd176584: dataIn1 = 32'd8397
; 
32'd176585: dataIn1 = 32'd8402
; 
32'd176586: dataIn1 = 32'd8403
; 
32'd176587: dataIn1 = 32'd5231
; 
32'd176588: dataIn1 = 32'd6464
; 
32'd176589: dataIn1 = 32'd8395
; 
32'd176590: dataIn1 = 32'd8398
; 
32'd176591: dataIn1 = 32'd8399
; 
32'd176592: dataIn1 = 32'd8416
; 
32'd176593: dataIn1 = 32'd8419
; 
32'd176594: dataIn1 = 32'd5231
; 
32'd176595: dataIn1 = 32'd6463
; 
32'd176596: dataIn1 = 32'd8395
; 
32'd176597: dataIn1 = 32'd8398
; 
32'd176598: dataIn1 = 32'd8399
; 
32'd176599: dataIn1 = 32'd8409
; 
32'd176600: dataIn1 = 32'd8412
; 
32'd176601: dataIn1 = 32'd5227
; 
32'd176602: dataIn1 = 32'd6464
; 
32'd176603: dataIn1 = 32'd8385
; 
32'd176604: dataIn1 = 32'd8396
; 
32'd176605: dataIn1 = 32'd8400
; 
32'd176606: dataIn1 = 32'd8401
; 
32'd176607: dataIn1 = 32'd8417
; 
32'd176608: dataIn1 = 32'd5227
; 
32'd176609: dataIn1 = 32'd6462
; 
32'd176610: dataIn1 = 32'd8379
; 
32'd176611: dataIn1 = 32'd8396
; 
32'd176612: dataIn1 = 32'd8400
; 
32'd176613: dataIn1 = 32'd8401
; 
32'd176614: dataIn1 = 32'd8405
; 
32'd176615: dataIn1 = 32'd5232
; 
32'd176616: dataIn1 = 32'd6463
; 
32'd176617: dataIn1 = 32'd8397
; 
32'd176618: dataIn1 = 32'd8402
; 
32'd176619: dataIn1 = 32'd8403
; 
32'd176620: dataIn1 = 32'd8411
; 
32'd176621: dataIn1 = 32'd8415
; 
32'd176622: dataIn1 = 32'd5232
; 
32'd176623: dataIn1 = 32'd6462
; 
32'd176624: dataIn1 = 32'd8397
; 
32'd176625: dataIn1 = 32'd8402
; 
32'd176626: dataIn1 = 32'd8403
; 
32'd176627: dataIn1 = 32'd8406
; 
32'd176628: dataIn1 = 32'd8408
; 
32'd176629: dataIn1 = 32'd6457
; 
32'd176630: dataIn1 = 32'd6465
; 
32'd176631: dataIn1 = 32'd8377
; 
32'd176632: dataIn1 = 32'd8404
; 
32'd176633: dataIn1 = 32'd8405
; 
32'd176634: dataIn1 = 32'd8406
; 
32'd176635: dataIn1 = 32'd8407
; 
32'd176636: dataIn1 = 32'd6457
; 
32'd176637: dataIn1 = 32'd6462
; 
32'd176638: dataIn1 = 32'd8379
; 
32'd176639: dataIn1 = 32'd8401
; 
32'd176640: dataIn1 = 32'd8404
; 
32'd176641: dataIn1 = 32'd8405
; 
32'd176642: dataIn1 = 32'd8406
; 
32'd176643: dataIn1 = 32'd6462
; 
32'd176644: dataIn1 = 32'd6465
; 
32'd176645: dataIn1 = 32'd8403
; 
32'd176646: dataIn1 = 32'd8404
; 
32'd176647: dataIn1 = 32'd8405
; 
32'd176648: dataIn1 = 32'd8406
; 
32'd176649: dataIn1 = 32'd8408
; 
32'd176650: dataIn1 = 32'd2724
; 
32'd176651: dataIn1 = 32'd6465
; 
32'd176652: dataIn1 = 32'd8377
; 
32'd176653: dataIn1 = 32'd8404
; 
32'd176654: dataIn1 = 32'd8407
; 
32'd176655: dataIn1 = 32'd8440
; 
32'd176656: dataIn1 = 32'd8493
; 
32'd176657: dataIn1 = 32'd5232
; 
32'd176658: dataIn1 = 32'd6465
; 
32'd176659: dataIn1 = 32'd8403
; 
32'd176660: dataIn1 = 32'd8406
; 
32'd176661: dataIn1 = 32'd8408
; 
32'd176662: dataIn1 = 32'd8492
; 
32'd176663: dataIn1 = 32'd8495
; 
32'd176664: dataIn1 = 32'd6463
; 
32'd176665: dataIn1 = 32'd6467
; 
32'd176666: dataIn1 = 32'd8399
; 
32'd176667: dataIn1 = 32'd8409
; 
32'd176668: dataIn1 = 32'd8410
; 
32'd176669: dataIn1 = 32'd8411
; 
32'd176670: dataIn1 = 32'd8412
; 
32'd176671: dataIn1 = 32'd6466
; 
32'd176672: dataIn1 = 32'd6467
; 
32'd176673: dataIn1 = 32'd8409
; 
32'd176674: dataIn1 = 32'd8410
; 
32'd176675: dataIn1 = 32'd8411
; 
32'd176676: dataIn1 = 32'd8413
; 
32'd176677: dataIn1 = 32'd8414
; 
32'd176678: dataIn1 = 32'd6463
; 
32'd176679: dataIn1 = 32'd6466
; 
32'd176680: dataIn1 = 32'd8402
; 
32'd176681: dataIn1 = 32'd8409
; 
32'd176682: dataIn1 = 32'd8410
; 
32'd176683: dataIn1 = 32'd8411
; 
32'd176684: dataIn1 = 32'd8415
; 
32'd176685: dataIn1 = 32'd5231
; 
32'd176686: dataIn1 = 32'd6467
; 
32'd176687: dataIn1 = 32'd8399
; 
32'd176688: dataIn1 = 32'd8409
; 
32'd176689: dataIn1 = 32'd8412
; 
32'd176690: dataIn1 = 32'd8574
; 
32'd176691: dataIn1 = 32'd8584
; 
32'd176692: dataIn1 = 32'd145
; 
32'd176693: dataIn1 = 32'd6467
; 
32'd176694: dataIn1 = 32'd8410
; 
32'd176695: dataIn1 = 32'd8413
; 
32'd176696: dataIn1 = 32'd8414
; 
32'd176697: dataIn1 = 32'd8585
; 
32'd176698: dataIn1 = 32'd8587
; 
32'd176699: dataIn1 = 32'd145
; 
32'd176700: dataIn1 = 32'd6466
; 
32'd176701: dataIn1 = 32'd8410
; 
32'd176702: dataIn1 = 32'd8413
; 
32'd176703: dataIn1 = 32'd8414
; 
32'd176704: dataIn1 = 32'd8497
; 
32'd176705: dataIn1 = 32'd8500
; 
32'd176706: dataIn1 = 32'd5232
; 
32'd176707: dataIn1 = 32'd6466
; 
32'd176708: dataIn1 = 32'd8402
; 
32'd176709: dataIn1 = 32'd8411
; 
32'd176710: dataIn1 = 32'd8415
; 
32'd176711: dataIn1 = 32'd8491
; 
32'd176712: dataIn1 = 32'd8498
; 
32'd176713: dataIn1 = 32'd6464
; 
32'd176714: dataIn1 = 32'd6468
; 
32'd176715: dataIn1 = 32'd8398
; 
32'd176716: dataIn1 = 32'd8416
; 
32'd176717: dataIn1 = 32'd8417
; 
32'd176718: dataIn1 = 32'd8418
; 
32'd176719: dataIn1 = 32'd8419
; 
32'd176720: dataIn1 = 32'd6458
; 
32'd176721: dataIn1 = 32'd6464
; 
32'd176722: dataIn1 = 32'd8385
; 
32'd176723: dataIn1 = 32'd8400
; 
32'd176724: dataIn1 = 32'd8416
; 
32'd176725: dataIn1 = 32'd8417
; 
32'd176726: dataIn1 = 32'd8418
; 
32'd176727: dataIn1 = 32'd6458
; 
32'd176728: dataIn1 = 32'd6468
; 
32'd176729: dataIn1 = 32'd8387
; 
32'd176730: dataIn1 = 32'd8416
; 
32'd176731: dataIn1 = 32'd8417
; 
32'd176732: dataIn1 = 32'd8418
; 
32'd176733: dataIn1 = 32'd8420
; 
32'd176734: dataIn1 = 32'd5231
; 
32'd176735: dataIn1 = 32'd6468
; 
32'd176736: dataIn1 = 32'd8398
; 
32'd176737: dataIn1 = 32'd8416
; 
32'd176738: dataIn1 = 32'd8419
; 
32'd176739: dataIn1 = 32'd8573
; 
32'd176740: dataIn1 = 32'd8589
; 
32'd176741: dataIn1 = 32'd2726
; 
32'd176742: dataIn1 = 32'd6468
; 
32'd176743: dataIn1 = 32'd8387
; 
32'd176744: dataIn1 = 32'd8418
; 
32'd176745: dataIn1 = 32'd8420
; 
32'd176746: dataIn1 = 32'd8552
; 
32'd176747: dataIn1 = 32'd8591
; 
32'd176748: dataIn1 = 32'd6456
; 
32'd176749: dataIn1 = 32'd6470
; 
32'd176750: dataIn1 = 32'd8378
; 
32'd176751: dataIn1 = 32'd8421
; 
32'd176752: dataIn1 = 32'd8422
; 
32'd176753: dataIn1 = 32'd8423
; 
32'd176754: dataIn1 = 32'd8424
; 
32'd176755: dataIn1 = 32'd6469
; 
32'd176756: dataIn1 = 32'd6470
; 
32'd176757: dataIn1 = 32'd8421
; 
32'd176758: dataIn1 = 32'd8422
; 
32'd176759: dataIn1 = 32'd8423
; 
32'd176760: dataIn1 = 32'd8425
; 
32'd176761: dataIn1 = 32'd8426
; 
32'd176762: dataIn1 = 32'd6456
; 
32'd176763: dataIn1 = 32'd6469
; 
32'd176764: dataIn1 = 32'd8380
; 
32'd176765: dataIn1 = 32'd8421
; 
32'd176766: dataIn1 = 32'd8422
; 
32'd176767: dataIn1 = 32'd8423
; 
32'd176768: dataIn1 = 32'd8427
; 
32'd176769: dataIn1 = 32'd2724
; 
32'd176770: dataIn1 = 32'd6470
; 
32'd176771: dataIn1 = 32'd8378
; 
32'd176772: dataIn1 = 32'd8421
; 
32'd176773: dataIn1 = 32'd8424
; 
32'd176774: dataIn1 = 32'd8441
; 
32'd176775: dataIn1 = 32'd8515
; 
32'd176776: dataIn1 = 32'd5234
; 
32'd176777: dataIn1 = 32'd6470
; 
32'd176778: dataIn1 = 32'd8422
; 
32'd176779: dataIn1 = 32'd8425
; 
32'd176780: dataIn1 = 32'd8426
; 
32'd176781: dataIn1 = 32'd8512
; 
32'd176782: dataIn1 = 32'd8516
; 
32'd176783: dataIn1 = 32'd5234
; 
32'd176784: dataIn1 = 32'd6469
; 
32'd176785: dataIn1 = 32'd6771
; 
32'd176786: dataIn1 = 32'd8422
; 
32'd176787: dataIn1 = 32'd8425
; 
32'd176788: dataIn1 = 32'd8426
; 
32'd176789: dataIn1 = 32'd5228
; 
32'd176790: dataIn1 = 32'd6469
; 
32'd176791: dataIn1 = 32'd6770
; 
32'd176792: dataIn1 = 32'd8380
; 
32'd176793: dataIn1 = 32'd8423
; 
32'd176794: dataIn1 = 32'd8427
; 
32'd176795: dataIn1 = 32'd6472
; 
32'd176796: dataIn1 = 32'd6473
; 
32'd176797: dataIn1 = 32'd8428
; 
32'd176798: dataIn1 = 32'd8429
; 
32'd176799: dataIn1 = 32'd8430
; 
32'd176800: dataIn1 = 32'd8431
; 
32'd176801: dataIn1 = 32'd8432
; 
32'd176802: dataIn1 = 32'd6471
; 
32'd176803: dataIn1 = 32'd6473
; 
32'd176804: dataIn1 = 32'd8428
; 
32'd176805: dataIn1 = 32'd8429
; 
32'd176806: dataIn1 = 32'd8430
; 
32'd176807: dataIn1 = 32'd8433
; 
32'd176808: dataIn1 = 32'd8434
; 
32'd176809: dataIn1 = 32'd6471
; 
32'd176810: dataIn1 = 32'd6472
; 
32'd176811: dataIn1 = 32'd8428
; 
32'd176812: dataIn1 = 32'd8429
; 
32'd176813: dataIn1 = 32'd8430
; 
32'd176814: dataIn1 = 32'd8435
; 
32'd176815: dataIn1 = 32'd8436
; 
32'd176816: dataIn1 = 32'd5235
; 
32'd176817: dataIn1 = 32'd6473
; 
32'd176818: dataIn1 = 32'd8428
; 
32'd176819: dataIn1 = 32'd8431
; 
32'd176820: dataIn1 = 32'd8432
; 
32'd176821: dataIn1 = 32'd8451
; 
32'd176822: dataIn1 = 32'd8454
; 
32'd176823: dataIn1 = 32'd5235
; 
32'd176824: dataIn1 = 32'd6472
; 
32'd176825: dataIn1 = 32'd8428
; 
32'd176826: dataIn1 = 32'd8431
; 
32'd176827: dataIn1 = 32'd8432
; 
32'd176828: dataIn1 = 32'd8444
; 
32'd176829: dataIn1 = 32'd8447
; 
32'd176830: dataIn1 = 32'd5236
; 
32'd176831: dataIn1 = 32'd6473
; 
32'd176832: dataIn1 = 32'd8429
; 
32'd176833: dataIn1 = 32'd8433
; 
32'd176834: dataIn1 = 32'd8434
; 
32'd176835: dataIn1 = 32'd8452
; 
32'd176836: dataIn1 = 32'd8455
; 
32'd176837: dataIn1 = 32'd5236
; 
32'd176838: dataIn1 = 32'd6471
; 
32'd176839: dataIn1 = 32'd8429
; 
32'd176840: dataIn1 = 32'd8433
; 
32'd176841: dataIn1 = 32'd8434
; 
32'd176842: dataIn1 = 32'd8438
; 
32'd176843: dataIn1 = 32'd8442
; 
32'd176844: dataIn1 = 32'd5237
; 
32'd176845: dataIn1 = 32'd6472
; 
32'd176846: dataIn1 = 32'd8430
; 
32'd176847: dataIn1 = 32'd8435
; 
32'd176848: dataIn1 = 32'd8436
; 
32'd176849: dataIn1 = 32'd8446
; 
32'd176850: dataIn1 = 32'd8450
; 
32'd176851: dataIn1 = 32'd5237
; 
32'd176852: dataIn1 = 32'd6471
; 
32'd176853: dataIn1 = 32'd8430
; 
32'd176854: dataIn1 = 32'd8435
; 
32'd176855: dataIn1 = 32'd8436
; 
32'd176856: dataIn1 = 32'd8439
; 
32'd176857: dataIn1 = 32'd8443
; 
32'd176858: dataIn1 = 32'd6474
; 
32'd176859: dataIn1 = 32'd6475
; 
32'd176860: dataIn1 = 32'd8437
; 
32'd176861: dataIn1 = 32'd8438
; 
32'd176862: dataIn1 = 32'd8439
; 
32'd176863: dataIn1 = 32'd8440
; 
32'd176864: dataIn1 = 32'd8441
; 
32'd176865: dataIn1 = 32'd6471
; 
32'd176866: dataIn1 = 32'd6475
; 
32'd176867: dataIn1 = 32'd8434
; 
32'd176868: dataIn1 = 32'd8437
; 
32'd176869: dataIn1 = 32'd8438
; 
32'd176870: dataIn1 = 32'd8439
; 
32'd176871: dataIn1 = 32'd8442
; 
32'd176872: dataIn1 = 32'd6471
; 
32'd176873: dataIn1 = 32'd6474
; 
32'd176874: dataIn1 = 32'd8436
; 
32'd176875: dataIn1 = 32'd8437
; 
32'd176876: dataIn1 = 32'd8438
; 
32'd176877: dataIn1 = 32'd8439
; 
32'd176878: dataIn1 = 32'd8443
; 
32'd176879: dataIn1 = 32'd2724
; 
32'd176880: dataIn1 = 32'd6475
; 
32'd176881: dataIn1 = 32'd8407
; 
32'd176882: dataIn1 = 32'd8437
; 
32'd176883: dataIn1 = 32'd8440
; 
32'd176884: dataIn1 = 32'd8441
; 
32'd176885: dataIn1 = 32'd8493
; 
32'd176886: dataIn1 = 32'd2724
; 
32'd176887: dataIn1 = 32'd6474
; 
32'd176888: dataIn1 = 32'd8424
; 
32'd176889: dataIn1 = 32'd8437
; 
32'd176890: dataIn1 = 32'd8440
; 
32'd176891: dataIn1 = 32'd8441
; 
32'd176892: dataIn1 = 32'd8515
; 
32'd176893: dataIn1 = 32'd5236
; 
32'd176894: dataIn1 = 32'd6475
; 
32'd176895: dataIn1 = 32'd8434
; 
32'd176896: dataIn1 = 32'd8438
; 
32'd176897: dataIn1 = 32'd8442
; 
32'd176898: dataIn1 = 32'd8490
; 
32'd176899: dataIn1 = 32'd8494
; 
32'd176900: dataIn1 = 32'd5237
; 
32'd176901: dataIn1 = 32'd6474
; 
32'd176902: dataIn1 = 32'd8436
; 
32'd176903: dataIn1 = 32'd8439
; 
32'd176904: dataIn1 = 32'd8443
; 
32'd176905: dataIn1 = 32'd8514
; 
32'd176906: dataIn1 = 32'd8517
; 
32'd176907: dataIn1 = 32'd6472
; 
32'd176908: dataIn1 = 32'd6477
; 
32'd176909: dataIn1 = 32'd8432
; 
32'd176910: dataIn1 = 32'd8444
; 
32'd176911: dataIn1 = 32'd8445
; 
32'd176912: dataIn1 = 32'd8446
; 
32'd176913: dataIn1 = 32'd8447
; 
32'd176914: dataIn1 = 32'd6476
; 
32'd176915: dataIn1 = 32'd6477
; 
32'd176916: dataIn1 = 32'd8444
; 
32'd176917: dataIn1 = 32'd8445
; 
32'd176918: dataIn1 = 32'd8446
; 
32'd176919: dataIn1 = 32'd8448
; 
32'd176920: dataIn1 = 32'd8449
; 
32'd176921: dataIn1 = 32'd6472
; 
32'd176922: dataIn1 = 32'd6476
; 
32'd176923: dataIn1 = 32'd8435
; 
32'd176924: dataIn1 = 32'd8444
; 
32'd176925: dataIn1 = 32'd8445
; 
32'd176926: dataIn1 = 32'd8446
; 
32'd176927: dataIn1 = 32'd8450
; 
32'd176928: dataIn1 = 32'd5235
; 
32'd176929: dataIn1 = 32'd6477
; 
32'd176930: dataIn1 = 32'd8432
; 
32'd176931: dataIn1 = 32'd8444
; 
32'd176932: dataIn1 = 32'd8447
; 
32'd176933: dataIn1 = 32'd8462
; 
32'd176934: dataIn1 = 32'd8474
; 
32'd176935: dataIn1 = 32'd2727
; 
32'd176936: dataIn1 = 32'd6477
; 
32'd176937: dataIn1 = 32'd8445
; 
32'd176938: dataIn1 = 32'd8448
; 
32'd176939: dataIn1 = 32'd8449
; 
32'd176940: dataIn1 = 32'd8475
; 
32'd176941: dataIn1 = 32'd8477
; 
32'd176942: dataIn1 = 32'd2727
; 
32'd176943: dataIn1 = 32'd6476
; 
32'd176944: dataIn1 = 32'd8445
; 
32'd176945: dataIn1 = 32'd8448
; 
32'd176946: dataIn1 = 32'd8449
; 
32'd176947: dataIn1 = 32'd8519
; 
32'd176948: dataIn1 = 32'd8522
; 
32'd176949: dataIn1 = 32'd5237
; 
32'd176950: dataIn1 = 32'd6476
; 
32'd176951: dataIn1 = 32'd8435
; 
32'd176952: dataIn1 = 32'd8446
; 
32'd176953: dataIn1 = 32'd8450
; 
32'd176954: dataIn1 = 32'd8513
; 
32'd176955: dataIn1 = 32'd8520
; 
32'd176956: dataIn1 = 32'd6473
; 
32'd176957: dataIn1 = 32'd6479
; 
32'd176958: dataIn1 = 32'd8431
; 
32'd176959: dataIn1 = 32'd8451
; 
32'd176960: dataIn1 = 32'd8452
; 
32'd176961: dataIn1 = 32'd8453
; 
32'd176962: dataIn1 = 32'd8454
; 
32'd176963: dataIn1 = 32'd6473
; 
32'd176964: dataIn1 = 32'd6478
; 
32'd176965: dataIn1 = 32'd8433
; 
32'd176966: dataIn1 = 32'd8451
; 
32'd176967: dataIn1 = 32'd8452
; 
32'd176968: dataIn1 = 32'd8453
; 
32'd176969: dataIn1 = 32'd8455
; 
32'd176970: dataIn1 = 32'd6478
; 
32'd176971: dataIn1 = 32'd6479
; 
32'd176972: dataIn1 = 32'd8451
; 
32'd176973: dataIn1 = 32'd8452
; 
32'd176974: dataIn1 = 32'd8453
; 
32'd176975: dataIn1 = 32'd8456
; 
32'd176976: dataIn1 = 32'd8457
; 
32'd176977: dataIn1 = 32'd5235
; 
32'd176978: dataIn1 = 32'd6479
; 
32'd176979: dataIn1 = 32'd8431
; 
32'd176980: dataIn1 = 32'd8451
; 
32'd176981: dataIn1 = 32'd8454
; 
32'd176982: dataIn1 = 32'd8461
; 
32'd176983: dataIn1 = 32'd8479
; 
32'd176984: dataIn1 = 32'd5236
; 
32'd176985: dataIn1 = 32'd6478
; 
32'd176986: dataIn1 = 32'd8433
; 
32'd176987: dataIn1 = 32'd8452
; 
32'd176988: dataIn1 = 32'd8455
; 
32'd176989: dataIn1 = 32'd8489
; 
32'd176990: dataIn1 = 32'd8502
; 
32'd176991: dataIn1 = 32'd1115
; 
32'd176992: dataIn1 = 32'd6479
; 
32'd176993: dataIn1 = 32'd8453
; 
32'd176994: dataIn1 = 32'd8456
; 
32'd176995: dataIn1 = 32'd8457
; 
32'd176996: dataIn1 = 32'd8481
; 
32'd176997: dataIn1 = 32'd8483
; 
32'd176998: dataIn1 = 32'd1115
; 
32'd176999: dataIn1 = 32'd6478
; 
32'd177000: dataIn1 = 32'd8453
; 
32'd177001: dataIn1 = 32'd8456
; 
32'd177002: dataIn1 = 32'd8457
; 
32'd177003: dataIn1 = 32'd8503
; 
32'd177004: dataIn1 = 32'd8505
; 
32'd177005: dataIn1 = 32'd6481
; 
32'd177006: dataIn1 = 32'd6482
; 
32'd177007: dataIn1 = 32'd8458
; 
32'd177008: dataIn1 = 32'd8459
; 
32'd177009: dataIn1 = 32'd8460
; 
32'd177010: dataIn1 = 32'd8461
; 
32'd177011: dataIn1 = 32'd8462
; 
32'd177012: dataIn1 = 32'd6480
; 
32'd177013: dataIn1 = 32'd6482
; 
32'd177014: dataIn1 = 32'd8458
; 
32'd177015: dataIn1 = 32'd8459
; 
32'd177016: dataIn1 = 32'd8460
; 
32'd177017: dataIn1 = 32'd8463
; 
32'd177018: dataIn1 = 32'd8464
; 
32'd177019: dataIn1 = 32'd6480
; 
32'd177020: dataIn1 = 32'd6481
; 
32'd177021: dataIn1 = 32'd8458
; 
32'd177022: dataIn1 = 32'd8459
; 
32'd177023: dataIn1 = 32'd8460
; 
32'd177024: dataIn1 = 32'd8465
; 
32'd177025: dataIn1 = 32'd8466
; 
32'd177026: dataIn1 = 32'd5235
; 
32'd177027: dataIn1 = 32'd6482
; 
32'd177028: dataIn1 = 32'd8454
; 
32'd177029: dataIn1 = 32'd8458
; 
32'd177030: dataIn1 = 32'd8461
; 
32'd177031: dataIn1 = 32'd8462
; 
32'd177032: dataIn1 = 32'd8479
; 
32'd177033: dataIn1 = 32'd5235
; 
32'd177034: dataIn1 = 32'd6481
; 
32'd177035: dataIn1 = 32'd8447
; 
32'd177036: dataIn1 = 32'd8458
; 
32'd177037: dataIn1 = 32'd8461
; 
32'd177038: dataIn1 = 32'd8462
; 
32'd177039: dataIn1 = 32'd8474
; 
32'd177040: dataIn1 = 32'd2676
; 
32'd177041: dataIn1 = 32'd6482
; 
32'd177042: dataIn1 = 32'd8459
; 
32'd177043: dataIn1 = 32'd8463
; 
32'd177044: dataIn1 = 32'd8464
; 
32'd177045: dataIn1 = 32'd8480
; 
32'd177046: dataIn1 = 32'd8482
; 
32'd177047: dataIn1 = 32'd2676
; 
32'd177048: dataIn1 = 32'd6480
; 
32'd177049: dataIn1 = 32'd8459
; 
32'd177050: dataIn1 = 32'd8463
; 
32'd177051: dataIn1 = 32'd8464
; 
32'd177052: dataIn1 = 32'd8468
; 
32'd177053: dataIn1 = 32'd8472
; 
32'd177054: dataIn1 = 32'd5238
; 
32'd177055: dataIn1 = 32'd6481
; 
32'd177056: dataIn1 = 32'd8460
; 
32'd177057: dataIn1 = 32'd8465
; 
32'd177058: dataIn1 = 32'd8466
; 
32'd177059: dataIn1 = 32'd8476
; 
32'd177060: dataIn1 = 32'd8478
; 
32'd177061: dataIn1 = 32'd5238
; 
32'd177062: dataIn1 = 32'd6480
; 
32'd177063: dataIn1 = 32'd8460
; 
32'd177064: dataIn1 = 32'd8465
; 
32'd177065: dataIn1 = 32'd8466
; 
32'd177066: dataIn1 = 32'd8469
; 
32'd177067: dataIn1 = 32'd8473
; 
32'd177068: dataIn1 = 32'd5053
; 
32'd177069: dataIn1 = 32'd6483
; 
32'd177070: dataIn1 = 32'd8467
; 
32'd177071: dataIn1 = 32'd8468
; 
32'd177072: dataIn1 = 32'd8469
; 
32'd177073: dataIn1 = 32'd8470
; 
32'd177074: dataIn1 = 32'd8471
; 
32'd177075: dataIn1 = 32'd5053
; 
32'd177076: dataIn1 = 32'd6480
; 
32'd177077: dataIn1 = 32'd8464
; 
32'd177078: dataIn1 = 32'd8467
; 
32'd177079: dataIn1 = 32'd8468
; 
32'd177080: dataIn1 = 32'd8469
; 
32'd177081: dataIn1 = 32'd8472
; 
32'd177082: dataIn1 = 32'd6480
; 
32'd177083: dataIn1 = 32'd6483
; 
32'd177084: dataIn1 = 32'd8466
; 
32'd177085: dataIn1 = 32'd8467
; 
32'd177086: dataIn1 = 32'd8468
; 
32'd177087: dataIn1 = 32'd8469
; 
32'd177088: dataIn1 = 32'd8473
; 
32'd177089: dataIn1 = 32'd10
; 
32'd177090: dataIn1 = 32'd4753
; 
32'd177091: dataIn1 = 32'd5053
; 
32'd177092: dataIn1 = 32'd8467
; 
32'd177093: dataIn1 = 32'd8470
; 
32'd177094: dataIn1 = 32'd8471
; 
32'd177095: dataIn1 = 32'd10
; 
32'd177096: dataIn1 = 32'd6483
; 
32'd177097: dataIn1 = 32'd8363
; 
32'd177098: dataIn1 = 32'd8467
; 
32'd177099: dataIn1 = 32'd8470
; 
32'd177100: dataIn1 = 32'd8471
; 
32'd177101: dataIn1 = 32'd9163
; 
32'd177102: dataIn1 = 32'd2676
; 
32'd177103: dataIn1 = 32'd5051
; 
32'd177104: dataIn1 = 32'd5053
; 
32'd177105: dataIn1 = 32'd8464
; 
32'd177106: dataIn1 = 32'd8468
; 
32'd177107: dataIn1 = 32'd8472
; 
32'd177108: dataIn1 = 32'd5238
; 
32'd177109: dataIn1 = 32'd6483
; 
32'd177110: dataIn1 = 32'd8466
; 
32'd177111: dataIn1 = 32'd8469
; 
32'd177112: dataIn1 = 32'd8473
; 
32'd177113: dataIn1 = 32'd9160
; 
32'd177114: dataIn1 = 32'd9164
; 
32'd177115: dataIn1 = 32'd6477
; 
32'd177116: dataIn1 = 32'd6481
; 
32'd177117: dataIn1 = 32'd8447
; 
32'd177118: dataIn1 = 32'd8462
; 
32'd177119: dataIn1 = 32'd8474
; 
32'd177120: dataIn1 = 32'd8475
; 
32'd177121: dataIn1 = 32'd8476
; 
32'd177122: dataIn1 = 32'd6477
; 
32'd177123: dataIn1 = 32'd6484
; 
32'd177124: dataIn1 = 32'd8448
; 
32'd177125: dataIn1 = 32'd8474
; 
32'd177126: dataIn1 = 32'd8475
; 
32'd177127: dataIn1 = 32'd8476
; 
32'd177128: dataIn1 = 32'd8477
; 
32'd177129: dataIn1 = 32'd6481
; 
32'd177130: dataIn1 = 32'd6484
; 
32'd177131: dataIn1 = 32'd8465
; 
32'd177132: dataIn1 = 32'd8474
; 
32'd177133: dataIn1 = 32'd8475
; 
32'd177134: dataIn1 = 32'd8476
; 
32'd177135: dataIn1 = 32'd8478
; 
32'd177136: dataIn1 = 32'd2727
; 
32'd177137: dataIn1 = 32'd6484
; 
32'd177138: dataIn1 = 32'd8448
; 
32'd177139: dataIn1 = 32'd8475
; 
32'd177140: dataIn1 = 32'd8477
; 
32'd177141: dataIn1 = 32'd9152
; 
32'd177142: dataIn1 = 32'd9171
; 
32'd177143: dataIn1 = 32'd5238
; 
32'd177144: dataIn1 = 32'd6484
; 
32'd177145: dataIn1 = 32'd8465
; 
32'd177146: dataIn1 = 32'd8476
; 
32'd177147: dataIn1 = 32'd8478
; 
32'd177148: dataIn1 = 32'd9159
; 
32'd177149: dataIn1 = 32'd9170
; 
32'd177150: dataIn1 = 32'd6479
; 
32'd177151: dataIn1 = 32'd6482
; 
32'd177152: dataIn1 = 32'd8454
; 
32'd177153: dataIn1 = 32'd8461
; 
32'd177154: dataIn1 = 32'd8479
; 
32'd177155: dataIn1 = 32'd8480
; 
32'd177156: dataIn1 = 32'd8481
; 
32'd177157: dataIn1 = 32'd5054
; 
32'd177158: dataIn1 = 32'd6482
; 
32'd177159: dataIn1 = 32'd8463
; 
32'd177160: dataIn1 = 32'd8479
; 
32'd177161: dataIn1 = 32'd8480
; 
32'd177162: dataIn1 = 32'd8481
; 
32'd177163: dataIn1 = 32'd8482
; 
32'd177164: dataIn1 = 32'd5054
; 
32'd177165: dataIn1 = 32'd6479
; 
32'd177166: dataIn1 = 32'd8456
; 
32'd177167: dataIn1 = 32'd8479
; 
32'd177168: dataIn1 = 32'd8480
; 
32'd177169: dataIn1 = 32'd8481
; 
32'd177170: dataIn1 = 32'd8483
; 
32'd177171: dataIn1 = 32'd2676
; 
32'd177172: dataIn1 = 32'd5052
; 
32'd177173: dataIn1 = 32'd5054
; 
32'd177174: dataIn1 = 32'd8463
; 
32'd177175: dataIn1 = 32'd8480
; 
32'd177176: dataIn1 = 32'd8482
; 
32'd177177: dataIn1 = 32'd1115
; 
32'd177178: dataIn1 = 32'd5043
; 
32'd177179: dataIn1 = 32'd5054
; 
32'd177180: dataIn1 = 32'd8456
; 
32'd177181: dataIn1 = 32'd8481
; 
32'd177182: dataIn1 = 32'd8483
; 
32'd177183: dataIn1 = 32'd6486
; 
32'd177184: dataIn1 = 32'd6487
; 
32'd177185: dataIn1 = 32'd8484
; 
32'd177186: dataIn1 = 32'd8485
; 
32'd177187: dataIn1 = 32'd8486
; 
32'd177188: dataIn1 = 32'd8487
; 
32'd177189: dataIn1 = 32'd8488
; 
32'd177190: dataIn1 = 32'd6485
; 
32'd177191: dataIn1 = 32'd6487
; 
32'd177192: dataIn1 = 32'd8484
; 
32'd177193: dataIn1 = 32'd8485
; 
32'd177194: dataIn1 = 32'd8486
; 
32'd177195: dataIn1 = 32'd8489
; 
32'd177196: dataIn1 = 32'd8490
; 
32'd177197: dataIn1 = 32'd6485
; 
32'd177198: dataIn1 = 32'd6486
; 
32'd177199: dataIn1 = 32'd8484
; 
32'd177200: dataIn1 = 32'd8485
; 
32'd177201: dataIn1 = 32'd8486
; 
32'd177202: dataIn1 = 32'd8491
; 
32'd177203: dataIn1 = 32'd8492
; 
32'd177204: dataIn1 = 32'd2675
; 
32'd177205: dataIn1 = 32'd6487
; 
32'd177206: dataIn1 = 32'd8484
; 
32'd177207: dataIn1 = 32'd8487
; 
32'd177208: dataIn1 = 32'd8488
; 
32'd177209: dataIn1 = 32'd8501
; 
32'd177210: dataIn1 = 32'd8504
; 
32'd177211: dataIn1 = 32'd2675
; 
32'd177212: dataIn1 = 32'd6486
; 
32'd177213: dataIn1 = 32'd8484
; 
32'd177214: dataIn1 = 32'd8487
; 
32'd177215: dataIn1 = 32'd8488
; 
32'd177216: dataIn1 = 32'd8496
; 
32'd177217: dataIn1 = 32'd8499
; 
32'd177218: dataIn1 = 32'd5236
; 
32'd177219: dataIn1 = 32'd6487
; 
32'd177220: dataIn1 = 32'd8455
; 
32'd177221: dataIn1 = 32'd8485
; 
32'd177222: dataIn1 = 32'd8489
; 
32'd177223: dataIn1 = 32'd8490
; 
32'd177224: dataIn1 = 32'd8502
; 
32'd177225: dataIn1 = 32'd5236
; 
32'd177226: dataIn1 = 32'd6485
; 
32'd177227: dataIn1 = 32'd8442
; 
32'd177228: dataIn1 = 32'd8485
; 
32'd177229: dataIn1 = 32'd8489
; 
32'd177230: dataIn1 = 32'd8490
; 
32'd177231: dataIn1 = 32'd8494
; 
32'd177232: dataIn1 = 32'd5232
; 
32'd177233: dataIn1 = 32'd6486
; 
32'd177234: dataIn1 = 32'd8415
; 
32'd177235: dataIn1 = 32'd8486
; 
32'd177236: dataIn1 = 32'd8491
; 
32'd177237: dataIn1 = 32'd8492
; 
32'd177238: dataIn1 = 32'd8498
; 
32'd177239: dataIn1 = 32'd5232
; 
32'd177240: dataIn1 = 32'd6485
; 
32'd177241: dataIn1 = 32'd8408
; 
32'd177242: dataIn1 = 32'd8486
; 
32'd177243: dataIn1 = 32'd8491
; 
32'd177244: dataIn1 = 32'd8492
; 
32'd177245: dataIn1 = 32'd8495
; 
32'd177246: dataIn1 = 32'd6465
; 
32'd177247: dataIn1 = 32'd6475
; 
32'd177248: dataIn1 = 32'd8407
; 
32'd177249: dataIn1 = 32'd8440
; 
32'd177250: dataIn1 = 32'd8493
; 
32'd177251: dataIn1 = 32'd8494
; 
32'd177252: dataIn1 = 32'd8495
; 
32'd177253: dataIn1 = 32'd6475
; 
32'd177254: dataIn1 = 32'd6485
; 
32'd177255: dataIn1 = 32'd8442
; 
32'd177256: dataIn1 = 32'd8490
; 
32'd177257: dataIn1 = 32'd8493
; 
32'd177258: dataIn1 = 32'd8494
; 
32'd177259: dataIn1 = 32'd8495
; 
32'd177260: dataIn1 = 32'd6465
; 
32'd177261: dataIn1 = 32'd6485
; 
32'd177262: dataIn1 = 32'd8408
; 
32'd177263: dataIn1 = 32'd8492
; 
32'd177264: dataIn1 = 32'd8493
; 
32'd177265: dataIn1 = 32'd8494
; 
32'd177266: dataIn1 = 32'd8495
; 
32'd177267: dataIn1 = 32'd5048
; 
32'd177268: dataIn1 = 32'd6486
; 
32'd177269: dataIn1 = 32'd8488
; 
32'd177270: dataIn1 = 32'd8496
; 
32'd177271: dataIn1 = 32'd8497
; 
32'd177272: dataIn1 = 32'd8498
; 
32'd177273: dataIn1 = 32'd8499
; 
32'd177274: dataIn1 = 32'd5048
; 
32'd177275: dataIn1 = 32'd6466
; 
32'd177276: dataIn1 = 32'd8414
; 
32'd177277: dataIn1 = 32'd8496
; 
32'd177278: dataIn1 = 32'd8497
; 
32'd177279: dataIn1 = 32'd8498
; 
32'd177280: dataIn1 = 32'd8500
; 
32'd177281: dataIn1 = 32'd6466
; 
32'd177282: dataIn1 = 32'd6486
; 
32'd177283: dataIn1 = 32'd8415
; 
32'd177284: dataIn1 = 32'd8491
; 
32'd177285: dataIn1 = 32'd8496
; 
32'd177286: dataIn1 = 32'd8497
; 
32'd177287: dataIn1 = 32'd8498
; 
32'd177288: dataIn1 = 32'd2675
; 
32'd177289: dataIn1 = 32'd5045
; 
32'd177290: dataIn1 = 32'd5048
; 
32'd177291: dataIn1 = 32'd8488
; 
32'd177292: dataIn1 = 32'd8496
; 
32'd177293: dataIn1 = 32'd8499
; 
32'd177294: dataIn1 = 32'd145
; 
32'd177295: dataIn1 = 32'd4759
; 
32'd177296: dataIn1 = 32'd5048
; 
32'd177297: dataIn1 = 32'd8414
; 
32'd177298: dataIn1 = 32'd8497
; 
32'd177299: dataIn1 = 32'd8500
; 
32'd177300: dataIn1 = 32'd5049
; 
32'd177301: dataIn1 = 32'd6487
; 
32'd177302: dataIn1 = 32'd8487
; 
32'd177303: dataIn1 = 32'd8501
; 
32'd177304: dataIn1 = 32'd8502
; 
32'd177305: dataIn1 = 32'd8503
; 
32'd177306: dataIn1 = 32'd8504
; 
32'd177307: dataIn1 = 32'd6478
; 
32'd177308: dataIn1 = 32'd6487
; 
32'd177309: dataIn1 = 32'd8455
; 
32'd177310: dataIn1 = 32'd8489
; 
32'd177311: dataIn1 = 32'd8501
; 
32'd177312: dataIn1 = 32'd8502
; 
32'd177313: dataIn1 = 32'd8503
; 
32'd177314: dataIn1 = 32'd5049
; 
32'd177315: dataIn1 = 32'd6478
; 
32'd177316: dataIn1 = 32'd8457
; 
32'd177317: dataIn1 = 32'd8501
; 
32'd177318: dataIn1 = 32'd8502
; 
32'd177319: dataIn1 = 32'd8503
; 
32'd177320: dataIn1 = 32'd8505
; 
32'd177321: dataIn1 = 32'd2675
; 
32'd177322: dataIn1 = 32'd5047
; 
32'd177323: dataIn1 = 32'd5049
; 
32'd177324: dataIn1 = 32'd8487
; 
32'd177325: dataIn1 = 32'd8501
; 
32'd177326: dataIn1 = 32'd8504
; 
32'd177327: dataIn1 = 32'd1115
; 
32'd177328: dataIn1 = 32'd5044
; 
32'd177329: dataIn1 = 32'd5049
; 
32'd177330: dataIn1 = 32'd8457
; 
32'd177331: dataIn1 = 32'd8503
; 
32'd177332: dataIn1 = 32'd8505
; 
32'd177333: dataIn1 = 32'd6489
; 
32'd177334: dataIn1 = 32'd6490
; 
32'd177335: dataIn1 = 32'd8506
; 
32'd177336: dataIn1 = 32'd8507
; 
32'd177337: dataIn1 = 32'd8508
; 
32'd177338: dataIn1 = 32'd8509
; 
32'd177339: dataIn1 = 32'd8510
; 
32'd177340: dataIn1 = 32'd6488
; 
32'd177341: dataIn1 = 32'd6490
; 
32'd177342: dataIn1 = 32'd8506
; 
32'd177343: dataIn1 = 32'd8507
; 
32'd177344: dataIn1 = 32'd8508
; 
32'd177345: dataIn1 = 32'd8511
; 
32'd177346: dataIn1 = 32'd8512
; 
32'd177347: dataIn1 = 32'd6488
; 
32'd177348: dataIn1 = 32'd6489
; 
32'd177349: dataIn1 = 32'd8506
; 
32'd177350: dataIn1 = 32'd8507
; 
32'd177351: dataIn1 = 32'd8508
; 
32'd177352: dataIn1 = 32'd8513
; 
32'd177353: dataIn1 = 32'd8514
; 
32'd177354: dataIn1 = 32'd5239
; 
32'd177355: dataIn1 = 32'd6490
; 
32'd177356: dataIn1 = 32'd6773
; 
32'd177357: dataIn1 = 32'd8506
; 
32'd177358: dataIn1 = 32'd8509
; 
32'd177359: dataIn1 = 32'd8510
; 
32'd177360: dataIn1 = 32'd5239
; 
32'd177361: dataIn1 = 32'd6489
; 
32'd177362: dataIn1 = 32'd8506
; 
32'd177363: dataIn1 = 32'd8509
; 
32'd177364: dataIn1 = 32'd8510
; 
32'd177365: dataIn1 = 32'd8518
; 
32'd177366: dataIn1 = 32'd8521
; 
32'd177367: dataIn1 = 32'd5234
; 
32'd177368: dataIn1 = 32'd6490
; 
32'd177369: dataIn1 = 32'd6772
; 
32'd177370: dataIn1 = 32'd8507
; 
32'd177371: dataIn1 = 32'd8511
; 
32'd177372: dataIn1 = 32'd8512
; 
32'd177373: dataIn1 = 32'd5234
; 
32'd177374: dataIn1 = 32'd6488
; 
32'd177375: dataIn1 = 32'd8425
; 
32'd177376: dataIn1 = 32'd8507
; 
32'd177377: dataIn1 = 32'd8511
; 
32'd177378: dataIn1 = 32'd8512
; 
32'd177379: dataIn1 = 32'd8516
; 
32'd177380: dataIn1 = 32'd5237
; 
32'd177381: dataIn1 = 32'd6489
; 
32'd177382: dataIn1 = 32'd8450
; 
32'd177383: dataIn1 = 32'd8508
; 
32'd177384: dataIn1 = 32'd8513
; 
32'd177385: dataIn1 = 32'd8514
; 
32'd177386: dataIn1 = 32'd8520
; 
32'd177387: dataIn1 = 32'd5237
; 
32'd177388: dataIn1 = 32'd6488
; 
32'd177389: dataIn1 = 32'd8443
; 
32'd177390: dataIn1 = 32'd8508
; 
32'd177391: dataIn1 = 32'd8513
; 
32'd177392: dataIn1 = 32'd8514
; 
32'd177393: dataIn1 = 32'd8517
; 
32'd177394: dataIn1 = 32'd6470
; 
32'd177395: dataIn1 = 32'd6474
; 
32'd177396: dataIn1 = 32'd8424
; 
32'd177397: dataIn1 = 32'd8441
; 
32'd177398: dataIn1 = 32'd8515
; 
32'd177399: dataIn1 = 32'd8516
; 
32'd177400: dataIn1 = 32'd8517
; 
32'd177401: dataIn1 = 32'd6470
; 
32'd177402: dataIn1 = 32'd6488
; 
32'd177403: dataIn1 = 32'd8425
; 
32'd177404: dataIn1 = 32'd8512
; 
32'd177405: dataIn1 = 32'd8515
; 
32'd177406: dataIn1 = 32'd8516
; 
32'd177407: dataIn1 = 32'd8517
; 
32'd177408: dataIn1 = 32'd6474
; 
32'd177409: dataIn1 = 32'd6488
; 
32'd177410: dataIn1 = 32'd8443
; 
32'd177411: dataIn1 = 32'd8514
; 
32'd177412: dataIn1 = 32'd8515
; 
32'd177413: dataIn1 = 32'd8516
; 
32'd177414: dataIn1 = 32'd8517
; 
32'd177415: dataIn1 = 32'd6489
; 
32'd177416: dataIn1 = 32'd6491
; 
32'd177417: dataIn1 = 32'd8510
; 
32'd177418: dataIn1 = 32'd8518
; 
32'd177419: dataIn1 = 32'd8519
; 
32'd177420: dataIn1 = 32'd8520
; 
32'd177421: dataIn1 = 32'd8521
; 
32'd177422: dataIn1 = 32'd6476
; 
32'd177423: dataIn1 = 32'd6491
; 
32'd177424: dataIn1 = 32'd8449
; 
32'd177425: dataIn1 = 32'd8518
; 
32'd177426: dataIn1 = 32'd8519
; 
32'd177427: dataIn1 = 32'd8520
; 
32'd177428: dataIn1 = 32'd8522
; 
32'd177429: dataIn1 = 32'd6476
; 
32'd177430: dataIn1 = 32'd6489
; 
32'd177431: dataIn1 = 32'd8450
; 
32'd177432: dataIn1 = 32'd8513
; 
32'd177433: dataIn1 = 32'd8518
; 
32'd177434: dataIn1 = 32'd8519
; 
32'd177435: dataIn1 = 32'd8520
; 
32'd177436: dataIn1 = 32'd5239
; 
32'd177437: dataIn1 = 32'd6491
; 
32'd177438: dataIn1 = 32'd8510
; 
32'd177439: dataIn1 = 32'd8518
; 
32'd177440: dataIn1 = 32'd8521
; 
32'd177441: dataIn1 = 32'd9172
; 
32'd177442: dataIn1 = 32'd9175
; 
32'd177443: dataIn1 = 32'd2727
; 
32'd177444: dataIn1 = 32'd6491
; 
32'd177445: dataIn1 = 32'd8449
; 
32'd177446: dataIn1 = 32'd8519
; 
32'd177447: dataIn1 = 32'd8522
; 
32'd177448: dataIn1 = 32'd9153
; 
32'd177449: dataIn1 = 32'd9174
; 
32'd177450: dataIn1 = 32'd6493
; 
32'd177451: dataIn1 = 32'd6494
; 
32'd177452: dataIn1 = 32'd8523
; 
32'd177453: dataIn1 = 32'd8524
; 
32'd177454: dataIn1 = 32'd8525
; 
32'd177455: dataIn1 = 32'd8526
; 
32'd177456: dataIn1 = 32'd8527
; 
32'd177457: dataIn1 = 32'd6492
; 
32'd177458: dataIn1 = 32'd6494
; 
32'd177459: dataIn1 = 32'd8523
; 
32'd177460: dataIn1 = 32'd8524
; 
32'd177461: dataIn1 = 32'd8525
; 
32'd177462: dataIn1 = 32'd8528
; 
32'd177463: dataIn1 = 32'd8529
; 
32'd177464: dataIn1 = 32'd6492
; 
32'd177465: dataIn1 = 32'd6493
; 
32'd177466: dataIn1 = 32'd8523
; 
32'd177467: dataIn1 = 32'd8524
; 
32'd177468: dataIn1 = 32'd8525
; 
32'd177469: dataIn1 = 32'd8530
; 
32'd177470: dataIn1 = 32'd8531
; 
32'd177471: dataIn1 = 32'd5240
; 
32'd177472: dataIn1 = 32'd6494
; 
32'd177473: dataIn1 = 32'd8523
; 
32'd177474: dataIn1 = 32'd8526
; 
32'd177475: dataIn1 = 32'd8527
; 
32'd177476: dataIn1 = 32'd8546
; 
32'd177477: dataIn1 = 32'd8549
; 
32'd177478: dataIn1 = 32'd5240
; 
32'd177479: dataIn1 = 32'd6493
; 
32'd177480: dataIn1 = 32'd8523
; 
32'd177481: dataIn1 = 32'd8526
; 
32'd177482: dataIn1 = 32'd8527
; 
32'd177483: dataIn1 = 32'd8539
; 
32'd177484: dataIn1 = 32'd8542
; 
32'd177485: dataIn1 = 32'd5241
; 
32'd177486: dataIn1 = 32'd6494
; 
32'd177487: dataIn1 = 32'd8524
; 
32'd177488: dataIn1 = 32'd8528
; 
32'd177489: dataIn1 = 32'd8529
; 
32'd177490: dataIn1 = 32'd8547
; 
32'd177491: dataIn1 = 32'd8550
; 
32'd177492: dataIn1 = 32'd5241
; 
32'd177493: dataIn1 = 32'd6492
; 
32'd177494: dataIn1 = 32'd8524
; 
32'd177495: dataIn1 = 32'd8528
; 
32'd177496: dataIn1 = 32'd8529
; 
32'd177497: dataIn1 = 32'd8533
; 
32'd177498: dataIn1 = 32'd8537
; 
32'd177499: dataIn1 = 32'd5242
; 
32'd177500: dataIn1 = 32'd6493
; 
32'd177501: dataIn1 = 32'd8525
; 
32'd177502: dataIn1 = 32'd8530
; 
32'd177503: dataIn1 = 32'd8531
; 
32'd177504: dataIn1 = 32'd8541
; 
32'd177505: dataIn1 = 32'd8545
; 
32'd177506: dataIn1 = 32'd5242
; 
32'd177507: dataIn1 = 32'd6492
; 
32'd177508: dataIn1 = 32'd8525
; 
32'd177509: dataIn1 = 32'd8530
; 
32'd177510: dataIn1 = 32'd8531
; 
32'd177511: dataIn1 = 32'd8534
; 
32'd177512: dataIn1 = 32'd8538
; 
32'd177513: dataIn1 = 32'd6495
; 
32'd177514: dataIn1 = 32'd6496
; 
32'd177515: dataIn1 = 32'd8532
; 
32'd177516: dataIn1 = 32'd8533
; 
32'd177517: dataIn1 = 32'd8534
; 
32'd177518: dataIn1 = 32'd8535
; 
32'd177519: dataIn1 = 32'd8536
; 
32'd177520: dataIn1 = 32'd6492
; 
32'd177521: dataIn1 = 32'd6496
; 
32'd177522: dataIn1 = 32'd8529
; 
32'd177523: dataIn1 = 32'd8532
; 
32'd177524: dataIn1 = 32'd8533
; 
32'd177525: dataIn1 = 32'd8534
; 
32'd177526: dataIn1 = 32'd8537
; 
32'd177527: dataIn1 = 32'd6492
; 
32'd177528: dataIn1 = 32'd6495
; 
32'd177529: dataIn1 = 32'd8531
; 
32'd177530: dataIn1 = 32'd8532
; 
32'd177531: dataIn1 = 32'd8533
; 
32'd177532: dataIn1 = 32'd8534
; 
32'd177533: dataIn1 = 32'd8538
; 
32'd177534: dataIn1 = 32'd1116
; 
32'd177535: dataIn1 = 32'd6496
; 
32'd177536: dataIn1 = 32'd8532
; 
32'd177537: dataIn1 = 32'd8535
; 
32'd177538: dataIn1 = 32'd8536
; 
32'd177539: dataIn1 = 32'd8579
; 
32'd177540: dataIn1 = 32'd8582
; 
32'd177541: dataIn1 = 32'd1116
; 
32'd177542: dataIn1 = 32'd6495
; 
32'd177543: dataIn1 = 32'd8532
; 
32'd177544: dataIn1 = 32'd8535
; 
32'd177545: dataIn1 = 32'd8536
; 
32'd177546: dataIn1 = 32'd8601
; 
32'd177547: dataIn1 = 32'd8604
; 
32'd177548: dataIn1 = 32'd5241
; 
32'd177549: dataIn1 = 32'd6496
; 
32'd177550: dataIn1 = 32'd8529
; 
32'd177551: dataIn1 = 32'd8533
; 
32'd177552: dataIn1 = 32'd8537
; 
32'd177553: dataIn1 = 32'd8576
; 
32'd177554: dataIn1 = 32'd8580
; 
32'd177555: dataIn1 = 32'd5242
; 
32'd177556: dataIn1 = 32'd6495
; 
32'd177557: dataIn1 = 32'd8531
; 
32'd177558: dataIn1 = 32'd8534
; 
32'd177559: dataIn1 = 32'd8538
; 
32'd177560: dataIn1 = 32'd8600
; 
32'd177561: dataIn1 = 32'd8603
; 
32'd177562: dataIn1 = 32'd6493
; 
32'd177563: dataIn1 = 32'd6498
; 
32'd177564: dataIn1 = 32'd8527
; 
32'd177565: dataIn1 = 32'd8539
; 
32'd177566: dataIn1 = 32'd8540
; 
32'd177567: dataIn1 = 32'd8541
; 
32'd177568: dataIn1 = 32'd8542
; 
32'd177569: dataIn1 = 32'd6497
; 
32'd177570: dataIn1 = 32'd6498
; 
32'd177571: dataIn1 = 32'd8539
; 
32'd177572: dataIn1 = 32'd8540
; 
32'd177573: dataIn1 = 32'd8541
; 
32'd177574: dataIn1 = 32'd8543
; 
32'd177575: dataIn1 = 32'd8544
; 
32'd177576: dataIn1 = 32'd6493
; 
32'd177577: dataIn1 = 32'd6497
; 
32'd177578: dataIn1 = 32'd8530
; 
32'd177579: dataIn1 = 32'd8539
; 
32'd177580: dataIn1 = 32'd8540
; 
32'd177581: dataIn1 = 32'd8541
; 
32'd177582: dataIn1 = 32'd8545
; 
32'd177583: dataIn1 = 32'd5240
; 
32'd177584: dataIn1 = 32'd6498
; 
32'd177585: dataIn1 = 32'd8527
; 
32'd177586: dataIn1 = 32'd8539
; 
32'd177587: dataIn1 = 32'd8542
; 
32'd177588: dataIn1 = 32'd8557
; 
32'd177589: dataIn1 = 32'd8562
; 
32'd177590: dataIn1 = 32'd2728
; 
32'd177591: dataIn1 = 32'd6498
; 
32'd177592: dataIn1 = 32'd8540
; 
32'd177593: dataIn1 = 32'd8543
; 
32'd177594: dataIn1 = 32'd8544
; 
32'd177595: dataIn1 = 32'd8563
; 
32'd177596: dataIn1 = 32'd8565
; 
32'd177597: dataIn1 = 32'd2728
; 
32'd177598: dataIn1 = 32'd6497
; 
32'd177599: dataIn1 = 32'd8540
; 
32'd177600: dataIn1 = 32'd8543
; 
32'd177601: dataIn1 = 32'd8544
; 
32'd177602: dataIn1 = 32'd8607
; 
32'd177603: dataIn1 = 32'd8610
; 
32'd177604: dataIn1 = 32'd5242
; 
32'd177605: dataIn1 = 32'd6497
; 
32'd177606: dataIn1 = 32'd8530
; 
32'd177607: dataIn1 = 32'd8541
; 
32'd177608: dataIn1 = 32'd8545
; 
32'd177609: dataIn1 = 32'd8599
; 
32'd177610: dataIn1 = 32'd8608
; 
32'd177611: dataIn1 = 32'd6494
; 
32'd177612: dataIn1 = 32'd6500
; 
32'd177613: dataIn1 = 32'd8526
; 
32'd177614: dataIn1 = 32'd8546
; 
32'd177615: dataIn1 = 32'd8547
; 
32'd177616: dataIn1 = 32'd8548
; 
32'd177617: dataIn1 = 32'd8549
; 
32'd177618: dataIn1 = 32'd6494
; 
32'd177619: dataIn1 = 32'd6499
; 
32'd177620: dataIn1 = 32'd8528
; 
32'd177621: dataIn1 = 32'd8546
; 
32'd177622: dataIn1 = 32'd8547
; 
32'd177623: dataIn1 = 32'd8548
; 
32'd177624: dataIn1 = 32'd8550
; 
32'd177625: dataIn1 = 32'd6499
; 
32'd177626: dataIn1 = 32'd6500
; 
32'd177627: dataIn1 = 32'd8546
; 
32'd177628: dataIn1 = 32'd8547
; 
32'd177629: dataIn1 = 32'd8548
; 
32'd177630: dataIn1 = 32'd8551
; 
32'd177631: dataIn1 = 32'd8552
; 
32'd177632: dataIn1 = 32'd5240
; 
32'd177633: dataIn1 = 32'd6500
; 
32'd177634: dataIn1 = 32'd8526
; 
32'd177635: dataIn1 = 32'd8546
; 
32'd177636: dataIn1 = 32'd8549
; 
32'd177637: dataIn1 = 32'd8556
; 
32'd177638: dataIn1 = 32'd8567
; 
32'd177639: dataIn1 = 32'd5241
; 
32'd177640: dataIn1 = 32'd6499
; 
32'd177641: dataIn1 = 32'd8528
; 
32'd177642: dataIn1 = 32'd8547
; 
32'd177643: dataIn1 = 32'd8550
; 
32'd177644: dataIn1 = 32'd8575
; 
32'd177645: dataIn1 = 32'd8590
; 
32'd177646: dataIn1 = 32'd2726
; 
32'd177647: dataIn1 = 32'd6500
; 
32'd177648: dataIn1 = 32'd8394
; 
32'd177649: dataIn1 = 32'd8548
; 
32'd177650: dataIn1 = 32'd8551
; 
32'd177651: dataIn1 = 32'd8552
; 
32'd177652: dataIn1 = 32'd8569
; 
32'd177653: dataIn1 = 32'd2726
; 
32'd177654: dataIn1 = 32'd6499
; 
32'd177655: dataIn1 = 32'd8420
; 
32'd177656: dataIn1 = 32'd8548
; 
32'd177657: dataIn1 = 32'd8551
; 
32'd177658: dataIn1 = 32'd8552
; 
32'd177659: dataIn1 = 32'd8591
; 
32'd177660: dataIn1 = 32'd6502
; 
32'd177661: dataIn1 = 32'd6503
; 
32'd177662: dataIn1 = 32'd8553
; 
32'd177663: dataIn1 = 32'd8554
; 
32'd177664: dataIn1 = 32'd8555
; 
32'd177665: dataIn1 = 32'd8556
; 
32'd177666: dataIn1 = 32'd8557
; 
32'd177667: dataIn1 = 32'd6501
; 
32'd177668: dataIn1 = 32'd6503
; 
32'd177669: dataIn1 = 32'd8553
; 
32'd177670: dataIn1 = 32'd8554
; 
32'd177671: dataIn1 = 32'd8555
; 
32'd177672: dataIn1 = 32'd8558
; 
32'd177673: dataIn1 = 32'd8559
; 
32'd177674: dataIn1 = 32'd6501
; 
32'd177675: dataIn1 = 32'd6502
; 
32'd177676: dataIn1 = 32'd8553
; 
32'd177677: dataIn1 = 32'd8554
; 
32'd177678: dataIn1 = 32'd8555
; 
32'd177679: dataIn1 = 32'd8560
; 
32'd177680: dataIn1 = 32'd8561
; 
32'd177681: dataIn1 = 32'd5240
; 
32'd177682: dataIn1 = 32'd6503
; 
32'd177683: dataIn1 = 32'd8549
; 
32'd177684: dataIn1 = 32'd8553
; 
32'd177685: dataIn1 = 32'd8556
; 
32'd177686: dataIn1 = 32'd8557
; 
32'd177687: dataIn1 = 32'd8567
; 
32'd177688: dataIn1 = 32'd5240
; 
32'd177689: dataIn1 = 32'd6502
; 
32'd177690: dataIn1 = 32'd8542
; 
32'd177691: dataIn1 = 32'd8553
; 
32'd177692: dataIn1 = 32'd8556
; 
32'd177693: dataIn1 = 32'd8557
; 
32'd177694: dataIn1 = 32'd8562
; 
32'd177695: dataIn1 = 32'd5229
; 
32'd177696: dataIn1 = 32'd6503
; 
32'd177697: dataIn1 = 32'd8393
; 
32'd177698: dataIn1 = 32'd8554
; 
32'd177699: dataIn1 = 32'd8558
; 
32'd177700: dataIn1 = 32'd8559
; 
32'd177701: dataIn1 = 32'd8568
; 
32'd177702: dataIn1 = 32'd5229
; 
32'd177703: dataIn1 = 32'd6501
; 
32'd177704: dataIn1 = 32'd6775
; 
32'd177705: dataIn1 = 32'd8554
; 
32'd177706: dataIn1 = 32'd8558
; 
32'd177707: dataIn1 = 32'd8559
; 
32'd177708: dataIn1 = 32'd5243
; 
32'd177709: dataIn1 = 32'd6502
; 
32'd177710: dataIn1 = 32'd8555
; 
32'd177711: dataIn1 = 32'd8560
; 
32'd177712: dataIn1 = 32'd8561
; 
32'd177713: dataIn1 = 32'd8564
; 
32'd177714: dataIn1 = 32'd8566
; 
32'd177715: dataIn1 = 32'd5243
; 
32'd177716: dataIn1 = 32'd6501
; 
32'd177717: dataIn1 = 32'd6774
; 
32'd177718: dataIn1 = 32'd8555
; 
32'd177719: dataIn1 = 32'd8560
; 
32'd177720: dataIn1 = 32'd8561
; 
32'd177721: dataIn1 = 32'd6498
; 
32'd177722: dataIn1 = 32'd6502
; 
32'd177723: dataIn1 = 32'd8542
; 
32'd177724: dataIn1 = 32'd8557
; 
32'd177725: dataIn1 = 32'd8562
; 
32'd177726: dataIn1 = 32'd8563
; 
32'd177727: dataIn1 = 32'd8564
; 
32'd177728: dataIn1 = 32'd6498
; 
32'd177729: dataIn1 = 32'd6504
; 
32'd177730: dataIn1 = 32'd8543
; 
32'd177731: dataIn1 = 32'd8562
; 
32'd177732: dataIn1 = 32'd8563
; 
32'd177733: dataIn1 = 32'd8564
; 
32'd177734: dataIn1 = 32'd8565
; 
32'd177735: dataIn1 = 32'd6502
; 
32'd177736: dataIn1 = 32'd6504
; 
32'd177737: dataIn1 = 32'd8560
; 
32'd177738: dataIn1 = 32'd8562
; 
32'd177739: dataIn1 = 32'd8563
; 
32'd177740: dataIn1 = 32'd8564
; 
32'd177741: dataIn1 = 32'd8566
; 
32'd177742: dataIn1 = 32'd2728
; 
32'd177743: dataIn1 = 32'd6504
; 
32'd177744: dataIn1 = 32'd8543
; 
32'd177745: dataIn1 = 32'd8563
; 
32'd177746: dataIn1 = 32'd8565
; 
32'd177747: dataIn1 = 32'd9195
; 
32'd177748: dataIn1 = 32'd9228
; 
32'd177749: dataIn1 = 32'd5243
; 
32'd177750: dataIn1 = 32'd6504
; 
32'd177751: dataIn1 = 32'd8560
; 
32'd177752: dataIn1 = 32'd8564
; 
32'd177753: dataIn1 = 32'd8566
; 
32'd177754: dataIn1 = 32'd9227
; 
32'd177755: dataIn1 = 32'd9230
; 
32'd177756: dataIn1 = 32'd6500
; 
32'd177757: dataIn1 = 32'd6503
; 
32'd177758: dataIn1 = 32'd8549
; 
32'd177759: dataIn1 = 32'd8556
; 
32'd177760: dataIn1 = 32'd8567
; 
32'd177761: dataIn1 = 32'd8568
; 
32'd177762: dataIn1 = 32'd8569
; 
32'd177763: dataIn1 = 32'd6460
; 
32'd177764: dataIn1 = 32'd6503
; 
32'd177765: dataIn1 = 32'd8393
; 
32'd177766: dataIn1 = 32'd8558
; 
32'd177767: dataIn1 = 32'd8567
; 
32'd177768: dataIn1 = 32'd8568
; 
32'd177769: dataIn1 = 32'd8569
; 
32'd177770: dataIn1 = 32'd6460
; 
32'd177771: dataIn1 = 32'd6500
; 
32'd177772: dataIn1 = 32'd8394
; 
32'd177773: dataIn1 = 32'd8551
; 
32'd177774: dataIn1 = 32'd8567
; 
32'd177775: dataIn1 = 32'd8568
; 
32'd177776: dataIn1 = 32'd8569
; 
32'd177777: dataIn1 = 32'd6506
; 
32'd177778: dataIn1 = 32'd6507
; 
32'd177779: dataIn1 = 32'd8570
; 
32'd177780: dataIn1 = 32'd8571
; 
32'd177781: dataIn1 = 32'd8572
; 
32'd177782: dataIn1 = 32'd8573
; 
32'd177783: dataIn1 = 32'd8574
; 
32'd177784: dataIn1 = 32'd6505
; 
32'd177785: dataIn1 = 32'd6507
; 
32'd177786: dataIn1 = 32'd8570
; 
32'd177787: dataIn1 = 32'd8571
; 
32'd177788: dataIn1 = 32'd8572
; 
32'd177789: dataIn1 = 32'd8575
; 
32'd177790: dataIn1 = 32'd8576
; 
32'd177791: dataIn1 = 32'd6505
; 
32'd177792: dataIn1 = 32'd6506
; 
32'd177793: dataIn1 = 32'd8570
; 
32'd177794: dataIn1 = 32'd8571
; 
32'd177795: dataIn1 = 32'd8572
; 
32'd177796: dataIn1 = 32'd8577
; 
32'd177797: dataIn1 = 32'd8578
; 
32'd177798: dataIn1 = 32'd5231
; 
32'd177799: dataIn1 = 32'd6507
; 
32'd177800: dataIn1 = 32'd8419
; 
32'd177801: dataIn1 = 32'd8570
; 
32'd177802: dataIn1 = 32'd8573
; 
32'd177803: dataIn1 = 32'd8574
; 
32'd177804: dataIn1 = 32'd8589
; 
32'd177805: dataIn1 = 32'd5231
; 
32'd177806: dataIn1 = 32'd6506
; 
32'd177807: dataIn1 = 32'd8412
; 
32'd177808: dataIn1 = 32'd8570
; 
32'd177809: dataIn1 = 32'd8573
; 
32'd177810: dataIn1 = 32'd8574
; 
32'd177811: dataIn1 = 32'd8584
; 
32'd177812: dataIn1 = 32'd5241
; 
32'd177813: dataIn1 = 32'd6507
; 
32'd177814: dataIn1 = 32'd8550
; 
32'd177815: dataIn1 = 32'd8571
; 
32'd177816: dataIn1 = 32'd8575
; 
32'd177817: dataIn1 = 32'd8576
; 
32'd177818: dataIn1 = 32'd8590
; 
32'd177819: dataIn1 = 32'd5241
; 
32'd177820: dataIn1 = 32'd6505
; 
32'd177821: dataIn1 = 32'd8537
; 
32'd177822: dataIn1 = 32'd8571
; 
32'd177823: dataIn1 = 32'd8575
; 
32'd177824: dataIn1 = 32'd8576
; 
32'd177825: dataIn1 = 32'd8580
; 
32'd177826: dataIn1 = 32'd2680
; 
32'd177827: dataIn1 = 32'd6506
; 
32'd177828: dataIn1 = 32'd8572
; 
32'd177829: dataIn1 = 32'd8577
; 
32'd177830: dataIn1 = 32'd8578
; 
32'd177831: dataIn1 = 32'd8586
; 
32'd177832: dataIn1 = 32'd8588
; 
32'd177833: dataIn1 = 32'd2680
; 
32'd177834: dataIn1 = 32'd6505
; 
32'd177835: dataIn1 = 32'd8572
; 
32'd177836: dataIn1 = 32'd8577
; 
32'd177837: dataIn1 = 32'd8578
; 
32'd177838: dataIn1 = 32'd8581
; 
32'd177839: dataIn1 = 32'd8583
; 
32'd177840: dataIn1 = 32'd5068
; 
32'd177841: dataIn1 = 32'd6496
; 
32'd177842: dataIn1 = 32'd8535
; 
32'd177843: dataIn1 = 32'd8579
; 
32'd177844: dataIn1 = 32'd8580
; 
32'd177845: dataIn1 = 32'd8581
; 
32'd177846: dataIn1 = 32'd8582
; 
32'd177847: dataIn1 = 32'd6496
; 
32'd177848: dataIn1 = 32'd6505
; 
32'd177849: dataIn1 = 32'd8537
; 
32'd177850: dataIn1 = 32'd8576
; 
32'd177851: dataIn1 = 32'd8579
; 
32'd177852: dataIn1 = 32'd8580
; 
32'd177853: dataIn1 = 32'd8581
; 
32'd177854: dataIn1 = 32'd5068
; 
32'd177855: dataIn1 = 32'd6505
; 
32'd177856: dataIn1 = 32'd8578
; 
32'd177857: dataIn1 = 32'd8579
; 
32'd177858: dataIn1 = 32'd8580
; 
32'd177859: dataIn1 = 32'd8581
; 
32'd177860: dataIn1 = 32'd8583
; 
32'd177861: dataIn1 = 32'd1116
; 
32'd177862: dataIn1 = 32'd5061
; 
32'd177863: dataIn1 = 32'd5068
; 
32'd177864: dataIn1 = 32'd8535
; 
32'd177865: dataIn1 = 32'd8579
; 
32'd177866: dataIn1 = 32'd8582
; 
32'd177867: dataIn1 = 32'd2680
; 
32'd177868: dataIn1 = 32'd5065
; 
32'd177869: dataIn1 = 32'd5068
; 
32'd177870: dataIn1 = 32'd8578
; 
32'd177871: dataIn1 = 32'd8581
; 
32'd177872: dataIn1 = 32'd8583
; 
32'd177873: dataIn1 = 32'd6467
; 
32'd177874: dataIn1 = 32'd6506
; 
32'd177875: dataIn1 = 32'd8412
; 
32'd177876: dataIn1 = 32'd8574
; 
32'd177877: dataIn1 = 32'd8584
; 
32'd177878: dataIn1 = 32'd8585
; 
32'd177879: dataIn1 = 32'd8586
; 
32'd177880: dataIn1 = 32'd5067
; 
32'd177881: dataIn1 = 32'd6467
; 
32'd177882: dataIn1 = 32'd8413
; 
32'd177883: dataIn1 = 32'd8584
; 
32'd177884: dataIn1 = 32'd8585
; 
32'd177885: dataIn1 = 32'd8586
; 
32'd177886: dataIn1 = 32'd8587
; 
32'd177887: dataIn1 = 32'd5067
; 
32'd177888: dataIn1 = 32'd6506
; 
32'd177889: dataIn1 = 32'd8577
; 
32'd177890: dataIn1 = 32'd8584
; 
32'd177891: dataIn1 = 32'd8585
; 
32'd177892: dataIn1 = 32'd8586
; 
32'd177893: dataIn1 = 32'd8588
; 
32'd177894: dataIn1 = 32'd145
; 
32'd177895: dataIn1 = 32'd4760
; 
32'd177896: dataIn1 = 32'd5067
; 
32'd177897: dataIn1 = 32'd8413
; 
32'd177898: dataIn1 = 32'd8585
; 
32'd177899: dataIn1 = 32'd8587
; 
32'd177900: dataIn1 = 32'd2680
; 
32'd177901: dataIn1 = 32'd5064
; 
32'd177902: dataIn1 = 32'd5067
; 
32'd177903: dataIn1 = 32'd8577
; 
32'd177904: dataIn1 = 32'd8586
; 
32'd177905: dataIn1 = 32'd8588
; 
32'd177906: dataIn1 = 32'd6468
; 
32'd177907: dataIn1 = 32'd6507
; 
32'd177908: dataIn1 = 32'd8419
; 
32'd177909: dataIn1 = 32'd8573
; 
32'd177910: dataIn1 = 32'd8589
; 
32'd177911: dataIn1 = 32'd8590
; 
32'd177912: dataIn1 = 32'd8591
; 
32'd177913: dataIn1 = 32'd6499
; 
32'd177914: dataIn1 = 32'd6507
; 
32'd177915: dataIn1 = 32'd8550
; 
32'd177916: dataIn1 = 32'd8575
; 
32'd177917: dataIn1 = 32'd8589
; 
32'd177918: dataIn1 = 32'd8590
; 
32'd177919: dataIn1 = 32'd8591
; 
32'd177920: dataIn1 = 32'd6468
; 
32'd177921: dataIn1 = 32'd6499
; 
32'd177922: dataIn1 = 32'd8420
; 
32'd177923: dataIn1 = 32'd8552
; 
32'd177924: dataIn1 = 32'd8589
; 
32'd177925: dataIn1 = 32'd8590
; 
32'd177926: dataIn1 = 32'd8591
; 
32'd177927: dataIn1 = 32'd6509
; 
32'd177928: dataIn1 = 32'd6510
; 
32'd177929: dataIn1 = 32'd8592
; 
32'd177930: dataIn1 = 32'd8593
; 
32'd177931: dataIn1 = 32'd8594
; 
32'd177932: dataIn1 = 32'd8595
; 
32'd177933: dataIn1 = 32'd8596
; 
32'd177934: dataIn1 = 32'd6508
; 
32'd177935: dataIn1 = 32'd6510
; 
32'd177936: dataIn1 = 32'd8592
; 
32'd177937: dataIn1 = 32'd8593
; 
32'd177938: dataIn1 = 32'd8594
; 
32'd177939: dataIn1 = 32'd8597
; 
32'd177940: dataIn1 = 32'd8598
; 
32'd177941: dataIn1 = 32'd6508
; 
32'd177942: dataIn1 = 32'd6509
; 
32'd177943: dataIn1 = 32'd8592
; 
32'd177944: dataIn1 = 32'd8593
; 
32'd177945: dataIn1 = 32'd8594
; 
32'd177946: dataIn1 = 32'd8599
; 
32'd177947: dataIn1 = 32'd8600
; 
32'd177948: dataIn1 = 32'd5244
; 
32'd177949: dataIn1 = 32'd6510
; 
32'd177950: dataIn1 = 32'd8592
; 
32'd177951: dataIn1 = 32'd8595
; 
32'd177952: dataIn1 = 32'd8596
; 
32'd177953: dataIn1 = 32'd8611
; 
32'd177954: dataIn1 = 32'd8614
; 
32'd177955: dataIn1 = 32'd5244
; 
32'd177956: dataIn1 = 32'd6509
; 
32'd177957: dataIn1 = 32'd8592
; 
32'd177958: dataIn1 = 32'd8595
; 
32'd177959: dataIn1 = 32'd8596
; 
32'd177960: dataIn1 = 32'd8606
; 
32'd177961: dataIn1 = 32'd8609
; 
32'd177962: dataIn1 = 32'd2681
; 
32'd177963: dataIn1 = 32'd6510
; 
32'd177964: dataIn1 = 32'd8593
; 
32'd177965: dataIn1 = 32'd8597
; 
32'd177966: dataIn1 = 32'd8598
; 
32'd177967: dataIn1 = 32'd8612
; 
32'd177968: dataIn1 = 32'd8615
; 
32'd177969: dataIn1 = 32'd2681
; 
32'd177970: dataIn1 = 32'd6508
; 
32'd177971: dataIn1 = 32'd8593
; 
32'd177972: dataIn1 = 32'd8597
; 
32'd177973: dataIn1 = 32'd8598
; 
32'd177974: dataIn1 = 32'd8602
; 
32'd177975: dataIn1 = 32'd8605
; 
32'd177976: dataIn1 = 32'd5242
; 
32'd177977: dataIn1 = 32'd6509
; 
32'd177978: dataIn1 = 32'd8545
; 
32'd177979: dataIn1 = 32'd8594
; 
32'd177980: dataIn1 = 32'd8599
; 
32'd177981: dataIn1 = 32'd8600
; 
32'd177982: dataIn1 = 32'd8608
; 
32'd177983: dataIn1 = 32'd5242
; 
32'd177984: dataIn1 = 32'd6508
; 
32'd177985: dataIn1 = 32'd8538
; 
32'd177986: dataIn1 = 32'd8594
; 
32'd177987: dataIn1 = 32'd8599
; 
32'd177988: dataIn1 = 32'd8600
; 
32'd177989: dataIn1 = 32'd8603
; 
32'd177990: dataIn1 = 32'd5072
; 
32'd177991: dataIn1 = 32'd6495
; 
32'd177992: dataIn1 = 32'd8536
; 
32'd177993: dataIn1 = 32'd8601
; 
32'd177994: dataIn1 = 32'd8602
; 
32'd177995: dataIn1 = 32'd8603
; 
32'd177996: dataIn1 = 32'd8604
; 
32'd177997: dataIn1 = 32'd5072
; 
32'd177998: dataIn1 = 32'd6508
; 
32'd177999: dataIn1 = 32'd8598
; 
32'd178000: dataIn1 = 32'd8601
; 
32'd178001: dataIn1 = 32'd8602
; 
32'd178002: dataIn1 = 32'd8603
; 
32'd178003: dataIn1 = 32'd8605
; 
32'd178004: dataIn1 = 32'd6495
; 
32'd178005: dataIn1 = 32'd6508
; 
32'd178006: dataIn1 = 32'd8538
; 
32'd178007: dataIn1 = 32'd8600
; 
32'd178008: dataIn1 = 32'd8601
; 
32'd178009: dataIn1 = 32'd8602
; 
32'd178010: dataIn1 = 32'd8603
; 
32'd178011: dataIn1 = 32'd1116
; 
32'd178012: dataIn1 = 32'd5060
; 
32'd178013: dataIn1 = 32'd5072
; 
32'd178014: dataIn1 = 32'd8536
; 
32'd178015: dataIn1 = 32'd8601
; 
32'd178016: dataIn1 = 32'd8604
; 
32'd178017: dataIn1 = 32'd2681
; 
32'd178018: dataIn1 = 32'd5070
; 
32'd178019: dataIn1 = 32'd5072
; 
32'd178020: dataIn1 = 32'd8598
; 
32'd178021: dataIn1 = 32'd8602
; 
32'd178022: dataIn1 = 32'd8605
; 
32'd178023: dataIn1 = 32'd6509
; 
32'd178024: dataIn1 = 32'd6511
; 
32'd178025: dataIn1 = 32'd8596
; 
32'd178026: dataIn1 = 32'd8606
; 
32'd178027: dataIn1 = 32'd8607
; 
32'd178028: dataIn1 = 32'd8608
; 
32'd178029: dataIn1 = 32'd8609
; 
32'd178030: dataIn1 = 32'd6497
; 
32'd178031: dataIn1 = 32'd6511
; 
32'd178032: dataIn1 = 32'd8544
; 
32'd178033: dataIn1 = 32'd8606
; 
32'd178034: dataIn1 = 32'd8607
; 
32'd178035: dataIn1 = 32'd8608
; 
32'd178036: dataIn1 = 32'd8610
; 
32'd178037: dataIn1 = 32'd6497
; 
32'd178038: dataIn1 = 32'd6509
; 
32'd178039: dataIn1 = 32'd8545
; 
32'd178040: dataIn1 = 32'd8599
; 
32'd178041: dataIn1 = 32'd8606
; 
32'd178042: dataIn1 = 32'd8607
; 
32'd178043: dataIn1 = 32'd8608
; 
32'd178044: dataIn1 = 32'd5244
; 
32'd178045: dataIn1 = 32'd6511
; 
32'd178046: dataIn1 = 32'd8596
; 
32'd178047: dataIn1 = 32'd8606
; 
32'd178048: dataIn1 = 32'd8609
; 
32'd178049: dataIn1 = 32'd9211
; 
32'd178050: dataIn1 = 32'd9218
; 
32'd178051: dataIn1 = 32'd2728
; 
32'd178052: dataIn1 = 32'd6511
; 
32'd178053: dataIn1 = 32'd8544
; 
32'd178054: dataIn1 = 32'd8607
; 
32'd178055: dataIn1 = 32'd8610
; 
32'd178056: dataIn1 = 32'd9194
; 
32'd178057: dataIn1 = 32'd9217
; 
32'd178058: dataIn1 = 32'd6510
; 
32'd178059: dataIn1 = 32'd6512
; 
32'd178060: dataIn1 = 32'd8595
; 
32'd178061: dataIn1 = 32'd8611
; 
32'd178062: dataIn1 = 32'd8612
; 
32'd178063: dataIn1 = 32'd8613
; 
32'd178064: dataIn1 = 32'd8614
; 
32'd178065: dataIn1 = 32'd5073
; 
32'd178066: dataIn1 = 32'd6510
; 
32'd178067: dataIn1 = 32'd8597
; 
32'd178068: dataIn1 = 32'd8611
; 
32'd178069: dataIn1 = 32'd8612
; 
32'd178070: dataIn1 = 32'd8613
; 
32'd178071: dataIn1 = 32'd8615
; 
32'd178072: dataIn1 = 32'd5073
; 
32'd178073: dataIn1 = 32'd6512
; 
32'd178074: dataIn1 = 32'd8611
; 
32'd178075: dataIn1 = 32'd8612
; 
32'd178076: dataIn1 = 32'd8613
; 
32'd178077: dataIn1 = 32'd8616
; 
32'd178078: dataIn1 = 32'd8617
; 
32'd178079: dataIn1 = 32'd5244
; 
32'd178080: dataIn1 = 32'd6512
; 
32'd178081: dataIn1 = 32'd8595
; 
32'd178082: dataIn1 = 32'd8611
; 
32'd178083: dataIn1 = 32'd8614
; 
32'd178084: dataIn1 = 32'd9212
; 
32'd178085: dataIn1 = 32'd9215
; 
32'd178086: dataIn1 = 32'd2681
; 
32'd178087: dataIn1 = 32'd5071
; 
32'd178088: dataIn1 = 32'd5073
; 
32'd178089: dataIn1 = 32'd8597
; 
32'd178090: dataIn1 = 32'd8612
; 
32'd178091: dataIn1 = 32'd8615
; 
32'd178092: dataIn1 = 32'd11
; 
32'd178093: dataIn1 = 32'd6512
; 
32'd178094: dataIn1 = 32'd8613
; 
32'd178095: dataIn1 = 32'd8616
; 
32'd178096: dataIn1 = 32'd8617
; 
32'd178097: dataIn1 = 32'd8724
; 
32'd178098: dataIn1 = 32'd9213
; 
32'd178099: dataIn1 = 32'd11
; 
32'd178100: dataIn1 = 32'd4770
; 
32'd178101: dataIn1 = 32'd5073
; 
32'd178102: dataIn1 = 32'd8613
; 
32'd178103: dataIn1 = 32'd8616
; 
32'd178104: dataIn1 = 32'd8617
; 
32'd178105: dataIn1 = 32'd6514
; 
32'd178106: dataIn1 = 32'd6515
; 
32'd178107: dataIn1 = 32'd8618
; 
32'd178108: dataIn1 = 32'd8619
; 
32'd178109: dataIn1 = 32'd8620
; 
32'd178110: dataIn1 = 32'd8621
; 
32'd178111: dataIn1 = 32'd8622
; 
32'd178112: dataIn1 = 32'd6513
; 
32'd178113: dataIn1 = 32'd6515
; 
32'd178114: dataIn1 = 32'd8618
; 
32'd178115: dataIn1 = 32'd8619
; 
32'd178116: dataIn1 = 32'd8620
; 
32'd178117: dataIn1 = 32'd8623
; 
32'd178118: dataIn1 = 32'd8624
; 
32'd178119: dataIn1 = 32'd6513
; 
32'd178120: dataIn1 = 32'd6514
; 
32'd178121: dataIn1 = 32'd8618
; 
32'd178122: dataIn1 = 32'd8619
; 
32'd178123: dataIn1 = 32'd8620
; 
32'd178124: dataIn1 = 32'd8625
; 
32'd178125: dataIn1 = 32'd8626
; 
32'd178126: dataIn1 = 32'd5245
; 
32'd178127: dataIn1 = 32'd6515
; 
32'd178128: dataIn1 = 32'd8618
; 
32'd178129: dataIn1 = 32'd8621
; 
32'd178130: dataIn1 = 32'd8622
; 
32'd178131: dataIn1 = 32'd8634
; 
32'd178132: dataIn1 = 32'd8637
; 
32'd178133: dataIn1 = 32'd5245
; 
32'd178134: dataIn1 = 32'd6514
; 
32'd178135: dataIn1 = 32'd6777
; 
32'd178136: dataIn1 = 32'd8618
; 
32'd178137: dataIn1 = 32'd8621
; 
32'd178138: dataIn1 = 32'd8622
; 
32'd178139: dataIn1 = 32'd5246
; 
32'd178140: dataIn1 = 32'd6515
; 
32'd178141: dataIn1 = 32'd8619
; 
32'd178142: dataIn1 = 32'd8623
; 
32'd178143: dataIn1 = 32'd8624
; 
32'd178144: dataIn1 = 32'd8635
; 
32'd178145: dataIn1 = 32'd8638
; 
32'd178146: dataIn1 = 32'd5246
; 
32'd178147: dataIn1 = 32'd6513
; 
32'd178148: dataIn1 = 32'd8619
; 
32'd178149: dataIn1 = 32'd8623
; 
32'd178150: dataIn1 = 32'd8624
; 
32'd178151: dataIn1 = 32'd8628
; 
32'd178152: dataIn1 = 32'd8632
; 
32'd178153: dataIn1 = 32'd5247
; 
32'd178154: dataIn1 = 32'd6514
; 
32'd178155: dataIn1 = 32'd6776
; 
32'd178156: dataIn1 = 32'd8620
; 
32'd178157: dataIn1 = 32'd8625
; 
32'd178158: dataIn1 = 32'd8626
; 
32'd178159: dataIn1 = 32'd5247
; 
32'd178160: dataIn1 = 32'd6513
; 
32'd178161: dataIn1 = 32'd8620
; 
32'd178162: dataIn1 = 32'd8625
; 
32'd178163: dataIn1 = 32'd8626
; 
32'd178164: dataIn1 = 32'd8629
; 
32'd178165: dataIn1 = 32'd8633
; 
32'd178166: dataIn1 = 32'd6516
; 
32'd178167: dataIn1 = 32'd6517
; 
32'd178168: dataIn1 = 32'd8627
; 
32'd178169: dataIn1 = 32'd8628
; 
32'd178170: dataIn1 = 32'd8629
; 
32'd178171: dataIn1 = 32'd8630
; 
32'd178172: dataIn1 = 32'd8631
; 
32'd178173: dataIn1 = 32'd6513
; 
32'd178174: dataIn1 = 32'd6517
; 
32'd178175: dataIn1 = 32'd8624
; 
32'd178176: dataIn1 = 32'd8627
; 
32'd178177: dataIn1 = 32'd8628
; 
32'd178178: dataIn1 = 32'd8629
; 
32'd178179: dataIn1 = 32'd8632
; 
32'd178180: dataIn1 = 32'd6513
; 
32'd178181: dataIn1 = 32'd6516
; 
32'd178182: dataIn1 = 32'd8626
; 
32'd178183: dataIn1 = 32'd8627
; 
32'd178184: dataIn1 = 32'd8628
; 
32'd178185: dataIn1 = 32'd8629
; 
32'd178186: dataIn1 = 32'd8633
; 
32'd178187: dataIn1 = 32'd2729
; 
32'd178188: dataIn1 = 32'd6517
; 
32'd178189: dataIn1 = 32'd8627
; 
32'd178190: dataIn1 = 32'd8630
; 
32'd178191: dataIn1 = 32'd8631
; 
32'd178192: dataIn1 = 32'd8657
; 
32'd178193: dataIn1 = 32'd8660
; 
32'd178194: dataIn1 = 32'd2729
; 
32'd178195: dataIn1 = 32'd6516
; 
32'd178196: dataIn1 = 32'd8627
; 
32'd178197: dataIn1 = 32'd8630
; 
32'd178198: dataIn1 = 32'd8631
; 
32'd178199: dataIn1 = 32'd8674
; 
32'd178200: dataIn1 = 32'd8677
; 
32'd178201: dataIn1 = 32'd5246
; 
32'd178202: dataIn1 = 32'd6517
; 
32'd178203: dataIn1 = 32'd8624
; 
32'd178204: dataIn1 = 32'd8628
; 
32'd178205: dataIn1 = 32'd8632
; 
32'd178206: dataIn1 = 32'd8654
; 
32'd178207: dataIn1 = 32'd8658
; 
32'd178208: dataIn1 = 32'd5247
; 
32'd178209: dataIn1 = 32'd6516
; 
32'd178210: dataIn1 = 32'd8626
; 
32'd178211: dataIn1 = 32'd8629
; 
32'd178212: dataIn1 = 32'd8633
; 
32'd178213: dataIn1 = 32'd8676
; 
32'd178214: dataIn1 = 32'd8680
; 
32'd178215: dataIn1 = 32'd6515
; 
32'd178216: dataIn1 = 32'd6519
; 
32'd178217: dataIn1 = 32'd8621
; 
32'd178218: dataIn1 = 32'd8634
; 
32'd178219: dataIn1 = 32'd8635
; 
32'd178220: dataIn1 = 32'd8636
; 
32'd178221: dataIn1 = 32'd8637
; 
32'd178222: dataIn1 = 32'd6515
; 
32'd178223: dataIn1 = 32'd6518
; 
32'd178224: dataIn1 = 32'd8623
; 
32'd178225: dataIn1 = 32'd8634
; 
32'd178226: dataIn1 = 32'd8635
; 
32'd178227: dataIn1 = 32'd8636
; 
32'd178228: dataIn1 = 32'd8638
; 
32'd178229: dataIn1 = 32'd6518
; 
32'd178230: dataIn1 = 32'd6519
; 
32'd178231: dataIn1 = 32'd8634
; 
32'd178232: dataIn1 = 32'd8635
; 
32'd178233: dataIn1 = 32'd8636
; 
32'd178234: dataIn1 = 32'd8639
; 
32'd178235: dataIn1 = 32'd8640
; 
32'd178236: dataIn1 = 32'd5245
; 
32'd178237: dataIn1 = 32'd6519
; 
32'd178238: dataIn1 = 32'd8621
; 
32'd178239: dataIn1 = 32'd8634
; 
32'd178240: dataIn1 = 32'd8637
; 
32'd178241: dataIn1 = 32'd8641
; 
32'd178242: dataIn1 = 32'd8644
; 
32'd178243: dataIn1 = 32'd5246
; 
32'd178244: dataIn1 = 32'd6518
; 
32'd178245: dataIn1 = 32'd8623
; 
32'd178246: dataIn1 = 32'd8635
; 
32'd178247: dataIn1 = 32'd8638
; 
32'd178248: dataIn1 = 32'd8653
; 
32'd178249: dataIn1 = 32'd8670
; 
32'd178250: dataIn1 = 32'd2731
; 
32'd178251: dataIn1 = 32'd6519
; 
32'd178252: dataIn1 = 32'd8636
; 
32'd178253: dataIn1 = 32'd8639
; 
32'd178254: dataIn1 = 32'd8640
; 
32'd178255: dataIn1 = 32'd8643
; 
32'd178256: dataIn1 = 32'd8647
; 
32'd178257: dataIn1 = 32'd2731
; 
32'd178258: dataIn1 = 32'd6518
; 
32'd178259: dataIn1 = 32'd8636
; 
32'd178260: dataIn1 = 32'd8639
; 
32'd178261: dataIn1 = 32'd8640
; 
32'd178262: dataIn1 = 32'd8671
; 
32'd178263: dataIn1 = 32'd8673
; 
32'd178264: dataIn1 = 32'd6519
; 
32'd178265: dataIn1 = 32'd6521
; 
32'd178266: dataIn1 = 32'd8637
; 
32'd178267: dataIn1 = 32'd8641
; 
32'd178268: dataIn1 = 32'd8642
; 
32'd178269: dataIn1 = 32'd8643
; 
32'd178270: dataIn1 = 32'd8644
; 
32'd178271: dataIn1 = 32'd6520
; 
32'd178272: dataIn1 = 32'd6521
; 
32'd178273: dataIn1 = 32'd8641
; 
32'd178274: dataIn1 = 32'd8642
; 
32'd178275: dataIn1 = 32'd8643
; 
32'd178276: dataIn1 = 32'd8645
; 
32'd178277: dataIn1 = 32'd8646
; 
32'd178278: dataIn1 = 32'd6519
; 
32'd178279: dataIn1 = 32'd6520
; 
32'd178280: dataIn1 = 32'd8639
; 
32'd178281: dataIn1 = 32'd8641
; 
32'd178282: dataIn1 = 32'd8642
; 
32'd178283: dataIn1 = 32'd8643
; 
32'd178284: dataIn1 = 32'd8647
; 
32'd178285: dataIn1 = 32'd5245
; 
32'd178286: dataIn1 = 32'd6521
; 
32'd178287: dataIn1 = 32'd6779
; 
32'd178288: dataIn1 = 32'd8637
; 
32'd178289: dataIn1 = 32'd8641
; 
32'd178290: dataIn1 = 32'd8644
; 
32'd178291: dataIn1 = 32'd5248
; 
32'd178292: dataIn1 = 32'd6521
; 
32'd178293: dataIn1 = 32'd6778
; 
32'd178294: dataIn1 = 32'd8642
; 
32'd178295: dataIn1 = 32'd8645
; 
32'd178296: dataIn1 = 32'd8646
; 
32'd178297: dataIn1 = 32'd5248
; 
32'd178298: dataIn1 = 32'd6520
; 
32'd178299: dataIn1 = 32'd8642
; 
32'd178300: dataIn1 = 32'd8645
; 
32'd178301: dataIn1 = 32'd8646
; 
32'd178302: dataIn1 = 32'd8811
; 
32'd178303: dataIn1 = 32'd8820
; 
32'd178304: dataIn1 = 32'd2731
; 
32'd178305: dataIn1 = 32'd6520
; 
32'd178306: dataIn1 = 32'd8639
; 
32'd178307: dataIn1 = 32'd8643
; 
32'd178308: dataIn1 = 32'd8647
; 
32'd178309: dataIn1 = 32'd8804
; 
32'd178310: dataIn1 = 32'd8821
; 
32'd178311: dataIn1 = 32'd6523
; 
32'd178312: dataIn1 = 32'd6524
; 
32'd178313: dataIn1 = 32'd8648
; 
32'd178314: dataIn1 = 32'd8649
; 
32'd178315: dataIn1 = 32'd8650
; 
32'd178316: dataIn1 = 32'd8651
; 
32'd178317: dataIn1 = 32'd8652
; 
32'd178318: dataIn1 = 32'd6522
; 
32'd178319: dataIn1 = 32'd6524
; 
32'd178320: dataIn1 = 32'd8648
; 
32'd178321: dataIn1 = 32'd8649
; 
32'd178322: dataIn1 = 32'd8650
; 
32'd178323: dataIn1 = 32'd8653
; 
32'd178324: dataIn1 = 32'd8654
; 
32'd178325: dataIn1 = 32'd6522
; 
32'd178326: dataIn1 = 32'd6523
; 
32'd178327: dataIn1 = 32'd8648
; 
32'd178328: dataIn1 = 32'd8649
; 
32'd178329: dataIn1 = 32'd8650
; 
32'd178330: dataIn1 = 32'd8655
; 
32'd178331: dataIn1 = 32'd8656
; 
32'd178332: dataIn1 = 32'd5250
; 
32'd178333: dataIn1 = 32'd6524
; 
32'd178334: dataIn1 = 32'd8648
; 
32'd178335: dataIn1 = 32'd8651
; 
32'd178336: dataIn1 = 32'd8652
; 
32'd178337: dataIn1 = 32'd8669
; 
32'd178338: dataIn1 = 32'd8672
; 
32'd178339: dataIn1 = 32'd5250
; 
32'd178340: dataIn1 = 32'd6523
; 
32'd178341: dataIn1 = 32'd8648
; 
32'd178342: dataIn1 = 32'd8651
; 
32'd178343: dataIn1 = 32'd8652
; 
32'd178344: dataIn1 = 32'd8662
; 
32'd178345: dataIn1 = 32'd8665
; 
32'd178346: dataIn1 = 32'd5246
; 
32'd178347: dataIn1 = 32'd6524
; 
32'd178348: dataIn1 = 32'd8638
; 
32'd178349: dataIn1 = 32'd8649
; 
32'd178350: dataIn1 = 32'd8653
; 
32'd178351: dataIn1 = 32'd8654
; 
32'd178352: dataIn1 = 32'd8670
; 
32'd178353: dataIn1 = 32'd5246
; 
32'd178354: dataIn1 = 32'd6522
; 
32'd178355: dataIn1 = 32'd8632
; 
32'd178356: dataIn1 = 32'd8649
; 
32'd178357: dataIn1 = 32'd8653
; 
32'd178358: dataIn1 = 32'd8654
; 
32'd178359: dataIn1 = 32'd8658
; 
32'd178360: dataIn1 = 32'd5251
; 
32'd178361: dataIn1 = 32'd6523
; 
32'd178362: dataIn1 = 32'd8650
; 
32'd178363: dataIn1 = 32'd8655
; 
32'd178364: dataIn1 = 32'd8656
; 
32'd178365: dataIn1 = 32'd8664
; 
32'd178366: dataIn1 = 32'd8668
; 
32'd178367: dataIn1 = 32'd5251
; 
32'd178368: dataIn1 = 32'd6522
; 
32'd178369: dataIn1 = 32'd8650
; 
32'd178370: dataIn1 = 32'd8655
; 
32'd178371: dataIn1 = 32'd8656
; 
32'd178372: dataIn1 = 32'd8659
; 
32'd178373: dataIn1 = 32'd8661
; 
32'd178374: dataIn1 = 32'd6517
; 
32'd178375: dataIn1 = 32'd6525
; 
32'd178376: dataIn1 = 32'd8630
; 
32'd178377: dataIn1 = 32'd8657
; 
32'd178378: dataIn1 = 32'd8658
; 
32'd178379: dataIn1 = 32'd8659
; 
32'd178380: dataIn1 = 32'd8660
; 
32'd178381: dataIn1 = 32'd6517
; 
32'd178382: dataIn1 = 32'd6522
; 
32'd178383: dataIn1 = 32'd8632
; 
32'd178384: dataIn1 = 32'd8654
; 
32'd178385: dataIn1 = 32'd8657
; 
32'd178386: dataIn1 = 32'd8658
; 
32'd178387: dataIn1 = 32'd8659
; 
32'd178388: dataIn1 = 32'd6522
; 
32'd178389: dataIn1 = 32'd6525
; 
32'd178390: dataIn1 = 32'd8656
; 
32'd178391: dataIn1 = 32'd8657
; 
32'd178392: dataIn1 = 32'd8658
; 
32'd178393: dataIn1 = 32'd8659
; 
32'd178394: dataIn1 = 32'd8661
; 
32'd178395: dataIn1 = 32'd2729
; 
32'd178396: dataIn1 = 32'd6525
; 
32'd178397: dataIn1 = 32'd8630
; 
32'd178398: dataIn1 = 32'd8657
; 
32'd178399: dataIn1 = 32'd8660
; 
32'd178400: dataIn1 = 32'd8693
; 
32'd178401: dataIn1 = 32'd8746
; 
32'd178402: dataIn1 = 32'd5251
; 
32'd178403: dataIn1 = 32'd6525
; 
32'd178404: dataIn1 = 32'd8656
; 
32'd178405: dataIn1 = 32'd8659
; 
32'd178406: dataIn1 = 32'd8661
; 
32'd178407: dataIn1 = 32'd8745
; 
32'd178408: dataIn1 = 32'd8748
; 
32'd178409: dataIn1 = 32'd6523
; 
32'd178410: dataIn1 = 32'd6527
; 
32'd178411: dataIn1 = 32'd8652
; 
32'd178412: dataIn1 = 32'd8662
; 
32'd178413: dataIn1 = 32'd8663
; 
32'd178414: dataIn1 = 32'd8664
; 
32'd178415: dataIn1 = 32'd8665
; 
32'd178416: dataIn1 = 32'd6526
; 
32'd178417: dataIn1 = 32'd6527
; 
32'd178418: dataIn1 = 32'd8662
; 
32'd178419: dataIn1 = 32'd8663
; 
32'd178420: dataIn1 = 32'd8664
; 
32'd178421: dataIn1 = 32'd8666
; 
32'd178422: dataIn1 = 32'd8667
; 
32'd178423: dataIn1 = 32'd6523
; 
32'd178424: dataIn1 = 32'd6526
; 
32'd178425: dataIn1 = 32'd8655
; 
32'd178426: dataIn1 = 32'd8662
; 
32'd178427: dataIn1 = 32'd8663
; 
32'd178428: dataIn1 = 32'd8664
; 
32'd178429: dataIn1 = 32'd8668
; 
32'd178430: dataIn1 = 32'd5250
; 
32'd178431: dataIn1 = 32'd6527
; 
32'd178432: dataIn1 = 32'd8652
; 
32'd178433: dataIn1 = 32'd8662
; 
32'd178434: dataIn1 = 32'd8665
; 
32'd178435: dataIn1 = 32'd8826
; 
32'd178436: dataIn1 = 32'd8836
; 
32'd178437: dataIn1 = 32'd148
; 
32'd178438: dataIn1 = 32'd6527
; 
32'd178439: dataIn1 = 32'd8663
; 
32'd178440: dataIn1 = 32'd8666
; 
32'd178441: dataIn1 = 32'd8667
; 
32'd178442: dataIn1 = 32'd8837
; 
32'd178443: dataIn1 = 32'd8839
; 
32'd178444: dataIn1 = 32'd148
; 
32'd178445: dataIn1 = 32'd6526
; 
32'd178446: dataIn1 = 32'd8663
; 
32'd178447: dataIn1 = 32'd8666
; 
32'd178448: dataIn1 = 32'd8667
; 
32'd178449: dataIn1 = 32'd8750
; 
32'd178450: dataIn1 = 32'd8753
; 
32'd178451: dataIn1 = 32'd5251
; 
32'd178452: dataIn1 = 32'd6526
; 
32'd178453: dataIn1 = 32'd8655
; 
32'd178454: dataIn1 = 32'd8664
; 
32'd178455: dataIn1 = 32'd8668
; 
32'd178456: dataIn1 = 32'd8744
; 
32'd178457: dataIn1 = 32'd8751
; 
32'd178458: dataIn1 = 32'd6524
; 
32'd178459: dataIn1 = 32'd6528
; 
32'd178460: dataIn1 = 32'd8651
; 
32'd178461: dataIn1 = 32'd8669
; 
32'd178462: dataIn1 = 32'd8670
; 
32'd178463: dataIn1 = 32'd8671
; 
32'd178464: dataIn1 = 32'd8672
; 
32'd178465: dataIn1 = 32'd6518
; 
32'd178466: dataIn1 = 32'd6524
; 
32'd178467: dataIn1 = 32'd8638
; 
32'd178468: dataIn1 = 32'd8653
; 
32'd178469: dataIn1 = 32'd8669
; 
32'd178470: dataIn1 = 32'd8670
; 
32'd178471: dataIn1 = 32'd8671
; 
32'd178472: dataIn1 = 32'd6518
; 
32'd178473: dataIn1 = 32'd6528
; 
32'd178474: dataIn1 = 32'd8640
; 
32'd178475: dataIn1 = 32'd8669
; 
32'd178476: dataIn1 = 32'd8670
; 
32'd178477: dataIn1 = 32'd8671
; 
32'd178478: dataIn1 = 32'd8673
; 
32'd178479: dataIn1 = 32'd5250
; 
32'd178480: dataIn1 = 32'd6528
; 
32'd178481: dataIn1 = 32'd8651
; 
32'd178482: dataIn1 = 32'd8669
; 
32'd178483: dataIn1 = 32'd8672
; 
32'd178484: dataIn1 = 32'd8825
; 
32'd178485: dataIn1 = 32'd8841
; 
32'd178486: dataIn1 = 32'd2731
; 
32'd178487: dataIn1 = 32'd6528
; 
32'd178488: dataIn1 = 32'd8640
; 
32'd178489: dataIn1 = 32'd8671
; 
32'd178490: dataIn1 = 32'd8673
; 
32'd178491: dataIn1 = 32'd8805
; 
32'd178492: dataIn1 = 32'd8843
; 
32'd178493: dataIn1 = 32'd6516
; 
32'd178494: dataIn1 = 32'd6530
; 
32'd178495: dataIn1 = 32'd8631
; 
32'd178496: dataIn1 = 32'd8674
; 
32'd178497: dataIn1 = 32'd8675
; 
32'd178498: dataIn1 = 32'd8676
; 
32'd178499: dataIn1 = 32'd8677
; 
32'd178500: dataIn1 = 32'd6529
; 
32'd178501: dataIn1 = 32'd6530
; 
32'd178502: dataIn1 = 32'd8674
; 
32'd178503: dataIn1 = 32'd8675
; 
32'd178504: dataIn1 = 32'd8676
; 
32'd178505: dataIn1 = 32'd8678
; 
32'd178506: dataIn1 = 32'd8679
; 
32'd178507: dataIn1 = 32'd6516
; 
32'd178508: dataIn1 = 32'd6529
; 
32'd178509: dataIn1 = 32'd8633
; 
32'd178510: dataIn1 = 32'd8674
; 
32'd178511: dataIn1 = 32'd8675
; 
32'd178512: dataIn1 = 32'd8676
; 
32'd178513: dataIn1 = 32'd8680
; 
32'd178514: dataIn1 = 32'd2729
; 
32'd178515: dataIn1 = 32'd6530
; 
32'd178516: dataIn1 = 32'd8631
; 
32'd178517: dataIn1 = 32'd8674
; 
32'd178518: dataIn1 = 32'd8677
; 
32'd178519: dataIn1 = 32'd8694
; 
32'd178520: dataIn1 = 32'd8768
; 
32'd178521: dataIn1 = 32'd5253
; 
32'd178522: dataIn1 = 32'd6530
; 
32'd178523: dataIn1 = 32'd8675
; 
32'd178524: dataIn1 = 32'd8678
; 
32'd178525: dataIn1 = 32'd8679
; 
32'd178526: dataIn1 = 32'd8765
; 
32'd178527: dataIn1 = 32'd8769
; 
32'd178528: dataIn1 = 32'd5253
; 
32'd178529: dataIn1 = 32'd6529
; 
32'd178530: dataIn1 = 32'd6781
; 
32'd178531: dataIn1 = 32'd8675
; 
32'd178532: dataIn1 = 32'd8678
; 
32'd178533: dataIn1 = 32'd8679
; 
32'd178534: dataIn1 = 32'd5247
; 
32'd178535: dataIn1 = 32'd6529
; 
32'd178536: dataIn1 = 32'd6780
; 
32'd178537: dataIn1 = 32'd8633
; 
32'd178538: dataIn1 = 32'd8676
; 
32'd178539: dataIn1 = 32'd8680
; 
32'd178540: dataIn1 = 32'd6532
; 
32'd178541: dataIn1 = 32'd6533
; 
32'd178542: dataIn1 = 32'd8681
; 
32'd178543: dataIn1 = 32'd8682
; 
32'd178544: dataIn1 = 32'd8683
; 
32'd178545: dataIn1 = 32'd8684
; 
32'd178546: dataIn1 = 32'd8685
; 
32'd178547: dataIn1 = 32'd6531
; 
32'd178548: dataIn1 = 32'd6533
; 
32'd178549: dataIn1 = 32'd8681
; 
32'd178550: dataIn1 = 32'd8682
; 
32'd178551: dataIn1 = 32'd8683
; 
32'd178552: dataIn1 = 32'd8686
; 
32'd178553: dataIn1 = 32'd8687
; 
32'd178554: dataIn1 = 32'd6531
; 
32'd178555: dataIn1 = 32'd6532
; 
32'd178556: dataIn1 = 32'd8681
; 
32'd178557: dataIn1 = 32'd8682
; 
32'd178558: dataIn1 = 32'd8683
; 
32'd178559: dataIn1 = 32'd8688
; 
32'd178560: dataIn1 = 32'd8689
; 
32'd178561: dataIn1 = 32'd5254
; 
32'd178562: dataIn1 = 32'd6533
; 
32'd178563: dataIn1 = 32'd8681
; 
32'd178564: dataIn1 = 32'd8684
; 
32'd178565: dataIn1 = 32'd8685
; 
32'd178566: dataIn1 = 32'd8704
; 
32'd178567: dataIn1 = 32'd8707
; 
32'd178568: dataIn1 = 32'd5254
; 
32'd178569: dataIn1 = 32'd6532
; 
32'd178570: dataIn1 = 32'd8681
; 
32'd178571: dataIn1 = 32'd8684
; 
32'd178572: dataIn1 = 32'd8685
; 
32'd178573: dataIn1 = 32'd8697
; 
32'd178574: dataIn1 = 32'd8700
; 
32'd178575: dataIn1 = 32'd5255
; 
32'd178576: dataIn1 = 32'd6533
; 
32'd178577: dataIn1 = 32'd8682
; 
32'd178578: dataIn1 = 32'd8686
; 
32'd178579: dataIn1 = 32'd8687
; 
32'd178580: dataIn1 = 32'd8705
; 
32'd178581: dataIn1 = 32'd8708
; 
32'd178582: dataIn1 = 32'd5255
; 
32'd178583: dataIn1 = 32'd6531
; 
32'd178584: dataIn1 = 32'd8682
; 
32'd178585: dataIn1 = 32'd8686
; 
32'd178586: dataIn1 = 32'd8687
; 
32'd178587: dataIn1 = 32'd8691
; 
32'd178588: dataIn1 = 32'd8695
; 
32'd178589: dataIn1 = 32'd5256
; 
32'd178590: dataIn1 = 32'd6532
; 
32'd178591: dataIn1 = 32'd8683
; 
32'd178592: dataIn1 = 32'd8688
; 
32'd178593: dataIn1 = 32'd8689
; 
32'd178594: dataIn1 = 32'd8699
; 
32'd178595: dataIn1 = 32'd8703
; 
32'd178596: dataIn1 = 32'd5256
; 
32'd178597: dataIn1 = 32'd6531
; 
32'd178598: dataIn1 = 32'd8683
; 
32'd178599: dataIn1 = 32'd8688
; 
32'd178600: dataIn1 = 32'd8689
; 
32'd178601: dataIn1 = 32'd8692
; 
32'd178602: dataIn1 = 32'd8696
; 
32'd178603: dataIn1 = 32'd6534
; 
32'd178604: dataIn1 = 32'd6535
; 
32'd178605: dataIn1 = 32'd8690
; 
32'd178606: dataIn1 = 32'd8691
; 
32'd178607: dataIn1 = 32'd8692
; 
32'd178608: dataIn1 = 32'd8693
; 
32'd178609: dataIn1 = 32'd8694
; 
32'd178610: dataIn1 = 32'd6531
; 
32'd178611: dataIn1 = 32'd6535
; 
32'd178612: dataIn1 = 32'd8687
; 
32'd178613: dataIn1 = 32'd8690
; 
32'd178614: dataIn1 = 32'd8691
; 
32'd178615: dataIn1 = 32'd8692
; 
32'd178616: dataIn1 = 32'd8695
; 
32'd178617: dataIn1 = 32'd6531
; 
32'd178618: dataIn1 = 32'd6534
; 
32'd178619: dataIn1 = 32'd8689
; 
32'd178620: dataIn1 = 32'd8690
; 
32'd178621: dataIn1 = 32'd8691
; 
32'd178622: dataIn1 = 32'd8692
; 
32'd178623: dataIn1 = 32'd8696
; 
32'd178624: dataIn1 = 32'd2729
; 
32'd178625: dataIn1 = 32'd6535
; 
32'd178626: dataIn1 = 32'd8660
; 
32'd178627: dataIn1 = 32'd8690
; 
32'd178628: dataIn1 = 32'd8693
; 
32'd178629: dataIn1 = 32'd8694
; 
32'd178630: dataIn1 = 32'd8746
; 
32'd178631: dataIn1 = 32'd2729
; 
32'd178632: dataIn1 = 32'd6534
; 
32'd178633: dataIn1 = 32'd8677
; 
32'd178634: dataIn1 = 32'd8690
; 
32'd178635: dataIn1 = 32'd8693
; 
32'd178636: dataIn1 = 32'd8694
; 
32'd178637: dataIn1 = 32'd8768
; 
32'd178638: dataIn1 = 32'd5255
; 
32'd178639: dataIn1 = 32'd6535
; 
32'd178640: dataIn1 = 32'd8687
; 
32'd178641: dataIn1 = 32'd8691
; 
32'd178642: dataIn1 = 32'd8695
; 
32'd178643: dataIn1 = 32'd8743
; 
32'd178644: dataIn1 = 32'd8747
; 
32'd178645: dataIn1 = 32'd5256
; 
32'd178646: dataIn1 = 32'd6534
; 
32'd178647: dataIn1 = 32'd8689
; 
32'd178648: dataIn1 = 32'd8692
; 
32'd178649: dataIn1 = 32'd8696
; 
32'd178650: dataIn1 = 32'd8767
; 
32'd178651: dataIn1 = 32'd8770
; 
32'd178652: dataIn1 = 32'd6532
; 
32'd178653: dataIn1 = 32'd6537
; 
32'd178654: dataIn1 = 32'd8685
; 
32'd178655: dataIn1 = 32'd8697
; 
32'd178656: dataIn1 = 32'd8698
; 
32'd178657: dataIn1 = 32'd8699
; 
32'd178658: dataIn1 = 32'd8700
; 
32'd178659: dataIn1 = 32'd6536
; 
32'd178660: dataIn1 = 32'd6537
; 
32'd178661: dataIn1 = 32'd8697
; 
32'd178662: dataIn1 = 32'd8698
; 
32'd178663: dataIn1 = 32'd8699
; 
32'd178664: dataIn1 = 32'd8701
; 
32'd178665: dataIn1 = 32'd8702
; 
32'd178666: dataIn1 = 32'd6532
; 
32'd178667: dataIn1 = 32'd6536
; 
32'd178668: dataIn1 = 32'd8688
; 
32'd178669: dataIn1 = 32'd8697
; 
32'd178670: dataIn1 = 32'd8698
; 
32'd178671: dataIn1 = 32'd8699
; 
32'd178672: dataIn1 = 32'd8703
; 
32'd178673: dataIn1 = 32'd5254
; 
32'd178674: dataIn1 = 32'd6537
; 
32'd178675: dataIn1 = 32'd8685
; 
32'd178676: dataIn1 = 32'd8697
; 
32'd178677: dataIn1 = 32'd8700
; 
32'd178678: dataIn1 = 32'd8715
; 
32'd178679: dataIn1 = 32'd8727
; 
32'd178680: dataIn1 = 32'd2732
; 
32'd178681: dataIn1 = 32'd6537
; 
32'd178682: dataIn1 = 32'd8698
; 
32'd178683: dataIn1 = 32'd8701
; 
32'd178684: dataIn1 = 32'd8702
; 
32'd178685: dataIn1 = 32'd8728
; 
32'd178686: dataIn1 = 32'd8730
; 
32'd178687: dataIn1 = 32'd2732
; 
32'd178688: dataIn1 = 32'd6536
; 
32'd178689: dataIn1 = 32'd8698
; 
32'd178690: dataIn1 = 32'd8701
; 
32'd178691: dataIn1 = 32'd8702
; 
32'd178692: dataIn1 = 32'd8772
; 
32'd178693: dataIn1 = 32'd8775
; 
32'd178694: dataIn1 = 32'd5256
; 
32'd178695: dataIn1 = 32'd6536
; 
32'd178696: dataIn1 = 32'd8688
; 
32'd178697: dataIn1 = 32'd8699
; 
32'd178698: dataIn1 = 32'd8703
; 
32'd178699: dataIn1 = 32'd8766
; 
32'd178700: dataIn1 = 32'd8773
; 
32'd178701: dataIn1 = 32'd6533
; 
32'd178702: dataIn1 = 32'd6539
; 
32'd178703: dataIn1 = 32'd8684
; 
32'd178704: dataIn1 = 32'd8704
; 
32'd178705: dataIn1 = 32'd8705
; 
32'd178706: dataIn1 = 32'd8706
; 
32'd178707: dataIn1 = 32'd8707
; 
32'd178708: dataIn1 = 32'd6533
; 
32'd178709: dataIn1 = 32'd6538
; 
32'd178710: dataIn1 = 32'd8686
; 
32'd178711: dataIn1 = 32'd8704
; 
32'd178712: dataIn1 = 32'd8705
; 
32'd178713: dataIn1 = 32'd8706
; 
32'd178714: dataIn1 = 32'd8708
; 
32'd178715: dataIn1 = 32'd6538
; 
32'd178716: dataIn1 = 32'd6539
; 
32'd178717: dataIn1 = 32'd8704
; 
32'd178718: dataIn1 = 32'd8705
; 
32'd178719: dataIn1 = 32'd8706
; 
32'd178720: dataIn1 = 32'd8709
; 
32'd178721: dataIn1 = 32'd8710
; 
32'd178722: dataIn1 = 32'd5254
; 
32'd178723: dataIn1 = 32'd6539
; 
32'd178724: dataIn1 = 32'd8684
; 
32'd178725: dataIn1 = 32'd8704
; 
32'd178726: dataIn1 = 32'd8707
; 
32'd178727: dataIn1 = 32'd8714
; 
32'd178728: dataIn1 = 32'd8732
; 
32'd178729: dataIn1 = 32'd5255
; 
32'd178730: dataIn1 = 32'd6538
; 
32'd178731: dataIn1 = 32'd8686
; 
32'd178732: dataIn1 = 32'd8705
; 
32'd178733: dataIn1 = 32'd8708
; 
32'd178734: dataIn1 = 32'd8742
; 
32'd178735: dataIn1 = 32'd8755
; 
32'd178736: dataIn1 = 32'd1117
; 
32'd178737: dataIn1 = 32'd6539
; 
32'd178738: dataIn1 = 32'd8706
; 
32'd178739: dataIn1 = 32'd8709
; 
32'd178740: dataIn1 = 32'd8710
; 
32'd178741: dataIn1 = 32'd8734
; 
32'd178742: dataIn1 = 32'd8736
; 
32'd178743: dataIn1 = 32'd1117
; 
32'd178744: dataIn1 = 32'd6538
; 
32'd178745: dataIn1 = 32'd8706
; 
32'd178746: dataIn1 = 32'd8709
; 
32'd178747: dataIn1 = 32'd8710
; 
32'd178748: dataIn1 = 32'd8756
; 
32'd178749: dataIn1 = 32'd8758
; 
32'd178750: dataIn1 = 32'd6541
; 
32'd178751: dataIn1 = 32'd6542
; 
32'd178752: dataIn1 = 32'd8711
; 
32'd178753: dataIn1 = 32'd8712
; 
32'd178754: dataIn1 = 32'd8713
; 
32'd178755: dataIn1 = 32'd8714
; 
32'd178756: dataIn1 = 32'd8715
; 
32'd178757: dataIn1 = 32'd6540
; 
32'd178758: dataIn1 = 32'd6542
; 
32'd178759: dataIn1 = 32'd8711
; 
32'd178760: dataIn1 = 32'd8712
; 
32'd178761: dataIn1 = 32'd8713
; 
32'd178762: dataIn1 = 32'd8716
; 
32'd178763: dataIn1 = 32'd8717
; 
32'd178764: dataIn1 = 32'd6540
; 
32'd178765: dataIn1 = 32'd6541
; 
32'd178766: dataIn1 = 32'd8711
; 
32'd178767: dataIn1 = 32'd8712
; 
32'd178768: dataIn1 = 32'd8713
; 
32'd178769: dataIn1 = 32'd8718
; 
32'd178770: dataIn1 = 32'd8719
; 
32'd178771: dataIn1 = 32'd5254
; 
32'd178772: dataIn1 = 32'd6542
; 
32'd178773: dataIn1 = 32'd8707
; 
32'd178774: dataIn1 = 32'd8711
; 
32'd178775: dataIn1 = 32'd8714
; 
32'd178776: dataIn1 = 32'd8715
; 
32'd178777: dataIn1 = 32'd8732
; 
32'd178778: dataIn1 = 32'd5254
; 
32'd178779: dataIn1 = 32'd6541
; 
32'd178780: dataIn1 = 32'd8700
; 
32'd178781: dataIn1 = 32'd8711
; 
32'd178782: dataIn1 = 32'd8714
; 
32'd178783: dataIn1 = 32'd8715
; 
32'd178784: dataIn1 = 32'd8727
; 
32'd178785: dataIn1 = 32'd2686
; 
32'd178786: dataIn1 = 32'd6542
; 
32'd178787: dataIn1 = 32'd8712
; 
32'd178788: dataIn1 = 32'd8716
; 
32'd178789: dataIn1 = 32'd8717
; 
32'd178790: dataIn1 = 32'd8733
; 
32'd178791: dataIn1 = 32'd8735
; 
32'd178792: dataIn1 = 32'd2686
; 
32'd178793: dataIn1 = 32'd6540
; 
32'd178794: dataIn1 = 32'd8712
; 
32'd178795: dataIn1 = 32'd8716
; 
32'd178796: dataIn1 = 32'd8717
; 
32'd178797: dataIn1 = 32'd8721
; 
32'd178798: dataIn1 = 32'd8725
; 
32'd178799: dataIn1 = 32'd5257
; 
32'd178800: dataIn1 = 32'd6541
; 
32'd178801: dataIn1 = 32'd8713
; 
32'd178802: dataIn1 = 32'd8718
; 
32'd178803: dataIn1 = 32'd8719
; 
32'd178804: dataIn1 = 32'd8729
; 
32'd178805: dataIn1 = 32'd8731
; 
32'd178806: dataIn1 = 32'd5257
; 
32'd178807: dataIn1 = 32'd6540
; 
32'd178808: dataIn1 = 32'd8713
; 
32'd178809: dataIn1 = 32'd8718
; 
32'd178810: dataIn1 = 32'd8719
; 
32'd178811: dataIn1 = 32'd8722
; 
32'd178812: dataIn1 = 32'd8726
; 
32'd178813: dataIn1 = 32'd5091
; 
32'd178814: dataIn1 = 32'd6543
; 
32'd178815: dataIn1 = 32'd8720
; 
32'd178816: dataIn1 = 32'd8721
; 
32'd178817: dataIn1 = 32'd8722
; 
32'd178818: dataIn1 = 32'd8723
; 
32'd178819: dataIn1 = 32'd8724
; 
32'd178820: dataIn1 = 32'd5091
; 
32'd178821: dataIn1 = 32'd6540
; 
32'd178822: dataIn1 = 32'd8717
; 
32'd178823: dataIn1 = 32'd8720
; 
32'd178824: dataIn1 = 32'd8721
; 
32'd178825: dataIn1 = 32'd8722
; 
32'd178826: dataIn1 = 32'd8725
; 
32'd178827: dataIn1 = 32'd6540
; 
32'd178828: dataIn1 = 32'd6543
; 
32'd178829: dataIn1 = 32'd8719
; 
32'd178830: dataIn1 = 32'd8720
; 
32'd178831: dataIn1 = 32'd8721
; 
32'd178832: dataIn1 = 32'd8722
; 
32'd178833: dataIn1 = 32'd8726
; 
32'd178834: dataIn1 = 32'd11
; 
32'd178835: dataIn1 = 32'd4771
; 
32'd178836: dataIn1 = 32'd5091
; 
32'd178837: dataIn1 = 32'd8720
; 
32'd178838: dataIn1 = 32'd8723
; 
32'd178839: dataIn1 = 32'd8724
; 
32'd178840: dataIn1 = 32'd11
; 
32'd178841: dataIn1 = 32'd6543
; 
32'd178842: dataIn1 = 32'd8616
; 
32'd178843: dataIn1 = 32'd8720
; 
32'd178844: dataIn1 = 32'd8723
; 
32'd178845: dataIn1 = 32'd8724
; 
32'd178846: dataIn1 = 32'd9213
; 
32'd178847: dataIn1 = 32'd2686
; 
32'd178848: dataIn1 = 32'd5089
; 
32'd178849: dataIn1 = 32'd5091
; 
32'd178850: dataIn1 = 32'd8717
; 
32'd178851: dataIn1 = 32'd8721
; 
32'd178852: dataIn1 = 32'd8725
; 
32'd178853: dataIn1 = 32'd5257
; 
32'd178854: dataIn1 = 32'd6543
; 
32'd178855: dataIn1 = 32'd8719
; 
32'd178856: dataIn1 = 32'd8722
; 
32'd178857: dataIn1 = 32'd8726
; 
32'd178858: dataIn1 = 32'd9210
; 
32'd178859: dataIn1 = 32'd9214
; 
32'd178860: dataIn1 = 32'd6537
; 
32'd178861: dataIn1 = 32'd6541
; 
32'd178862: dataIn1 = 32'd8700
; 
32'd178863: dataIn1 = 32'd8715
; 
32'd178864: dataIn1 = 32'd8727
; 
32'd178865: dataIn1 = 32'd8728
; 
32'd178866: dataIn1 = 32'd8729
; 
32'd178867: dataIn1 = 32'd6537
; 
32'd178868: dataIn1 = 32'd6544
; 
32'd178869: dataIn1 = 32'd8701
; 
32'd178870: dataIn1 = 32'd8727
; 
32'd178871: dataIn1 = 32'd8728
; 
32'd178872: dataIn1 = 32'd8729
; 
32'd178873: dataIn1 = 32'd8730
; 
32'd178874: dataIn1 = 32'd6541
; 
32'd178875: dataIn1 = 32'd6544
; 
32'd178876: dataIn1 = 32'd8718
; 
32'd178877: dataIn1 = 32'd8727
; 
32'd178878: dataIn1 = 32'd8728
; 
32'd178879: dataIn1 = 32'd8729
; 
32'd178880: dataIn1 = 32'd8731
; 
32'd178881: dataIn1 = 32'd2732
; 
32'd178882: dataIn1 = 32'd6544
; 
32'd178883: dataIn1 = 32'd8701
; 
32'd178884: dataIn1 = 32'd8728
; 
32'd178885: dataIn1 = 32'd8730
; 
32'd178886: dataIn1 = 32'd9202
; 
32'd178887: dataIn1 = 32'd9221
; 
32'd178888: dataIn1 = 32'd5257
; 
32'd178889: dataIn1 = 32'd6544
; 
32'd178890: dataIn1 = 32'd8718
; 
32'd178891: dataIn1 = 32'd8729
; 
32'd178892: dataIn1 = 32'd8731
; 
32'd178893: dataIn1 = 32'd9209
; 
32'd178894: dataIn1 = 32'd9220
; 
32'd178895: dataIn1 = 32'd6539
; 
32'd178896: dataIn1 = 32'd6542
; 
32'd178897: dataIn1 = 32'd8707
; 
32'd178898: dataIn1 = 32'd8714
; 
32'd178899: dataIn1 = 32'd8732
; 
32'd178900: dataIn1 = 32'd8733
; 
32'd178901: dataIn1 = 32'd8734
; 
32'd178902: dataIn1 = 32'd5092
; 
32'd178903: dataIn1 = 32'd6542
; 
32'd178904: dataIn1 = 32'd8716
; 
32'd178905: dataIn1 = 32'd8732
; 
32'd178906: dataIn1 = 32'd8733
; 
32'd178907: dataIn1 = 32'd8734
; 
32'd178908: dataIn1 = 32'd8735
; 
32'd178909: dataIn1 = 32'd5092
; 
32'd178910: dataIn1 = 32'd6539
; 
32'd178911: dataIn1 = 32'd8709
; 
32'd178912: dataIn1 = 32'd8732
; 
32'd178913: dataIn1 = 32'd8733
; 
32'd178914: dataIn1 = 32'd8734
; 
32'd178915: dataIn1 = 32'd8736
; 
32'd178916: dataIn1 = 32'd2686
; 
32'd178917: dataIn1 = 32'd5090
; 
32'd178918: dataIn1 = 32'd5092
; 
32'd178919: dataIn1 = 32'd8716
; 
32'd178920: dataIn1 = 32'd8733
; 
32'd178921: dataIn1 = 32'd8735
; 
32'd178922: dataIn1 = 32'd1117
; 
32'd178923: dataIn1 = 32'd5081
; 
32'd178924: dataIn1 = 32'd5092
; 
32'd178925: dataIn1 = 32'd8709
; 
32'd178926: dataIn1 = 32'd8734
; 
32'd178927: dataIn1 = 32'd8736
; 
32'd178928: dataIn1 = 32'd6546
; 
32'd178929: dataIn1 = 32'd6547
; 
32'd178930: dataIn1 = 32'd8737
; 
32'd178931: dataIn1 = 32'd8738
; 
32'd178932: dataIn1 = 32'd8739
; 
32'd178933: dataIn1 = 32'd8740
; 
32'd178934: dataIn1 = 32'd8741
; 
32'd178935: dataIn1 = 32'd6545
; 
32'd178936: dataIn1 = 32'd6547
; 
32'd178937: dataIn1 = 32'd8737
; 
32'd178938: dataIn1 = 32'd8738
; 
32'd178939: dataIn1 = 32'd8739
; 
32'd178940: dataIn1 = 32'd8742
; 
32'd178941: dataIn1 = 32'd8743
; 
32'd178942: dataIn1 = 32'd6545
; 
32'd178943: dataIn1 = 32'd6546
; 
32'd178944: dataIn1 = 32'd8737
; 
32'd178945: dataIn1 = 32'd8738
; 
32'd178946: dataIn1 = 32'd8739
; 
32'd178947: dataIn1 = 32'd8744
; 
32'd178948: dataIn1 = 32'd8745
; 
32'd178949: dataIn1 = 32'd2685
; 
32'd178950: dataIn1 = 32'd6547
; 
32'd178951: dataIn1 = 32'd8737
; 
32'd178952: dataIn1 = 32'd8740
; 
32'd178953: dataIn1 = 32'd8741
; 
32'd178954: dataIn1 = 32'd8754
; 
32'd178955: dataIn1 = 32'd8757
; 
32'd178956: dataIn1 = 32'd2685
; 
32'd178957: dataIn1 = 32'd6546
; 
32'd178958: dataIn1 = 32'd8737
; 
32'd178959: dataIn1 = 32'd8740
; 
32'd178960: dataIn1 = 32'd8741
; 
32'd178961: dataIn1 = 32'd8749
; 
32'd178962: dataIn1 = 32'd8752
; 
32'd178963: dataIn1 = 32'd5255
; 
32'd178964: dataIn1 = 32'd6547
; 
32'd178965: dataIn1 = 32'd8708
; 
32'd178966: dataIn1 = 32'd8738
; 
32'd178967: dataIn1 = 32'd8742
; 
32'd178968: dataIn1 = 32'd8743
; 
32'd178969: dataIn1 = 32'd8755
; 
32'd178970: dataIn1 = 32'd5255
; 
32'd178971: dataIn1 = 32'd6545
; 
32'd178972: dataIn1 = 32'd8695
; 
32'd178973: dataIn1 = 32'd8738
; 
32'd178974: dataIn1 = 32'd8742
; 
32'd178975: dataIn1 = 32'd8743
; 
32'd178976: dataIn1 = 32'd8747
; 
32'd178977: dataIn1 = 32'd5251
; 
32'd178978: dataIn1 = 32'd6546
; 
32'd178979: dataIn1 = 32'd8668
; 
32'd178980: dataIn1 = 32'd8739
; 
32'd178981: dataIn1 = 32'd8744
; 
32'd178982: dataIn1 = 32'd8745
; 
32'd178983: dataIn1 = 32'd8751
; 
32'd178984: dataIn1 = 32'd5251
; 
32'd178985: dataIn1 = 32'd6545
; 
32'd178986: dataIn1 = 32'd8661
; 
32'd178987: dataIn1 = 32'd8739
; 
32'd178988: dataIn1 = 32'd8744
; 
32'd178989: dataIn1 = 32'd8745
; 
32'd178990: dataIn1 = 32'd8748
; 
32'd178991: dataIn1 = 32'd6525
; 
32'd178992: dataIn1 = 32'd6535
; 
32'd178993: dataIn1 = 32'd8660
; 
32'd178994: dataIn1 = 32'd8693
; 
32'd178995: dataIn1 = 32'd8746
; 
32'd178996: dataIn1 = 32'd8747
; 
32'd178997: dataIn1 = 32'd8748
; 
32'd178998: dataIn1 = 32'd6535
; 
32'd178999: dataIn1 = 32'd6545
; 
32'd179000: dataIn1 = 32'd8695
; 
32'd179001: dataIn1 = 32'd8743
; 
32'd179002: dataIn1 = 32'd8746
; 
32'd179003: dataIn1 = 32'd8747
; 
32'd179004: dataIn1 = 32'd8748
; 
32'd179005: dataIn1 = 32'd6525
; 
32'd179006: dataIn1 = 32'd6545
; 
32'd179007: dataIn1 = 32'd8661
; 
32'd179008: dataIn1 = 32'd8745
; 
32'd179009: dataIn1 = 32'd8746
; 
32'd179010: dataIn1 = 32'd8747
; 
32'd179011: dataIn1 = 32'd8748
; 
32'd179012: dataIn1 = 32'd5086
; 
32'd179013: dataIn1 = 32'd6546
; 
32'd179014: dataIn1 = 32'd8741
; 
32'd179015: dataIn1 = 32'd8749
; 
32'd179016: dataIn1 = 32'd8750
; 
32'd179017: dataIn1 = 32'd8751
; 
32'd179018: dataIn1 = 32'd8752
; 
32'd179019: dataIn1 = 32'd5086
; 
32'd179020: dataIn1 = 32'd6526
; 
32'd179021: dataIn1 = 32'd8667
; 
32'd179022: dataIn1 = 32'd8749
; 
32'd179023: dataIn1 = 32'd8750
; 
32'd179024: dataIn1 = 32'd8751
; 
32'd179025: dataIn1 = 32'd8753
; 
32'd179026: dataIn1 = 32'd6526
; 
32'd179027: dataIn1 = 32'd6546
; 
32'd179028: dataIn1 = 32'd8668
; 
32'd179029: dataIn1 = 32'd8744
; 
32'd179030: dataIn1 = 32'd8749
; 
32'd179031: dataIn1 = 32'd8750
; 
32'd179032: dataIn1 = 32'd8751
; 
32'd179033: dataIn1 = 32'd2685
; 
32'd179034: dataIn1 = 32'd5083
; 
32'd179035: dataIn1 = 32'd5086
; 
32'd179036: dataIn1 = 32'd8741
; 
32'd179037: dataIn1 = 32'd8749
; 
32'd179038: dataIn1 = 32'd8752
; 
32'd179039: dataIn1 = 32'd148
; 
32'd179040: dataIn1 = 32'd4777
; 
32'd179041: dataIn1 = 32'd5086
; 
32'd179042: dataIn1 = 32'd8667
; 
32'd179043: dataIn1 = 32'd8750
; 
32'd179044: dataIn1 = 32'd8753
; 
32'd179045: dataIn1 = 32'd5087
; 
32'd179046: dataIn1 = 32'd6547
; 
32'd179047: dataIn1 = 32'd8740
; 
32'd179048: dataIn1 = 32'd8754
; 
32'd179049: dataIn1 = 32'd8755
; 
32'd179050: dataIn1 = 32'd8756
; 
32'd179051: dataIn1 = 32'd8757
; 
32'd179052: dataIn1 = 32'd6538
; 
32'd179053: dataIn1 = 32'd6547
; 
32'd179054: dataIn1 = 32'd8708
; 
32'd179055: dataIn1 = 32'd8742
; 
32'd179056: dataIn1 = 32'd8754
; 
32'd179057: dataIn1 = 32'd8755
; 
32'd179058: dataIn1 = 32'd8756
; 
32'd179059: dataIn1 = 32'd5087
; 
32'd179060: dataIn1 = 32'd6538
; 
32'd179061: dataIn1 = 32'd8710
; 
32'd179062: dataIn1 = 32'd8754
; 
32'd179063: dataIn1 = 32'd8755
; 
32'd179064: dataIn1 = 32'd8756
; 
32'd179065: dataIn1 = 32'd8758
; 
32'd179066: dataIn1 = 32'd2685
; 
32'd179067: dataIn1 = 32'd5085
; 
32'd179068: dataIn1 = 32'd5087
; 
32'd179069: dataIn1 = 32'd8740
; 
32'd179070: dataIn1 = 32'd8754
; 
32'd179071: dataIn1 = 32'd8757
; 
32'd179072: dataIn1 = 32'd1117
; 
32'd179073: dataIn1 = 32'd5082
; 
32'd179074: dataIn1 = 32'd5087
; 
32'd179075: dataIn1 = 32'd8710
; 
32'd179076: dataIn1 = 32'd8756
; 
32'd179077: dataIn1 = 32'd8758
; 
32'd179078: dataIn1 = 32'd6549
; 
32'd179079: dataIn1 = 32'd6550
; 
32'd179080: dataIn1 = 32'd8759
; 
32'd179081: dataIn1 = 32'd8760
; 
32'd179082: dataIn1 = 32'd8761
; 
32'd179083: dataIn1 = 32'd8762
; 
32'd179084: dataIn1 = 32'd8763
; 
32'd179085: dataIn1 = 32'd6548
; 
32'd179086: dataIn1 = 32'd6550
; 
32'd179087: dataIn1 = 32'd8759
; 
32'd179088: dataIn1 = 32'd8760
; 
32'd179089: dataIn1 = 32'd8761
; 
32'd179090: dataIn1 = 32'd8764
; 
32'd179091: dataIn1 = 32'd8765
; 
32'd179092: dataIn1 = 32'd6548
; 
32'd179093: dataIn1 = 32'd6549
; 
32'd179094: dataIn1 = 32'd8759
; 
32'd179095: dataIn1 = 32'd8760
; 
32'd179096: dataIn1 = 32'd8761
; 
32'd179097: dataIn1 = 32'd8766
; 
32'd179098: dataIn1 = 32'd8767
; 
32'd179099: dataIn1 = 32'd5258
; 
32'd179100: dataIn1 = 32'd6550
; 
32'd179101: dataIn1 = 32'd6783
; 
32'd179102: dataIn1 = 32'd8759
; 
32'd179103: dataIn1 = 32'd8762
; 
32'd179104: dataIn1 = 32'd8763
; 
32'd179105: dataIn1 = 32'd5258
; 
32'd179106: dataIn1 = 32'd6549
; 
32'd179107: dataIn1 = 32'd8759
; 
32'd179108: dataIn1 = 32'd8762
; 
32'd179109: dataIn1 = 32'd8763
; 
32'd179110: dataIn1 = 32'd8771
; 
32'd179111: dataIn1 = 32'd8774
; 
32'd179112: dataIn1 = 32'd5253
; 
32'd179113: dataIn1 = 32'd6550
; 
32'd179114: dataIn1 = 32'd6782
; 
32'd179115: dataIn1 = 32'd8760
; 
32'd179116: dataIn1 = 32'd8764
; 
32'd179117: dataIn1 = 32'd8765
; 
32'd179118: dataIn1 = 32'd5253
; 
32'd179119: dataIn1 = 32'd6548
; 
32'd179120: dataIn1 = 32'd8678
; 
32'd179121: dataIn1 = 32'd8760
; 
32'd179122: dataIn1 = 32'd8764
; 
32'd179123: dataIn1 = 32'd8765
; 
32'd179124: dataIn1 = 32'd8769
; 
32'd179125: dataIn1 = 32'd5256
; 
32'd179126: dataIn1 = 32'd6549
; 
32'd179127: dataIn1 = 32'd8703
; 
32'd179128: dataIn1 = 32'd8761
; 
32'd179129: dataIn1 = 32'd8766
; 
32'd179130: dataIn1 = 32'd8767
; 
32'd179131: dataIn1 = 32'd8773
; 
32'd179132: dataIn1 = 32'd5256
; 
32'd179133: dataIn1 = 32'd6548
; 
32'd179134: dataIn1 = 32'd8696
; 
32'd179135: dataIn1 = 32'd8761
; 
32'd179136: dataIn1 = 32'd8766
; 
32'd179137: dataIn1 = 32'd8767
; 
32'd179138: dataIn1 = 32'd8770
; 
32'd179139: dataIn1 = 32'd6530
; 
32'd179140: dataIn1 = 32'd6534
; 
32'd179141: dataIn1 = 32'd8677
; 
32'd179142: dataIn1 = 32'd8694
; 
32'd179143: dataIn1 = 32'd8768
; 
32'd179144: dataIn1 = 32'd8769
; 
32'd179145: dataIn1 = 32'd8770
; 
32'd179146: dataIn1 = 32'd6530
; 
32'd179147: dataIn1 = 32'd6548
; 
32'd179148: dataIn1 = 32'd8678
; 
32'd179149: dataIn1 = 32'd8765
; 
32'd179150: dataIn1 = 32'd8768
; 
32'd179151: dataIn1 = 32'd8769
; 
32'd179152: dataIn1 = 32'd8770
; 
32'd179153: dataIn1 = 32'd6534
; 
32'd179154: dataIn1 = 32'd6548
; 
32'd179155: dataIn1 = 32'd8696
; 
32'd179156: dataIn1 = 32'd8767
; 
32'd179157: dataIn1 = 32'd8768
; 
32'd179158: dataIn1 = 32'd8769
; 
32'd179159: dataIn1 = 32'd8770
; 
32'd179160: dataIn1 = 32'd6549
; 
32'd179161: dataIn1 = 32'd6551
; 
32'd179162: dataIn1 = 32'd8763
; 
32'd179163: dataIn1 = 32'd8771
; 
32'd179164: dataIn1 = 32'd8772
; 
32'd179165: dataIn1 = 32'd8773
; 
32'd179166: dataIn1 = 32'd8774
; 
32'd179167: dataIn1 = 32'd6536
; 
32'd179168: dataIn1 = 32'd6551
; 
32'd179169: dataIn1 = 32'd8702
; 
32'd179170: dataIn1 = 32'd8771
; 
32'd179171: dataIn1 = 32'd8772
; 
32'd179172: dataIn1 = 32'd8773
; 
32'd179173: dataIn1 = 32'd8775
; 
32'd179174: dataIn1 = 32'd6536
; 
32'd179175: dataIn1 = 32'd6549
; 
32'd179176: dataIn1 = 32'd8703
; 
32'd179177: dataIn1 = 32'd8766
; 
32'd179178: dataIn1 = 32'd8771
; 
32'd179179: dataIn1 = 32'd8772
; 
32'd179180: dataIn1 = 32'd8773
; 
32'd179181: dataIn1 = 32'd5258
; 
32'd179182: dataIn1 = 32'd6551
; 
32'd179183: dataIn1 = 32'd8763
; 
32'd179184: dataIn1 = 32'd8771
; 
32'd179185: dataIn1 = 32'd8774
; 
32'd179186: dataIn1 = 32'd9222
; 
32'd179187: dataIn1 = 32'd9225
; 
32'd179188: dataIn1 = 32'd2732
; 
32'd179189: dataIn1 = 32'd6551
; 
32'd179190: dataIn1 = 32'd8702
; 
32'd179191: dataIn1 = 32'd8772
; 
32'd179192: dataIn1 = 32'd8775
; 
32'd179193: dataIn1 = 32'd9203
; 
32'd179194: dataIn1 = 32'd9224
; 
32'd179195: dataIn1 = 32'd6553
; 
32'd179196: dataIn1 = 32'd6554
; 
32'd179197: dataIn1 = 32'd8776
; 
32'd179198: dataIn1 = 32'd8777
; 
32'd179199: dataIn1 = 32'd8778
; 
32'd179200: dataIn1 = 32'd8779
; 
32'd179201: dataIn1 = 32'd8780
; 
32'd179202: dataIn1 = 32'd6552
; 
32'd179203: dataIn1 = 32'd6554
; 
32'd179204: dataIn1 = 32'd8776
; 
32'd179205: dataIn1 = 32'd8777
; 
32'd179206: dataIn1 = 32'd8778
; 
32'd179207: dataIn1 = 32'd8781
; 
32'd179208: dataIn1 = 32'd8782
; 
32'd179209: dataIn1 = 32'd6552
; 
32'd179210: dataIn1 = 32'd6553
; 
32'd179211: dataIn1 = 32'd8776
; 
32'd179212: dataIn1 = 32'd8777
; 
32'd179213: dataIn1 = 32'd8778
; 
32'd179214: dataIn1 = 32'd8783
; 
32'd179215: dataIn1 = 32'd8784
; 
32'd179216: dataIn1 = 32'd5259
; 
32'd179217: dataIn1 = 32'd6554
; 
32'd179218: dataIn1 = 32'd8776
; 
32'd179219: dataIn1 = 32'd8779
; 
32'd179220: dataIn1 = 32'd8780
; 
32'd179221: dataIn1 = 32'd8799
; 
32'd179222: dataIn1 = 32'd8802
; 
32'd179223: dataIn1 = 32'd5259
; 
32'd179224: dataIn1 = 32'd6553
; 
32'd179225: dataIn1 = 32'd8776
; 
32'd179226: dataIn1 = 32'd8779
; 
32'd179227: dataIn1 = 32'd8780
; 
32'd179228: dataIn1 = 32'd8792
; 
32'd179229: dataIn1 = 32'd8795
; 
32'd179230: dataIn1 = 32'd5260
; 
32'd179231: dataIn1 = 32'd6554
; 
32'd179232: dataIn1 = 32'd8777
; 
32'd179233: dataIn1 = 32'd8781
; 
32'd179234: dataIn1 = 32'd8782
; 
32'd179235: dataIn1 = 32'd8800
; 
32'd179236: dataIn1 = 32'd8803
; 
32'd179237: dataIn1 = 32'd5260
; 
32'd179238: dataIn1 = 32'd6552
; 
32'd179239: dataIn1 = 32'd8777
; 
32'd179240: dataIn1 = 32'd8781
; 
32'd179241: dataIn1 = 32'd8782
; 
32'd179242: dataIn1 = 32'd8786
; 
32'd179243: dataIn1 = 32'd8790
; 
32'd179244: dataIn1 = 32'd5261
; 
32'd179245: dataIn1 = 32'd6553
; 
32'd179246: dataIn1 = 32'd8778
; 
32'd179247: dataIn1 = 32'd8783
; 
32'd179248: dataIn1 = 32'd8784
; 
32'd179249: dataIn1 = 32'd8794
; 
32'd179250: dataIn1 = 32'd8798
; 
32'd179251: dataIn1 = 32'd5261
; 
32'd179252: dataIn1 = 32'd6552
; 
32'd179253: dataIn1 = 32'd8778
; 
32'd179254: dataIn1 = 32'd8783
; 
32'd179255: dataIn1 = 32'd8784
; 
32'd179256: dataIn1 = 32'd8787
; 
32'd179257: dataIn1 = 32'd8791
; 
32'd179258: dataIn1 = 32'd6555
; 
32'd179259: dataIn1 = 32'd6556
; 
32'd179260: dataIn1 = 32'd8785
; 
32'd179261: dataIn1 = 32'd8786
; 
32'd179262: dataIn1 = 32'd8787
; 
32'd179263: dataIn1 = 32'd8788
; 
32'd179264: dataIn1 = 32'd8789
; 
32'd179265: dataIn1 = 32'd6552
; 
32'd179266: dataIn1 = 32'd6556
; 
32'd179267: dataIn1 = 32'd8782
; 
32'd179268: dataIn1 = 32'd8785
; 
32'd179269: dataIn1 = 32'd8786
; 
32'd179270: dataIn1 = 32'd8787
; 
32'd179271: dataIn1 = 32'd8790
; 
32'd179272: dataIn1 = 32'd6552
; 
32'd179273: dataIn1 = 32'd6555
; 
32'd179274: dataIn1 = 32'd8784
; 
32'd179275: dataIn1 = 32'd8785
; 
32'd179276: dataIn1 = 32'd8786
; 
32'd179277: dataIn1 = 32'd8787
; 
32'd179278: dataIn1 = 32'd8791
; 
32'd179279: dataIn1 = 32'd1118
; 
32'd179280: dataIn1 = 32'd6556
; 
32'd179281: dataIn1 = 32'd8785
; 
32'd179282: dataIn1 = 32'd8788
; 
32'd179283: dataIn1 = 32'd8789
; 
32'd179284: dataIn1 = 32'd8831
; 
32'd179285: dataIn1 = 32'd8834
; 
32'd179286: dataIn1 = 32'd1118
; 
32'd179287: dataIn1 = 32'd6555
; 
32'd179288: dataIn1 = 32'd8785
; 
32'd179289: dataIn1 = 32'd8788
; 
32'd179290: dataIn1 = 32'd8789
; 
32'd179291: dataIn1 = 32'd8853
; 
32'd179292: dataIn1 = 32'd8856
; 
32'd179293: dataIn1 = 32'd5260
; 
32'd179294: dataIn1 = 32'd6556
; 
32'd179295: dataIn1 = 32'd8782
; 
32'd179296: dataIn1 = 32'd8786
; 
32'd179297: dataIn1 = 32'd8790
; 
32'd179298: dataIn1 = 32'd8828
; 
32'd179299: dataIn1 = 32'd8832
; 
32'd179300: dataIn1 = 32'd5261
; 
32'd179301: dataIn1 = 32'd6555
; 
32'd179302: dataIn1 = 32'd8784
; 
32'd179303: dataIn1 = 32'd8787
; 
32'd179304: dataIn1 = 32'd8791
; 
32'd179305: dataIn1 = 32'd8852
; 
32'd179306: dataIn1 = 32'd8855
; 
32'd179307: dataIn1 = 32'd6553
; 
32'd179308: dataIn1 = 32'd6558
; 
32'd179309: dataIn1 = 32'd8780
; 
32'd179310: dataIn1 = 32'd8792
; 
32'd179311: dataIn1 = 32'd8793
; 
32'd179312: dataIn1 = 32'd8794
; 
32'd179313: dataIn1 = 32'd8795
; 
32'd179314: dataIn1 = 32'd6557
; 
32'd179315: dataIn1 = 32'd6558
; 
32'd179316: dataIn1 = 32'd8792
; 
32'd179317: dataIn1 = 32'd8793
; 
32'd179318: dataIn1 = 32'd8794
; 
32'd179319: dataIn1 = 32'd8796
; 
32'd179320: dataIn1 = 32'd8797
; 
32'd179321: dataIn1 = 32'd6553
; 
32'd179322: dataIn1 = 32'd6557
; 
32'd179323: dataIn1 = 32'd8783
; 
32'd179324: dataIn1 = 32'd8792
; 
32'd179325: dataIn1 = 32'd8793
; 
32'd179326: dataIn1 = 32'd8794
; 
32'd179327: dataIn1 = 32'd8798
; 
32'd179328: dataIn1 = 32'd5259
; 
32'd179329: dataIn1 = 32'd6558
; 
32'd179330: dataIn1 = 32'd8780
; 
32'd179331: dataIn1 = 32'd8792
; 
32'd179332: dataIn1 = 32'd8795
; 
32'd179333: dataIn1 = 32'd8810
; 
32'd179334: dataIn1 = 32'd8815
; 
32'd179335: dataIn1 = 32'd2733
; 
32'd179336: dataIn1 = 32'd6558
; 
32'd179337: dataIn1 = 32'd8793
; 
32'd179338: dataIn1 = 32'd8796
; 
32'd179339: dataIn1 = 32'd8797
; 
32'd179340: dataIn1 = 32'd8816
; 
32'd179341: dataIn1 = 32'd9276
; 
32'd179342: dataIn1 = 32'd2733
; 
32'd179343: dataIn1 = 32'd6557
; 
32'd179344: dataIn1 = 32'd8793
; 
32'd179345: dataIn1 = 32'd8796
; 
32'd179346: dataIn1 = 32'd8797
; 
32'd179347: dataIn1 = 32'd8859
; 
32'd179348: dataIn1 = 32'd8862
; 
32'd179349: dataIn1 = 32'd5261
; 
32'd179350: dataIn1 = 32'd6557
; 
32'd179351: dataIn1 = 32'd8783
; 
32'd179352: dataIn1 = 32'd8794
; 
32'd179353: dataIn1 = 32'd8798
; 
32'd179354: dataIn1 = 32'd8851
; 
32'd179355: dataIn1 = 32'd8860
; 
32'd179356: dataIn1 = 32'd6554
; 
32'd179357: dataIn1 = 32'd6560
; 
32'd179358: dataIn1 = 32'd8779
; 
32'd179359: dataIn1 = 32'd8799
; 
32'd179360: dataIn1 = 32'd8800
; 
32'd179361: dataIn1 = 32'd8801
; 
32'd179362: dataIn1 = 32'd8802
; 
32'd179363: dataIn1 = 32'd6554
; 
32'd179364: dataIn1 = 32'd6559
; 
32'd179365: dataIn1 = 32'd8781
; 
32'd179366: dataIn1 = 32'd8799
; 
32'd179367: dataIn1 = 32'd8800
; 
32'd179368: dataIn1 = 32'd8801
; 
32'd179369: dataIn1 = 32'd8803
; 
32'd179370: dataIn1 = 32'd6559
; 
32'd179371: dataIn1 = 32'd6560
; 
32'd179372: dataIn1 = 32'd8799
; 
32'd179373: dataIn1 = 32'd8800
; 
32'd179374: dataIn1 = 32'd8801
; 
32'd179375: dataIn1 = 32'd8804
; 
32'd179376: dataIn1 = 32'd8805
; 
32'd179377: dataIn1 = 32'd5259
; 
32'd179378: dataIn1 = 32'd6560
; 
32'd179379: dataIn1 = 32'd8779
; 
32'd179380: dataIn1 = 32'd8799
; 
32'd179381: dataIn1 = 32'd8802
; 
32'd179382: dataIn1 = 32'd8809
; 
32'd179383: dataIn1 = 32'd8819
; 
32'd179384: dataIn1 = 32'd5260
; 
32'd179385: dataIn1 = 32'd6559
; 
32'd179386: dataIn1 = 32'd8781
; 
32'd179387: dataIn1 = 32'd8800
; 
32'd179388: dataIn1 = 32'd8803
; 
32'd179389: dataIn1 = 32'd8827
; 
32'd179390: dataIn1 = 32'd8842
; 
32'd179391: dataIn1 = 32'd2731
; 
32'd179392: dataIn1 = 32'd6560
; 
32'd179393: dataIn1 = 32'd8647
; 
32'd179394: dataIn1 = 32'd8801
; 
32'd179395: dataIn1 = 32'd8804
; 
32'd179396: dataIn1 = 32'd8805
; 
32'd179397: dataIn1 = 32'd8821
; 
32'd179398: dataIn1 = 32'd2731
; 
32'd179399: dataIn1 = 32'd6559
; 
32'd179400: dataIn1 = 32'd8673
; 
32'd179401: dataIn1 = 32'd8801
; 
32'd179402: dataIn1 = 32'd8804
; 
32'd179403: dataIn1 = 32'd8805
; 
32'd179404: dataIn1 = 32'd8843
; 
32'd179405: dataIn1 = 32'd6562
; 
32'd179406: dataIn1 = 32'd6563
; 
32'd179407: dataIn1 = 32'd8806
; 
32'd179408: dataIn1 = 32'd8807
; 
32'd179409: dataIn1 = 32'd8808
; 
32'd179410: dataIn1 = 32'd8809
; 
32'd179411: dataIn1 = 32'd8810
; 
32'd179412: dataIn1 = 32'd6561
; 
32'd179413: dataIn1 = 32'd6563
; 
32'd179414: dataIn1 = 32'd8806
; 
32'd179415: dataIn1 = 32'd8807
; 
32'd179416: dataIn1 = 32'd8808
; 
32'd179417: dataIn1 = 32'd8811
; 
32'd179418: dataIn1 = 32'd8812
; 
32'd179419: dataIn1 = 32'd6561
; 
32'd179420: dataIn1 = 32'd6562
; 
32'd179421: dataIn1 = 32'd8806
; 
32'd179422: dataIn1 = 32'd8807
; 
32'd179423: dataIn1 = 32'd8808
; 
32'd179424: dataIn1 = 32'd8813
; 
32'd179425: dataIn1 = 32'd8814
; 
32'd179426: dataIn1 = 32'd5259
; 
32'd179427: dataIn1 = 32'd6563
; 
32'd179428: dataIn1 = 32'd8802
; 
32'd179429: dataIn1 = 32'd8806
; 
32'd179430: dataIn1 = 32'd8809
; 
32'd179431: dataIn1 = 32'd8810
; 
32'd179432: dataIn1 = 32'd8819
; 
32'd179433: dataIn1 = 32'd5259
; 
32'd179434: dataIn1 = 32'd6562
; 
32'd179435: dataIn1 = 32'd8795
; 
32'd179436: dataIn1 = 32'd8806
; 
32'd179437: dataIn1 = 32'd8809
; 
32'd179438: dataIn1 = 32'd8810
; 
32'd179439: dataIn1 = 32'd8815
; 
32'd179440: dataIn1 = 32'd5248
; 
32'd179441: dataIn1 = 32'd6563
; 
32'd179442: dataIn1 = 32'd8646
; 
32'd179443: dataIn1 = 32'd8807
; 
32'd179444: dataIn1 = 32'd8811
; 
32'd179445: dataIn1 = 32'd8812
; 
32'd179446: dataIn1 = 32'd8820
; 
32'd179447: dataIn1 = 32'd5248
; 
32'd179448: dataIn1 = 32'd6561
; 
32'd179449: dataIn1 = 32'd6785
; 
32'd179450: dataIn1 = 32'd8807
; 
32'd179451: dataIn1 = 32'd8811
; 
32'd179452: dataIn1 = 32'd8812
; 
32'd179453: dataIn1 = 32'd5262
; 
32'd179454: dataIn1 = 32'd6562
; 
32'd179455: dataIn1 = 32'd8808
; 
32'd179456: dataIn1 = 32'd8813
; 
32'd179457: dataIn1 = 32'd8814
; 
32'd179458: dataIn1 = 32'd8817
; 
32'd179459: dataIn1 = 32'd8818
; 
32'd179460: dataIn1 = 32'd5262
; 
32'd179461: dataIn1 = 32'd6561
; 
32'd179462: dataIn1 = 32'd6784
; 
32'd179463: dataIn1 = 32'd8808
; 
32'd179464: dataIn1 = 32'd8813
; 
32'd179465: dataIn1 = 32'd8814
; 
32'd179466: dataIn1 = 32'd6558
; 
32'd179467: dataIn1 = 32'd6562
; 
32'd179468: dataIn1 = 32'd8795
; 
32'd179469: dataIn1 = 32'd8810
; 
32'd179470: dataIn1 = 32'd8815
; 
32'd179471: dataIn1 = 32'd8816
; 
32'd179472: dataIn1 = 32'd8817
; 
32'd179473: dataIn1 = 32'd6558
; 
32'd179474: dataIn1 = 32'd6564
; 
32'd179475: dataIn1 = 32'd8796
; 
32'd179476: dataIn1 = 32'd8815
; 
32'd179477: dataIn1 = 32'd8816
; 
32'd179478: dataIn1 = 32'd8817
; 
32'd179479: dataIn1 = 32'd9276
; 
32'd179480: dataIn1 = 32'd6562
; 
32'd179481: dataIn1 = 32'd6564
; 
32'd179482: dataIn1 = 32'd8813
; 
32'd179483: dataIn1 = 32'd8815
; 
32'd179484: dataIn1 = 32'd8816
; 
32'd179485: dataIn1 = 32'd8817
; 
32'd179486: dataIn1 = 32'd8818
; 
32'd179487: dataIn1 = 32'd5262
; 
32'd179488: dataIn1 = 32'd6564
; 
32'd179489: dataIn1 = 32'd8813
; 
32'd179490: dataIn1 = 32'd8817
; 
32'd179491: dataIn1 = 32'd8818
; 
32'd179492: dataIn1 = 32'd9442
; 
32'd179493: dataIn1 = 32'd9447
; 
32'd179494: dataIn1 = 32'd6560
; 
32'd179495: dataIn1 = 32'd6563
; 
32'd179496: dataIn1 = 32'd8802
; 
32'd179497: dataIn1 = 32'd8809
; 
32'd179498: dataIn1 = 32'd8819
; 
32'd179499: dataIn1 = 32'd8820
; 
32'd179500: dataIn1 = 32'd8821
; 
32'd179501: dataIn1 = 32'd6520
; 
32'd179502: dataIn1 = 32'd6563
; 
32'd179503: dataIn1 = 32'd8646
; 
32'd179504: dataIn1 = 32'd8811
; 
32'd179505: dataIn1 = 32'd8819
; 
32'd179506: dataIn1 = 32'd8820
; 
32'd179507: dataIn1 = 32'd8821
; 
32'd179508: dataIn1 = 32'd6520
; 
32'd179509: dataIn1 = 32'd6560
; 
32'd179510: dataIn1 = 32'd8647
; 
32'd179511: dataIn1 = 32'd8804
; 
32'd179512: dataIn1 = 32'd8819
; 
32'd179513: dataIn1 = 32'd8820
; 
32'd179514: dataIn1 = 32'd8821
; 
32'd179515: dataIn1 = 32'd6566
; 
32'd179516: dataIn1 = 32'd6567
; 
32'd179517: dataIn1 = 32'd8822
; 
32'd179518: dataIn1 = 32'd8823
; 
32'd179519: dataIn1 = 32'd8824
; 
32'd179520: dataIn1 = 32'd8825
; 
32'd179521: dataIn1 = 32'd8826
; 
32'd179522: dataIn1 = 32'd6565
; 
32'd179523: dataIn1 = 32'd6567
; 
32'd179524: dataIn1 = 32'd8822
; 
32'd179525: dataIn1 = 32'd8823
; 
32'd179526: dataIn1 = 32'd8824
; 
32'd179527: dataIn1 = 32'd8827
; 
32'd179528: dataIn1 = 32'd8828
; 
32'd179529: dataIn1 = 32'd6565
; 
32'd179530: dataIn1 = 32'd6566
; 
32'd179531: dataIn1 = 32'd8822
; 
32'd179532: dataIn1 = 32'd8823
; 
32'd179533: dataIn1 = 32'd8824
; 
32'd179534: dataIn1 = 32'd8829
; 
32'd179535: dataIn1 = 32'd8830
; 
32'd179536: dataIn1 = 32'd5250
; 
32'd179537: dataIn1 = 32'd6567
; 
32'd179538: dataIn1 = 32'd8672
; 
32'd179539: dataIn1 = 32'd8822
; 
32'd179540: dataIn1 = 32'd8825
; 
32'd179541: dataIn1 = 32'd8826
; 
32'd179542: dataIn1 = 32'd8841
; 
32'd179543: dataIn1 = 32'd5250
; 
32'd179544: dataIn1 = 32'd6566
; 
32'd179545: dataIn1 = 32'd8665
; 
32'd179546: dataIn1 = 32'd8822
; 
32'd179547: dataIn1 = 32'd8825
; 
32'd179548: dataIn1 = 32'd8826
; 
32'd179549: dataIn1 = 32'd8836
; 
32'd179550: dataIn1 = 32'd5260
; 
32'd179551: dataIn1 = 32'd6567
; 
32'd179552: dataIn1 = 32'd8803
; 
32'd179553: dataIn1 = 32'd8823
; 
32'd179554: dataIn1 = 32'd8827
; 
32'd179555: dataIn1 = 32'd8828
; 
32'd179556: dataIn1 = 32'd8842
; 
32'd179557: dataIn1 = 32'd5260
; 
32'd179558: dataIn1 = 32'd6565
; 
32'd179559: dataIn1 = 32'd8790
; 
32'd179560: dataIn1 = 32'd8823
; 
32'd179561: dataIn1 = 32'd8827
; 
32'd179562: dataIn1 = 32'd8828
; 
32'd179563: dataIn1 = 32'd8832
; 
32'd179564: dataIn1 = 32'd2690
; 
32'd179565: dataIn1 = 32'd6566
; 
32'd179566: dataIn1 = 32'd8824
; 
32'd179567: dataIn1 = 32'd8829
; 
32'd179568: dataIn1 = 32'd8830
; 
32'd179569: dataIn1 = 32'd8838
; 
32'd179570: dataIn1 = 32'd8840
; 
32'd179571: dataIn1 = 32'd2690
; 
32'd179572: dataIn1 = 32'd6565
; 
32'd179573: dataIn1 = 32'd8824
; 
32'd179574: dataIn1 = 32'd8829
; 
32'd179575: dataIn1 = 32'd8830
; 
32'd179576: dataIn1 = 32'd8833
; 
32'd179577: dataIn1 = 32'd8835
; 
32'd179578: dataIn1 = 32'd5106
; 
32'd179579: dataIn1 = 32'd6556
; 
32'd179580: dataIn1 = 32'd8788
; 
32'd179581: dataIn1 = 32'd8831
; 
32'd179582: dataIn1 = 32'd8832
; 
32'd179583: dataIn1 = 32'd8833
; 
32'd179584: dataIn1 = 32'd8834
; 
32'd179585: dataIn1 = 32'd6556
; 
32'd179586: dataIn1 = 32'd6565
; 
32'd179587: dataIn1 = 32'd8790
; 
32'd179588: dataIn1 = 32'd8828
; 
32'd179589: dataIn1 = 32'd8831
; 
32'd179590: dataIn1 = 32'd8832
; 
32'd179591: dataIn1 = 32'd8833
; 
32'd179592: dataIn1 = 32'd5106
; 
32'd179593: dataIn1 = 32'd6565
; 
32'd179594: dataIn1 = 32'd8830
; 
32'd179595: dataIn1 = 32'd8831
; 
32'd179596: dataIn1 = 32'd8832
; 
32'd179597: dataIn1 = 32'd8833
; 
32'd179598: dataIn1 = 32'd8835
; 
32'd179599: dataIn1 = 32'd1118
; 
32'd179600: dataIn1 = 32'd5099
; 
32'd179601: dataIn1 = 32'd5106
; 
32'd179602: dataIn1 = 32'd8788
; 
32'd179603: dataIn1 = 32'd8831
; 
32'd179604: dataIn1 = 32'd8834
; 
32'd179605: dataIn1 = 32'd2690
; 
32'd179606: dataIn1 = 32'd5103
; 
32'd179607: dataIn1 = 32'd5106
; 
32'd179608: dataIn1 = 32'd8830
; 
32'd179609: dataIn1 = 32'd8833
; 
32'd179610: dataIn1 = 32'd8835
; 
32'd179611: dataIn1 = 32'd6527
; 
32'd179612: dataIn1 = 32'd6566
; 
32'd179613: dataIn1 = 32'd8665
; 
32'd179614: dataIn1 = 32'd8826
; 
32'd179615: dataIn1 = 32'd8836
; 
32'd179616: dataIn1 = 32'd8837
; 
32'd179617: dataIn1 = 32'd8838
; 
32'd179618: dataIn1 = 32'd5105
; 
32'd179619: dataIn1 = 32'd6527
; 
32'd179620: dataIn1 = 32'd8666
; 
32'd179621: dataIn1 = 32'd8836
; 
32'd179622: dataIn1 = 32'd8837
; 
32'd179623: dataIn1 = 32'd8838
; 
32'd179624: dataIn1 = 32'd8839
; 
32'd179625: dataIn1 = 32'd5105
; 
32'd179626: dataIn1 = 32'd6566
; 
32'd179627: dataIn1 = 32'd8829
; 
32'd179628: dataIn1 = 32'd8836
; 
32'd179629: dataIn1 = 32'd8837
; 
32'd179630: dataIn1 = 32'd8838
; 
32'd179631: dataIn1 = 32'd8840
; 
32'd179632: dataIn1 = 32'd148
; 
32'd179633: dataIn1 = 32'd4778
; 
32'd179634: dataIn1 = 32'd5105
; 
32'd179635: dataIn1 = 32'd8666
; 
32'd179636: dataIn1 = 32'd8837
; 
32'd179637: dataIn1 = 32'd8839
; 
32'd179638: dataIn1 = 32'd2690
; 
32'd179639: dataIn1 = 32'd5102
; 
32'd179640: dataIn1 = 32'd5105
; 
32'd179641: dataIn1 = 32'd8829
; 
32'd179642: dataIn1 = 32'd8838
; 
32'd179643: dataIn1 = 32'd8840
; 
32'd179644: dataIn1 = 32'd6528
; 
32'd179645: dataIn1 = 32'd6567
; 
32'd179646: dataIn1 = 32'd8672
; 
32'd179647: dataIn1 = 32'd8825
; 
32'd179648: dataIn1 = 32'd8841
; 
32'd179649: dataIn1 = 32'd8842
; 
32'd179650: dataIn1 = 32'd8843
; 
32'd179651: dataIn1 = 32'd6559
; 
32'd179652: dataIn1 = 32'd6567
; 
32'd179653: dataIn1 = 32'd8803
; 
32'd179654: dataIn1 = 32'd8827
; 
32'd179655: dataIn1 = 32'd8841
; 
32'd179656: dataIn1 = 32'd8842
; 
32'd179657: dataIn1 = 32'd8843
; 
32'd179658: dataIn1 = 32'd6528
; 
32'd179659: dataIn1 = 32'd6559
; 
32'd179660: dataIn1 = 32'd8673
; 
32'd179661: dataIn1 = 32'd8805
; 
32'd179662: dataIn1 = 32'd8841
; 
32'd179663: dataIn1 = 32'd8842
; 
32'd179664: dataIn1 = 32'd8843
; 
32'd179665: dataIn1 = 32'd6569
; 
32'd179666: dataIn1 = 32'd6570
; 
32'd179667: dataIn1 = 32'd8844
; 
32'd179668: dataIn1 = 32'd8845
; 
32'd179669: dataIn1 = 32'd8846
; 
32'd179670: dataIn1 = 32'd8847
; 
32'd179671: dataIn1 = 32'd8848
; 
32'd179672: dataIn1 = 32'd6568
; 
32'd179673: dataIn1 = 32'd6570
; 
32'd179674: dataIn1 = 32'd8844
; 
32'd179675: dataIn1 = 32'd8845
; 
32'd179676: dataIn1 = 32'd8846
; 
32'd179677: dataIn1 = 32'd8849
; 
32'd179678: dataIn1 = 32'd8850
; 
32'd179679: dataIn1 = 32'd6568
; 
32'd179680: dataIn1 = 32'd6569
; 
32'd179681: dataIn1 = 32'd8844
; 
32'd179682: dataIn1 = 32'd8845
; 
32'd179683: dataIn1 = 32'd8846
; 
32'd179684: dataIn1 = 32'd8851
; 
32'd179685: dataIn1 = 32'd8852
; 
32'd179686: dataIn1 = 32'd5263
; 
32'd179687: dataIn1 = 32'd6570
; 
32'd179688: dataIn1 = 32'd8844
; 
32'd179689: dataIn1 = 32'd8847
; 
32'd179690: dataIn1 = 32'd8848
; 
32'd179691: dataIn1 = 32'd8863
; 
32'd179692: dataIn1 = 32'd8866
; 
32'd179693: dataIn1 = 32'd5263
; 
32'd179694: dataIn1 = 32'd6569
; 
32'd179695: dataIn1 = 32'd8844
; 
32'd179696: dataIn1 = 32'd8847
; 
32'd179697: dataIn1 = 32'd8848
; 
32'd179698: dataIn1 = 32'd8858
; 
32'd179699: dataIn1 = 32'd8861
; 
32'd179700: dataIn1 = 32'd2691
; 
32'd179701: dataIn1 = 32'd6570
; 
32'd179702: dataIn1 = 32'd8845
; 
32'd179703: dataIn1 = 32'd8849
; 
32'd179704: dataIn1 = 32'd8850
; 
32'd179705: dataIn1 = 32'd8864
; 
32'd179706: dataIn1 = 32'd8867
; 
32'd179707: dataIn1 = 32'd2691
; 
32'd179708: dataIn1 = 32'd6568
; 
32'd179709: dataIn1 = 32'd8845
; 
32'd179710: dataIn1 = 32'd8849
; 
32'd179711: dataIn1 = 32'd8850
; 
32'd179712: dataIn1 = 32'd8854
; 
32'd179713: dataIn1 = 32'd8857
; 
32'd179714: dataIn1 = 32'd5261
; 
32'd179715: dataIn1 = 32'd6569
; 
32'd179716: dataIn1 = 32'd8798
; 
32'd179717: dataIn1 = 32'd8846
; 
32'd179718: dataIn1 = 32'd8851
; 
32'd179719: dataIn1 = 32'd8852
; 
32'd179720: dataIn1 = 32'd8860
; 
32'd179721: dataIn1 = 32'd5261
; 
32'd179722: dataIn1 = 32'd6568
; 
32'd179723: dataIn1 = 32'd8791
; 
32'd179724: dataIn1 = 32'd8846
; 
32'd179725: dataIn1 = 32'd8851
; 
32'd179726: dataIn1 = 32'd8852
; 
32'd179727: dataIn1 = 32'd8855
; 
32'd179728: dataIn1 = 32'd5110
; 
32'd179729: dataIn1 = 32'd6555
; 
32'd179730: dataIn1 = 32'd8789
; 
32'd179731: dataIn1 = 32'd8853
; 
32'd179732: dataIn1 = 32'd8854
; 
32'd179733: dataIn1 = 32'd8855
; 
32'd179734: dataIn1 = 32'd8856
; 
32'd179735: dataIn1 = 32'd5110
; 
32'd179736: dataIn1 = 32'd6568
; 
32'd179737: dataIn1 = 32'd8850
; 
32'd179738: dataIn1 = 32'd8853
; 
32'd179739: dataIn1 = 32'd8854
; 
32'd179740: dataIn1 = 32'd8855
; 
32'd179741: dataIn1 = 32'd8857
; 
32'd179742: dataIn1 = 32'd6555
; 
32'd179743: dataIn1 = 32'd6568
; 
32'd179744: dataIn1 = 32'd8791
; 
32'd179745: dataIn1 = 32'd8852
; 
32'd179746: dataIn1 = 32'd8853
; 
32'd179747: dataIn1 = 32'd8854
; 
32'd179748: dataIn1 = 32'd8855
; 
32'd179749: dataIn1 = 32'd1118
; 
32'd179750: dataIn1 = 32'd5098
; 
32'd179751: dataIn1 = 32'd5110
; 
32'd179752: dataIn1 = 32'd8789
; 
32'd179753: dataIn1 = 32'd8853
; 
32'd179754: dataIn1 = 32'd8856
; 
32'd179755: dataIn1 = 32'd2691
; 
32'd179756: dataIn1 = 32'd5108
; 
32'd179757: dataIn1 = 32'd5110
; 
32'd179758: dataIn1 = 32'd8850
; 
32'd179759: dataIn1 = 32'd8854
; 
32'd179760: dataIn1 = 32'd8857
; 
32'd179761: dataIn1 = 32'd6569
; 
32'd179762: dataIn1 = 32'd6571
; 
32'd179763: dataIn1 = 32'd8848
; 
32'd179764: dataIn1 = 32'd8858
; 
32'd179765: dataIn1 = 32'd8859
; 
32'd179766: dataIn1 = 32'd8860
; 
32'd179767: dataIn1 = 32'd8861
; 
32'd179768: dataIn1 = 32'd6557
; 
32'd179769: dataIn1 = 32'd6571
; 
32'd179770: dataIn1 = 32'd8797
; 
32'd179771: dataIn1 = 32'd8858
; 
32'd179772: dataIn1 = 32'd8859
; 
32'd179773: dataIn1 = 32'd8860
; 
32'd179774: dataIn1 = 32'd8862
; 
32'd179775: dataIn1 = 32'd6557
; 
32'd179776: dataIn1 = 32'd6569
; 
32'd179777: dataIn1 = 32'd8798
; 
32'd179778: dataIn1 = 32'd8851
; 
32'd179779: dataIn1 = 32'd8858
; 
32'd179780: dataIn1 = 32'd8859
; 
32'd179781: dataIn1 = 32'd8860
; 
32'd179782: dataIn1 = 32'd5263
; 
32'd179783: dataIn1 = 32'd6571
; 
32'd179784: dataIn1 = 32'd8848
; 
32'd179785: dataIn1 = 32'd8858
; 
32'd179786: dataIn1 = 32'd8861
; 
32'd179787: dataIn1 = 32'd9421
; 
32'd179788: dataIn1 = 32'd9429
; 
32'd179789: dataIn1 = 32'd2733
; 
32'd179790: dataIn1 = 32'd6571
; 
32'd179791: dataIn1 = 32'd8797
; 
32'd179792: dataIn1 = 32'd8859
; 
32'd179793: dataIn1 = 32'd8862
; 
32'd179794: dataIn1 = 32'd9404
; 
32'd179795: dataIn1 = 32'd9428
; 
32'd179796: dataIn1 = 32'd6570
; 
32'd179797: dataIn1 = 32'd6572
; 
32'd179798: dataIn1 = 32'd8847
; 
32'd179799: dataIn1 = 32'd8863
; 
32'd179800: dataIn1 = 32'd8864
; 
32'd179801: dataIn1 = 32'd8865
; 
32'd179802: dataIn1 = 32'd8866
; 
32'd179803: dataIn1 = 32'd5111
; 
32'd179804: dataIn1 = 32'd6570
; 
32'd179805: dataIn1 = 32'd8849
; 
32'd179806: dataIn1 = 32'd8863
; 
32'd179807: dataIn1 = 32'd8864
; 
32'd179808: dataIn1 = 32'd8865
; 
32'd179809: dataIn1 = 32'd8867
; 
32'd179810: dataIn1 = 32'd5111
; 
32'd179811: dataIn1 = 32'd6572
; 
32'd179812: dataIn1 = 32'd8863
; 
32'd179813: dataIn1 = 32'd8864
; 
32'd179814: dataIn1 = 32'd8865
; 
32'd179815: dataIn1 = 32'd8868
; 
32'd179816: dataIn1 = 32'd8869
; 
32'd179817: dataIn1 = 32'd5263
; 
32'd179818: dataIn1 = 32'd6572
; 
32'd179819: dataIn1 = 32'd8847
; 
32'd179820: dataIn1 = 32'd8863
; 
32'd179821: dataIn1 = 32'd8866
; 
32'd179822: dataIn1 = 32'd9422
; 
32'd179823: dataIn1 = 32'd9425
; 
32'd179824: dataIn1 = 32'd2691
; 
32'd179825: dataIn1 = 32'd5109
; 
32'd179826: dataIn1 = 32'd5111
; 
32'd179827: dataIn1 = 32'd8849
; 
32'd179828: dataIn1 = 32'd8864
; 
32'd179829: dataIn1 = 32'd8867
; 
32'd179830: dataIn1 = 32'd12
; 
32'd179831: dataIn1 = 32'd6572
; 
32'd179832: dataIn1 = 32'd8865
; 
32'd179833: dataIn1 = 32'd8868
; 
32'd179834: dataIn1 = 32'd8869
; 
32'd179835: dataIn1 = 32'd9423
; 
32'd179836: dataIn1 = 32'd9448
; 
32'd179837: dataIn1 = 32'd12
; 
32'd179838: dataIn1 = 32'd4788
; 
32'd179839: dataIn1 = 32'd5111
; 
32'd179840: dataIn1 = 32'd8865
; 
32'd179841: dataIn1 = 32'd8868
; 
32'd179842: dataIn1 = 32'd8869
; 
32'd179843: dataIn1 = 32'd6574
; 
32'd179844: dataIn1 = 32'd6575
; 
32'd179845: dataIn1 = 32'd8870
; 
32'd179846: dataIn1 = 32'd8871
; 
32'd179847: dataIn1 = 32'd8872
; 
32'd179848: dataIn1 = 32'd8873
; 
32'd179849: dataIn1 = 32'd8874
; 
32'd179850: dataIn1 = 32'd6573
; 
32'd179851: dataIn1 = 32'd6575
; 
32'd179852: dataIn1 = 32'd8870
; 
32'd179853: dataIn1 = 32'd8871
; 
32'd179854: dataIn1 = 32'd8872
; 
32'd179855: dataIn1 = 32'd8875
; 
32'd179856: dataIn1 = 32'd8876
; 
32'd179857: dataIn1 = 32'd6573
; 
32'd179858: dataIn1 = 32'd6574
; 
32'd179859: dataIn1 = 32'd8870
; 
32'd179860: dataIn1 = 32'd8871
; 
32'd179861: dataIn1 = 32'd8872
; 
32'd179862: dataIn1 = 32'd8877
; 
32'd179863: dataIn1 = 32'd8878
; 
32'd179864: dataIn1 = 32'd5264
; 
32'd179865: dataIn1 = 32'd6575
; 
32'd179866: dataIn1 = 32'd8870
; 
32'd179867: dataIn1 = 32'd8873
; 
32'd179868: dataIn1 = 32'd8874
; 
32'd179869: dataIn1 = 32'd8886
; 
32'd179870: dataIn1 = 32'd8889
; 
32'd179871: dataIn1 = 32'd5264
; 
32'd179872: dataIn1 = 32'd6574
; 
32'd179873: dataIn1 = 32'd8870
; 
32'd179874: dataIn1 = 32'd8873
; 
32'd179875: dataIn1 = 32'd8874
; 
32'd179876: dataIn1 = 32'd8879
; 
32'd179877: dataIn1 = 32'd8882
; 
32'd179878: dataIn1 = 32'd5265
; 
32'd179879: dataIn1 = 32'd6575
; 
32'd179880: dataIn1 = 32'd8871
; 
32'd179881: dataIn1 = 32'd8875
; 
32'd179882: dataIn1 = 32'd8876
; 
32'd179883: dataIn1 = 32'd8887
; 
32'd179884: dataIn1 = 32'd8890
; 
32'd179885: dataIn1 = 32'd5265
; 
32'd179886: dataIn1 = 32'd6573
; 
32'd179887: dataIn1 = 32'd6577
; 
32'd179888: dataIn1 = 32'd8871
; 
32'd179889: dataIn1 = 32'd8875
; 
32'd179890: dataIn1 = 32'd8876
; 
32'd179891: dataIn1 = 32'd5266
; 
32'd179892: dataIn1 = 32'd6574
; 
32'd179893: dataIn1 = 32'd8872
; 
32'd179894: dataIn1 = 32'd8877
; 
32'd179895: dataIn1 = 32'd8878
; 
32'd179896: dataIn1 = 32'd8881
; 
32'd179897: dataIn1 = 32'd8885
; 
32'd179898: dataIn1 = 32'd5266
; 
32'd179899: dataIn1 = 32'd6573
; 
32'd179900: dataIn1 = 32'd6576
; 
32'd179901: dataIn1 = 32'd8872
; 
32'd179902: dataIn1 = 32'd8877
; 
32'd179903: dataIn1 = 32'd8878
; 
32'd179904: dataIn1 = 32'd6574
; 
32'd179905: dataIn1 = 32'd6579
; 
32'd179906: dataIn1 = 32'd8874
; 
32'd179907: dataIn1 = 32'd8879
; 
32'd179908: dataIn1 = 32'd8880
; 
32'd179909: dataIn1 = 32'd8881
; 
32'd179910: dataIn1 = 32'd8882
; 
32'd179911: dataIn1 = 32'd6578
; 
32'd179912: dataIn1 = 32'd6579
; 
32'd179913: dataIn1 = 32'd8879
; 
32'd179914: dataIn1 = 32'd8880
; 
32'd179915: dataIn1 = 32'd8881
; 
32'd179916: dataIn1 = 32'd8883
; 
32'd179917: dataIn1 = 32'd8884
; 
32'd179918: dataIn1 = 32'd6574
; 
32'd179919: dataIn1 = 32'd6578
; 
32'd179920: dataIn1 = 32'd8877
; 
32'd179921: dataIn1 = 32'd8879
; 
32'd179922: dataIn1 = 32'd8880
; 
32'd179923: dataIn1 = 32'd8881
; 
32'd179924: dataIn1 = 32'd8885
; 
32'd179925: dataIn1 = 32'd5264
; 
32'd179926: dataIn1 = 32'd6579
; 
32'd179927: dataIn1 = 32'd8874
; 
32'd179928: dataIn1 = 32'd8879
; 
32'd179929: dataIn1 = 32'd8882
; 
32'd179930: dataIn1 = 32'd8897
; 
32'd179931: dataIn1 = 32'd8905
; 
32'd179932: dataIn1 = 32'd2696
; 
32'd179933: dataIn1 = 32'd6579
; 
32'd179934: dataIn1 = 32'd7219
; 
32'd179935: dataIn1 = 32'd8880
; 
32'd179936: dataIn1 = 32'd8883
; 
32'd179937: dataIn1 = 32'd8884
; 
32'd179938: dataIn1 = 32'd8906
; 
32'd179939: dataIn1 = 32'd2696
; 
32'd179940: dataIn1 = 32'd6578
; 
32'd179941: dataIn1 = 32'd7198
; 
32'd179942: dataIn1 = 32'd8880
; 
32'd179943: dataIn1 = 32'd8883
; 
32'd179944: dataIn1 = 32'd8884
; 
32'd179945: dataIn1 = 32'd8917
; 
32'd179946: dataIn1 = 32'd5266
; 
32'd179947: dataIn1 = 32'd6578
; 
32'd179948: dataIn1 = 32'd8877
; 
32'd179949: dataIn1 = 32'd8881
; 
32'd179950: dataIn1 = 32'd8885
; 
32'd179951: dataIn1 = 32'd8918
; 
32'd179952: dataIn1 = 32'd8920
; 
32'd179953: dataIn1 = 32'd6575
; 
32'd179954: dataIn1 = 32'd6581
; 
32'd179955: dataIn1 = 32'd8873
; 
32'd179956: dataIn1 = 32'd8886
; 
32'd179957: dataIn1 = 32'd8887
; 
32'd179958: dataIn1 = 32'd8888
; 
32'd179959: dataIn1 = 32'd8889
; 
32'd179960: dataIn1 = 32'd6575
; 
32'd179961: dataIn1 = 32'd6580
; 
32'd179962: dataIn1 = 32'd8875
; 
32'd179963: dataIn1 = 32'd8886
; 
32'd179964: dataIn1 = 32'd8887
; 
32'd179965: dataIn1 = 32'd8888
; 
32'd179966: dataIn1 = 32'd8890
; 
32'd179967: dataIn1 = 32'd6580
; 
32'd179968: dataIn1 = 32'd6581
; 
32'd179969: dataIn1 = 32'd8886
; 
32'd179970: dataIn1 = 32'd8887
; 
32'd179971: dataIn1 = 32'd8888
; 
32'd179972: dataIn1 = 32'd8891
; 
32'd179973: dataIn1 = 32'd8892
; 
32'd179974: dataIn1 = 32'd5264
; 
32'd179975: dataIn1 = 32'd6581
; 
32'd179976: dataIn1 = 32'd8873
; 
32'd179977: dataIn1 = 32'd8886
; 
32'd179978: dataIn1 = 32'd8889
; 
32'd179979: dataIn1 = 32'd8896
; 
32'd179980: dataIn1 = 32'd8908
; 
32'd179981: dataIn1 = 32'd5265
; 
32'd179982: dataIn1 = 32'd6580
; 
32'd179983: dataIn1 = 32'd8875
; 
32'd179984: dataIn1 = 32'd8887
; 
32'd179985: dataIn1 = 32'd8890
; 
32'd179986: dataIn1 = 32'd8912
; 
32'd179987: dataIn1 = 32'd8915
; 
32'd179988: dataIn1 = 32'd2322
; 
32'd179989: dataIn1 = 32'd6581
; 
32'd179990: dataIn1 = 32'd6949
; 
32'd179991: dataIn1 = 32'd8888
; 
32'd179992: dataIn1 = 32'd8891
; 
32'd179993: dataIn1 = 32'd8892
; 
32'd179994: dataIn1 = 32'd8910
; 
32'd179995: dataIn1 = 32'd2322
; 
32'd179996: dataIn1 = 32'd6580
; 
32'd179997: dataIn1 = 32'd6988
; 
32'd179998: dataIn1 = 32'd8888
; 
32'd179999: dataIn1 = 32'd8891
; 
32'd180000: dataIn1 = 32'd8892
; 
32'd180001: dataIn1 = 32'd8913
; 
32'd180002: dataIn1 = 32'd6583
; 
32'd180003: dataIn1 = 32'd6584
; 
32'd180004: dataIn1 = 32'd8893
; 
32'd180005: dataIn1 = 32'd8894
; 
32'd180006: dataIn1 = 32'd8895
; 
32'd180007: dataIn1 = 32'd8896
; 
32'd180008: dataIn1 = 32'd8897
; 
32'd180009: dataIn1 = 32'd6582
; 
32'd180010: dataIn1 = 32'd6584
; 
32'd180011: dataIn1 = 32'd8893
; 
32'd180012: dataIn1 = 32'd8894
; 
32'd180013: dataIn1 = 32'd8895
; 
32'd180014: dataIn1 = 32'd8898
; 
32'd180015: dataIn1 = 32'd8899
; 
32'd180016: dataIn1 = 32'd6582
; 
32'd180017: dataIn1 = 32'd6583
; 
32'd180018: dataIn1 = 32'd8893
; 
32'd180019: dataIn1 = 32'd8894
; 
32'd180020: dataIn1 = 32'd8895
; 
32'd180021: dataIn1 = 32'd8900
; 
32'd180022: dataIn1 = 32'd8901
; 
32'd180023: dataIn1 = 32'd5264
; 
32'd180024: dataIn1 = 32'd6584
; 
32'd180025: dataIn1 = 32'd8889
; 
32'd180026: dataIn1 = 32'd8893
; 
32'd180027: dataIn1 = 32'd8896
; 
32'd180028: dataIn1 = 32'd8897
; 
32'd180029: dataIn1 = 32'd8908
; 
32'd180030: dataIn1 = 32'd5264
; 
32'd180031: dataIn1 = 32'd6583
; 
32'd180032: dataIn1 = 32'd8882
; 
32'd180033: dataIn1 = 32'd8893
; 
32'd180034: dataIn1 = 32'd8896
; 
32'd180035: dataIn1 = 32'd8897
; 
32'd180036: dataIn1 = 32'd8905
; 
32'd180037: dataIn1 = 32'd3975
; 
32'd180038: dataIn1 = 32'd6584
; 
32'd180039: dataIn1 = 32'd6950
; 
32'd180040: dataIn1 = 32'd8894
; 
32'd180041: dataIn1 = 32'd8898
; 
32'd180042: dataIn1 = 32'd8899
; 
32'd180043: dataIn1 = 32'd8909
; 
32'd180044: dataIn1 = 32'd3975
; 
32'd180045: dataIn1 = 32'd6582
; 
32'd180046: dataIn1 = 32'd6944
; 
32'd180047: dataIn1 = 32'd8894
; 
32'd180048: dataIn1 = 32'd8898
; 
32'd180049: dataIn1 = 32'd8899
; 
32'd180050: dataIn1 = 32'd8903
; 
32'd180051: dataIn1 = 32'd5130
; 
32'd180052: dataIn1 = 32'd6583
; 
32'd180053: dataIn1 = 32'd7218
; 
32'd180054: dataIn1 = 32'd8895
; 
32'd180055: dataIn1 = 32'd8900
; 
32'd180056: dataIn1 = 32'd8901
; 
32'd180057: dataIn1 = 32'd8907
; 
32'd180058: dataIn1 = 32'd5130
; 
32'd180059: dataIn1 = 32'd6582
; 
32'd180060: dataIn1 = 32'd7221
; 
32'd180061: dataIn1 = 32'd8895
; 
32'd180062: dataIn1 = 32'd8900
; 
32'd180063: dataIn1 = 32'd8901
; 
32'd180064: dataIn1 = 32'd8904
; 
32'd180065: dataIn1 = 32'd4
; 
32'd180066: dataIn1 = 32'd5861
; 
32'd180067: dataIn1 = 32'd6140
; 
32'd180068: dataIn1 = 32'd8902
; 
32'd180069: dataIn1 = 32'd8903
; 
32'd180070: dataIn1 = 32'd8904
; 
32'd180071: dataIn1 = 32'd5861
; 
32'd180072: dataIn1 = 32'd6582
; 
32'd180073: dataIn1 = 32'd6944
; 
32'd180074: dataIn1 = 32'd8899
; 
32'd180075: dataIn1 = 32'd8902
; 
32'd180076: dataIn1 = 32'd8903
; 
32'd180077: dataIn1 = 32'd8904
; 
32'd180078: dataIn1 = 32'd6140
; 
32'd180079: dataIn1 = 32'd6582
; 
32'd180080: dataIn1 = 32'd7221
; 
32'd180081: dataIn1 = 32'd8901
; 
32'd180082: dataIn1 = 32'd8902
; 
32'd180083: dataIn1 = 32'd8903
; 
32'd180084: dataIn1 = 32'd8904
; 
32'd180085: dataIn1 = 32'd6579
; 
32'd180086: dataIn1 = 32'd6583
; 
32'd180087: dataIn1 = 32'd8882
; 
32'd180088: dataIn1 = 32'd8897
; 
32'd180089: dataIn1 = 32'd8905
; 
32'd180090: dataIn1 = 32'd8906
; 
32'd180091: dataIn1 = 32'd8907
; 
32'd180092: dataIn1 = 32'd6139
; 
32'd180093: dataIn1 = 32'd6579
; 
32'd180094: dataIn1 = 32'd7219
; 
32'd180095: dataIn1 = 32'd8883
; 
32'd180096: dataIn1 = 32'd8905
; 
32'd180097: dataIn1 = 32'd8906
; 
32'd180098: dataIn1 = 32'd8907
; 
32'd180099: dataIn1 = 32'd6139
; 
32'd180100: dataIn1 = 32'd6583
; 
32'd180101: dataIn1 = 32'd7218
; 
32'd180102: dataIn1 = 32'd8900
; 
32'd180103: dataIn1 = 32'd8905
; 
32'd180104: dataIn1 = 32'd8906
; 
32'd180105: dataIn1 = 32'd8907
; 
32'd180106: dataIn1 = 32'd6581
; 
32'd180107: dataIn1 = 32'd6584
; 
32'd180108: dataIn1 = 32'd8889
; 
32'd180109: dataIn1 = 32'd8896
; 
32'd180110: dataIn1 = 32'd8908
; 
32'd180111: dataIn1 = 32'd8909
; 
32'd180112: dataIn1 = 32'd8910
; 
32'd180113: dataIn1 = 32'd5862
; 
32'd180114: dataIn1 = 32'd6584
; 
32'd180115: dataIn1 = 32'd6950
; 
32'd180116: dataIn1 = 32'd8898
; 
32'd180117: dataIn1 = 32'd8908
; 
32'd180118: dataIn1 = 32'd8909
; 
32'd180119: dataIn1 = 32'd8910
; 
32'd180120: dataIn1 = 32'd5862
; 
32'd180121: dataIn1 = 32'd6581
; 
32'd180122: dataIn1 = 32'd6949
; 
32'd180123: dataIn1 = 32'd8891
; 
32'd180124: dataIn1 = 32'd8908
; 
32'd180125: dataIn1 = 32'd8909
; 
32'd180126: dataIn1 = 32'd8910
; 
32'd180127: dataIn1 = 32'd5869
; 
32'd180128: dataIn1 = 32'd6587
; 
32'd180129: dataIn1 = 32'd6987
; 
32'd180130: dataIn1 = 32'd8911
; 
32'd180131: dataIn1 = 32'd8912
; 
32'd180132: dataIn1 = 32'd8913
; 
32'd180133: dataIn1 = 32'd8914
; 
32'd180134: dataIn1 = 32'd6580
; 
32'd180135: dataIn1 = 32'd6587
; 
32'd180136: dataIn1 = 32'd8890
; 
32'd180137: dataIn1 = 32'd8911
; 
32'd180138: dataIn1 = 32'd8912
; 
32'd180139: dataIn1 = 32'd8913
; 
32'd180140: dataIn1 = 32'd8915
; 
32'd180141: dataIn1 = 32'd5869
; 
32'd180142: dataIn1 = 32'd6580
; 
32'd180143: dataIn1 = 32'd6988
; 
32'd180144: dataIn1 = 32'd8892
; 
32'd180145: dataIn1 = 32'd8911
; 
32'd180146: dataIn1 = 32'd8912
; 
32'd180147: dataIn1 = 32'd8913
; 
32'd180148: dataIn1 = 32'd3976
; 
32'd180149: dataIn1 = 32'd6586
; 
32'd180150: dataIn1 = 32'd6587
; 
32'd180151: dataIn1 = 32'd6987
; 
32'd180152: dataIn1 = 32'd8911
; 
32'd180153: dataIn1 = 32'd8914
; 
32'd180154: dataIn1 = 32'd5265
; 
32'd180155: dataIn1 = 32'd6585
; 
32'd180156: dataIn1 = 32'd6587
; 
32'd180157: dataIn1 = 32'd8890
; 
32'd180158: dataIn1 = 32'd8912
; 
32'd180159: dataIn1 = 32'd8915
; 
32'd180160: dataIn1 = 32'd6132
; 
32'd180161: dataIn1 = 32'd6591
; 
32'd180162: dataIn1 = 32'd7199
; 
32'd180163: dataIn1 = 32'd8916
; 
32'd180164: dataIn1 = 32'd8917
; 
32'd180165: dataIn1 = 32'd8918
; 
32'd180166: dataIn1 = 32'd8919
; 
32'd180167: dataIn1 = 32'd6132
; 
32'd180168: dataIn1 = 32'd6578
; 
32'd180169: dataIn1 = 32'd7198
; 
32'd180170: dataIn1 = 32'd8884
; 
32'd180171: dataIn1 = 32'd8916
; 
32'd180172: dataIn1 = 32'd8917
; 
32'd180173: dataIn1 = 32'd8918
; 
32'd180174: dataIn1 = 32'd6578
; 
32'd180175: dataIn1 = 32'd6591
; 
32'd180176: dataIn1 = 32'd8885
; 
32'd180177: dataIn1 = 32'd8916
; 
32'd180178: dataIn1 = 32'd8917
; 
32'd180179: dataIn1 = 32'd8918
; 
32'd180180: dataIn1 = 32'd8920
; 
32'd180181: dataIn1 = 32'd5129
; 
32'd180182: dataIn1 = 32'd6591
; 
32'd180183: dataIn1 = 32'd6592
; 
32'd180184: dataIn1 = 32'd7199
; 
32'd180185: dataIn1 = 32'd8916
; 
32'd180186: dataIn1 = 32'd8919
; 
32'd180187: dataIn1 = 32'd5266
; 
32'd180188: dataIn1 = 32'd6590
; 
32'd180189: dataIn1 = 32'd6591
; 
32'd180190: dataIn1 = 32'd8885
; 
32'd180191: dataIn1 = 32'd8918
; 
32'd180192: dataIn1 = 32'd8920
; 
32'd180193: dataIn1 = 32'd5888
; 
32'd180194: dataIn1 = 32'd6164
; 
32'd180195: dataIn1 = 32'd8921
; 
32'd180196: dataIn1 = 32'd8922
; 
32'd180197: dataIn1 = 32'd8923
; 
32'd180198: dataIn1 = 32'd8924
; 
32'd180199: dataIn1 = 32'd8925
; 
32'd180200: dataIn1 = 32'd6164
; 
32'd180201: dataIn1 = 32'd6595
; 
32'd180202: dataIn1 = 32'd8921
; 
32'd180203: dataIn1 = 32'd8922
; 
32'd180204: dataIn1 = 32'd8923
; 
32'd180205: dataIn1 = 32'd9746
; 
32'd180206: dataIn1 = 32'd9767
; 
32'd180207: dataIn1 = 32'd5888
; 
32'd180208: dataIn1 = 32'd6595
; 
32'd180209: dataIn1 = 32'd7054
; 
32'd180210: dataIn1 = 32'd8921
; 
32'd180211: dataIn1 = 32'd8922
; 
32'd180212: dataIn1 = 32'd8923
; 
32'd180213: dataIn1 = 32'd8926
; 
32'd180214: dataIn1 = 32'd5
; 
32'd180215: dataIn1 = 32'd6055
; 
32'd180216: dataIn1 = 32'd6164
; 
32'd180217: dataIn1 = 32'd7256
; 
32'd180218: dataIn1 = 32'd8921
; 
32'd180219: dataIn1 = 32'd8924
; 
32'd180220: dataIn1 = 32'd8925
; 
32'd180221: dataIn1 = 32'd5
; 
32'd180222: dataIn1 = 32'd5826
; 
32'd180223: dataIn1 = 32'd5888
; 
32'd180224: dataIn1 = 32'd7053
; 
32'd180225: dataIn1 = 32'd8921
; 
32'd180226: dataIn1 = 32'd8924
; 
32'd180227: dataIn1 = 32'd8925
; 
32'd180228: dataIn1 = 32'd3985
; 
32'd180229: dataIn1 = 32'd6595
; 
32'd180230: dataIn1 = 32'd7054
; 
32'd180231: dataIn1 = 32'd8923
; 
32'd180232: dataIn1 = 32'd8926
; 
32'd180233: dataIn1 = 32'd9744
; 
32'd180234: dataIn1 = 32'd9768
; 
32'd180235: dataIn1 = 32'd6600
; 
32'd180236: dataIn1 = 32'd6601
; 
32'd180237: dataIn1 = 32'd8927
; 
32'd180238: dataIn1 = 32'd8928
; 
32'd180239: dataIn1 = 32'd8929
; 
32'd180240: dataIn1 = 32'd8930
; 
32'd180241: dataIn1 = 32'd8931
; 
32'd180242: dataIn1 = 32'd6599
; 
32'd180243: dataIn1 = 32'd6601
; 
32'd180244: dataIn1 = 32'd8927
; 
32'd180245: dataIn1 = 32'd8928
; 
32'd180246: dataIn1 = 32'd8929
; 
32'd180247: dataIn1 = 32'd8932
; 
32'd180248: dataIn1 = 32'd8933
; 
32'd180249: dataIn1 = 32'd6599
; 
32'd180250: dataIn1 = 32'd6600
; 
32'd180251: dataIn1 = 32'd8927
; 
32'd180252: dataIn1 = 32'd8928
; 
32'd180253: dataIn1 = 32'd8929
; 
32'd180254: dataIn1 = 32'd8934
; 
32'd180255: dataIn1 = 32'd8935
; 
32'd180256: dataIn1 = 32'd5274
; 
32'd180257: dataIn1 = 32'd6601
; 
32'd180258: dataIn1 = 32'd8927
; 
32'd180259: dataIn1 = 32'd8930
; 
32'd180260: dataIn1 = 32'd8931
; 
32'd180261: dataIn1 = 32'd8943
; 
32'd180262: dataIn1 = 32'd8946
; 
32'd180263: dataIn1 = 32'd5274
; 
32'd180264: dataIn1 = 32'd6600
; 
32'd180265: dataIn1 = 32'd8927
; 
32'd180266: dataIn1 = 32'd8930
; 
32'd180267: dataIn1 = 32'd8931
; 
32'd180268: dataIn1 = 32'd8936
; 
32'd180269: dataIn1 = 32'd8939
; 
32'd180270: dataIn1 = 32'd5275
; 
32'd180271: dataIn1 = 32'd6601
; 
32'd180272: dataIn1 = 32'd8928
; 
32'd180273: dataIn1 = 32'd8932
; 
32'd180274: dataIn1 = 32'd8933
; 
32'd180275: dataIn1 = 32'd8944
; 
32'd180276: dataIn1 = 32'd8947
; 
32'd180277: dataIn1 = 32'd5275
; 
32'd180278: dataIn1 = 32'd6599
; 
32'd180279: dataIn1 = 32'd8928
; 
32'd180280: dataIn1 = 32'd8932
; 
32'd180281: dataIn1 = 32'd8933
; 
32'd180282: dataIn1 = 32'd9278
; 
32'd180283: dataIn1 = 32'd5276
; 
32'd180284: dataIn1 = 32'd6600
; 
32'd180285: dataIn1 = 32'd8929
; 
32'd180286: dataIn1 = 32'd8934
; 
32'd180287: dataIn1 = 32'd8935
; 
32'd180288: dataIn1 = 32'd8938
; 
32'd180289: dataIn1 = 32'd8942
; 
32'd180290: dataIn1 = 32'd5276
; 
32'd180291: dataIn1 = 32'd6599
; 
32'd180292: dataIn1 = 32'd8929
; 
32'd180293: dataIn1 = 32'd8934
; 
32'd180294: dataIn1 = 32'd8935
; 
32'd180295: dataIn1 = 32'd9277
; 
32'd180296: dataIn1 = 32'd6600
; 
32'd180297: dataIn1 = 32'd6603
; 
32'd180298: dataIn1 = 32'd8931
; 
32'd180299: dataIn1 = 32'd8936
; 
32'd180300: dataIn1 = 32'd8937
; 
32'd180301: dataIn1 = 32'd8938
; 
32'd180302: dataIn1 = 32'd8939
; 
32'd180303: dataIn1 = 32'd6602
; 
32'd180304: dataIn1 = 32'd6603
; 
32'd180305: dataIn1 = 32'd8936
; 
32'd180306: dataIn1 = 32'd8937
; 
32'd180307: dataIn1 = 32'd8938
; 
32'd180308: dataIn1 = 32'd8940
; 
32'd180309: dataIn1 = 32'd8941
; 
32'd180310: dataIn1 = 32'd6600
; 
32'd180311: dataIn1 = 32'd6602
; 
32'd180312: dataIn1 = 32'd8934
; 
32'd180313: dataIn1 = 32'd8936
; 
32'd180314: dataIn1 = 32'd8937
; 
32'd180315: dataIn1 = 32'd8938
; 
32'd180316: dataIn1 = 32'd8942
; 
32'd180317: dataIn1 = 32'd5274
; 
32'd180318: dataIn1 = 32'd6603
; 
32'd180319: dataIn1 = 32'd8931
; 
32'd180320: dataIn1 = 32'd8936
; 
32'd180321: dataIn1 = 32'd8939
; 
32'd180322: dataIn1 = 32'd8954
; 
32'd180323: dataIn1 = 32'd8964
; 
32'd180324: dataIn1 = 32'd2703
; 
32'd180325: dataIn1 = 32'd6603
; 
32'd180326: dataIn1 = 32'd7351
; 
32'd180327: dataIn1 = 32'd8937
; 
32'd180328: dataIn1 = 32'd8940
; 
32'd180329: dataIn1 = 32'd8941
; 
32'd180330: dataIn1 = 32'd8965
; 
32'd180331: dataIn1 = 32'd2703
; 
32'd180332: dataIn1 = 32'd6602
; 
32'd180333: dataIn1 = 32'd7316
; 
32'd180334: dataIn1 = 32'd8937
; 
32'd180335: dataIn1 = 32'd8940
; 
32'd180336: dataIn1 = 32'd8941
; 
32'd180337: dataIn1 = 32'd8975
; 
32'd180338: dataIn1 = 32'd5276
; 
32'd180339: dataIn1 = 32'd6602
; 
32'd180340: dataIn1 = 32'd6610
; 
32'd180341: dataIn1 = 32'd8934
; 
32'd180342: dataIn1 = 32'd8938
; 
32'd180343: dataIn1 = 32'd8942
; 
32'd180344: dataIn1 = 32'd6601
; 
32'd180345: dataIn1 = 32'd6605
; 
32'd180346: dataIn1 = 32'd8930
; 
32'd180347: dataIn1 = 32'd8943
; 
32'd180348: dataIn1 = 32'd8944
; 
32'd180349: dataIn1 = 32'd8945
; 
32'd180350: dataIn1 = 32'd8946
; 
32'd180351: dataIn1 = 32'd6601
; 
32'd180352: dataIn1 = 32'd6604
; 
32'd180353: dataIn1 = 32'd8932
; 
32'd180354: dataIn1 = 32'd8943
; 
32'd180355: dataIn1 = 32'd8944
; 
32'd180356: dataIn1 = 32'd8945
; 
32'd180357: dataIn1 = 32'd8947
; 
32'd180358: dataIn1 = 32'd6604
; 
32'd180359: dataIn1 = 32'd6605
; 
32'd180360: dataIn1 = 32'd8943
; 
32'd180361: dataIn1 = 32'd8944
; 
32'd180362: dataIn1 = 32'd8945
; 
32'd180363: dataIn1 = 32'd8948
; 
32'd180364: dataIn1 = 32'd8949
; 
32'd180365: dataIn1 = 32'd5274
; 
32'd180366: dataIn1 = 32'd6605
; 
32'd180367: dataIn1 = 32'd8930
; 
32'd180368: dataIn1 = 32'd8943
; 
32'd180369: dataIn1 = 32'd8946
; 
32'd180370: dataIn1 = 32'd8953
; 
32'd180371: dataIn1 = 32'd8967
; 
32'd180372: dataIn1 = 32'd5275
; 
32'd180373: dataIn1 = 32'd6604
; 
32'd180374: dataIn1 = 32'd8932
; 
32'd180375: dataIn1 = 32'd8944
; 
32'd180376: dataIn1 = 32'd8947
; 
32'd180377: dataIn1 = 32'd8971
; 
32'd180378: dataIn1 = 32'd8974
; 
32'd180379: dataIn1 = 32'd2707
; 
32'd180380: dataIn1 = 32'd6605
; 
32'd180381: dataIn1 = 32'd7466
; 
32'd180382: dataIn1 = 32'd8945
; 
32'd180383: dataIn1 = 32'd8948
; 
32'd180384: dataIn1 = 32'd8949
; 
32'd180385: dataIn1 = 32'd8969
; 
32'd180386: dataIn1 = 32'd2707
; 
32'd180387: dataIn1 = 32'd6604
; 
32'd180388: dataIn1 = 32'd7511
; 
32'd180389: dataIn1 = 32'd8945
; 
32'd180390: dataIn1 = 32'd8948
; 
32'd180391: dataIn1 = 32'd8949
; 
32'd180392: dataIn1 = 32'd8972
; 
32'd180393: dataIn1 = 32'd6607
; 
32'd180394: dataIn1 = 32'd6608
; 
32'd180395: dataIn1 = 32'd8950
; 
32'd180396: dataIn1 = 32'd8951
; 
32'd180397: dataIn1 = 32'd8952
; 
32'd180398: dataIn1 = 32'd8953
; 
32'd180399: dataIn1 = 32'd8954
; 
32'd180400: dataIn1 = 32'd6606
; 
32'd180401: dataIn1 = 32'd6608
; 
32'd180402: dataIn1 = 32'd8950
; 
32'd180403: dataIn1 = 32'd8951
; 
32'd180404: dataIn1 = 32'd8952
; 
32'd180405: dataIn1 = 32'd8955
; 
32'd180406: dataIn1 = 32'd8956
; 
32'd180407: dataIn1 = 32'd6606
; 
32'd180408: dataIn1 = 32'd6607
; 
32'd180409: dataIn1 = 32'd8950
; 
32'd180410: dataIn1 = 32'd8951
; 
32'd180411: dataIn1 = 32'd8952
; 
32'd180412: dataIn1 = 32'd8957
; 
32'd180413: dataIn1 = 32'd8958
; 
32'd180414: dataIn1 = 32'd5274
; 
32'd180415: dataIn1 = 32'd6608
; 
32'd180416: dataIn1 = 32'd8946
; 
32'd180417: dataIn1 = 32'd8950
; 
32'd180418: dataIn1 = 32'd8953
; 
32'd180419: dataIn1 = 32'd8954
; 
32'd180420: dataIn1 = 32'd8967
; 
32'd180421: dataIn1 = 32'd5274
; 
32'd180422: dataIn1 = 32'd6607
; 
32'd180423: dataIn1 = 32'd8939
; 
32'd180424: dataIn1 = 32'd8950
; 
32'd180425: dataIn1 = 32'd8953
; 
32'd180426: dataIn1 = 32'd8954
; 
32'd180427: dataIn1 = 32'd8964
; 
32'd180428: dataIn1 = 32'd5162
; 
32'd180429: dataIn1 = 32'd6608
; 
32'd180430: dataIn1 = 32'd7467
; 
32'd180431: dataIn1 = 32'd8951
; 
32'd180432: dataIn1 = 32'd8955
; 
32'd180433: dataIn1 = 32'd8956
; 
32'd180434: dataIn1 = 32'd8968
; 
32'd180435: dataIn1 = 32'd5162
; 
32'd180436: dataIn1 = 32'd6606
; 
32'd180437: dataIn1 = 32'd7462
; 
32'd180438: dataIn1 = 32'd8951
; 
32'd180439: dataIn1 = 32'd8955
; 
32'd180440: dataIn1 = 32'd8956
; 
32'd180441: dataIn1 = 32'd8960
; 
32'd180442: dataIn1 = 32'd5149
; 
32'd180443: dataIn1 = 32'd6607
; 
32'd180444: dataIn1 = 32'd7350
; 
32'd180445: dataIn1 = 32'd8952
; 
32'd180446: dataIn1 = 32'd8957
; 
32'd180447: dataIn1 = 32'd8958
; 
32'd180448: dataIn1 = 32'd8966
; 
32'd180449: dataIn1 = 32'd5149
; 
32'd180450: dataIn1 = 32'd6606
; 
32'd180451: dataIn1 = 32'd7355
; 
32'd180452: dataIn1 = 32'd8952
; 
32'd180453: dataIn1 = 32'd8957
; 
32'd180454: dataIn1 = 32'd8958
; 
32'd180455: dataIn1 = 32'd8961
; 
32'd180456: dataIn1 = 32'd6188
; 
32'd180457: dataIn1 = 32'd6219
; 
32'd180458: dataIn1 = 32'd8959
; 
32'd180459: dataIn1 = 32'd8960
; 
32'd180460: dataIn1 = 32'd8961
; 
32'd180461: dataIn1 = 32'd8962
; 
32'd180462: dataIn1 = 32'd8963
; 
32'd180463: dataIn1 = 32'd6219
; 
32'd180464: dataIn1 = 32'd6606
; 
32'd180465: dataIn1 = 32'd7462
; 
32'd180466: dataIn1 = 32'd8956
; 
32'd180467: dataIn1 = 32'd8959
; 
32'd180468: dataIn1 = 32'd8960
; 
32'd180469: dataIn1 = 32'd8961
; 
32'd180470: dataIn1 = 32'd6188
; 
32'd180471: dataIn1 = 32'd6606
; 
32'd180472: dataIn1 = 32'd7355
; 
32'd180473: dataIn1 = 32'd8958
; 
32'd180474: dataIn1 = 32'd8959
; 
32'd180475: dataIn1 = 32'd8960
; 
32'd180476: dataIn1 = 32'd8961
; 
32'd180477: dataIn1 = 32'd6
; 
32'd180478: dataIn1 = 32'd6065
; 
32'd180479: dataIn1 = 32'd6219
; 
32'd180480: dataIn1 = 32'd7458
; 
32'd180481: dataIn1 = 32'd8959
; 
32'd180482: dataIn1 = 32'd8962
; 
32'd180483: dataIn1 = 32'd8963
; 
32'd180484: dataIn1 = 32'd6
; 
32'd180485: dataIn1 = 32'd5995
; 
32'd180486: dataIn1 = 32'd6188
; 
32'd180487: dataIn1 = 32'd7354
; 
32'd180488: dataIn1 = 32'd8959
; 
32'd180489: dataIn1 = 32'd8962
; 
32'd180490: dataIn1 = 32'd8963
; 
32'd180491: dataIn1 = 32'd6603
; 
32'd180492: dataIn1 = 32'd6607
; 
32'd180493: dataIn1 = 32'd8939
; 
32'd180494: dataIn1 = 32'd8954
; 
32'd180495: dataIn1 = 32'd8964
; 
32'd180496: dataIn1 = 32'd8965
; 
32'd180497: dataIn1 = 32'd8966
; 
32'd180498: dataIn1 = 32'd6187
; 
32'd180499: dataIn1 = 32'd6603
; 
32'd180500: dataIn1 = 32'd7351
; 
32'd180501: dataIn1 = 32'd8940
; 
32'd180502: dataIn1 = 32'd8964
; 
32'd180503: dataIn1 = 32'd8965
; 
32'd180504: dataIn1 = 32'd8966
; 
32'd180505: dataIn1 = 32'd6187
; 
32'd180506: dataIn1 = 32'd6607
; 
32'd180507: dataIn1 = 32'd7350
; 
32'd180508: dataIn1 = 32'd8957
; 
32'd180509: dataIn1 = 32'd8964
; 
32'd180510: dataIn1 = 32'd8965
; 
32'd180511: dataIn1 = 32'd8966
; 
32'd180512: dataIn1 = 32'd6605
; 
32'd180513: dataIn1 = 32'd6608
; 
32'd180514: dataIn1 = 32'd8946
; 
32'd180515: dataIn1 = 32'd8953
; 
32'd180516: dataIn1 = 32'd8967
; 
32'd180517: dataIn1 = 32'd8968
; 
32'd180518: dataIn1 = 32'd8969
; 
32'd180519: dataIn1 = 32'd6220
; 
32'd180520: dataIn1 = 32'd6608
; 
32'd180521: dataIn1 = 32'd7467
; 
32'd180522: dataIn1 = 32'd8955
; 
32'd180523: dataIn1 = 32'd8967
; 
32'd180524: dataIn1 = 32'd8968
; 
32'd180525: dataIn1 = 32'd8969
; 
32'd180526: dataIn1 = 32'd6220
; 
32'd180527: dataIn1 = 32'd6605
; 
32'd180528: dataIn1 = 32'd7466
; 
32'd180529: dataIn1 = 32'd8948
; 
32'd180530: dataIn1 = 32'd8967
; 
32'd180531: dataIn1 = 32'd8968
; 
32'd180532: dataIn1 = 32'd8969
; 
32'd180533: dataIn1 = 32'd6227
; 
32'd180534: dataIn1 = 32'd6609
; 
32'd180535: dataIn1 = 32'd7510
; 
32'd180536: dataIn1 = 32'd8970
; 
32'd180537: dataIn1 = 32'd8971
; 
32'd180538: dataIn1 = 32'd8972
; 
32'd180539: dataIn1 = 32'd8973
; 
32'd180540: dataIn1 = 32'd6604
; 
32'd180541: dataIn1 = 32'd6609
; 
32'd180542: dataIn1 = 32'd8947
; 
32'd180543: dataIn1 = 32'd8970
; 
32'd180544: dataIn1 = 32'd8971
; 
32'd180545: dataIn1 = 32'd8972
; 
32'd180546: dataIn1 = 32'd8974
; 
32'd180547: dataIn1 = 32'd6227
; 
32'd180548: dataIn1 = 32'd6604
; 
32'd180549: dataIn1 = 32'd7511
; 
32'd180550: dataIn1 = 32'd8949
; 
32'd180551: dataIn1 = 32'd8970
; 
32'd180552: dataIn1 = 32'd8971
; 
32'd180553: dataIn1 = 32'd8972
; 
32'd180554: dataIn1 = 32'd5163
; 
32'd180555: dataIn1 = 32'd6609
; 
32'd180556: dataIn1 = 32'd7510
; 
32'd180557: dataIn1 = 32'd8970
; 
32'd180558: dataIn1 = 32'd8973
; 
32'd180559: dataIn1 = 32'd9280
; 
32'd180560: dataIn1 = 32'd5275
; 
32'd180561: dataIn1 = 32'd6609
; 
32'd180562: dataIn1 = 32'd8947
; 
32'd180563: dataIn1 = 32'd8971
; 
32'd180564: dataIn1 = 32'd8974
; 
32'd180565: dataIn1 = 32'd9279
; 
32'd180566: dataIn1 = 32'd6180
; 
32'd180567: dataIn1 = 32'd6602
; 
32'd180568: dataIn1 = 32'd6610
; 
32'd180569: dataIn1 = 32'd7316
; 
32'd180570: dataIn1 = 32'd8941
; 
32'd180571: dataIn1 = 32'd8975
; 
32'd180572: dataIn1 = 32'd6612
; 
32'd180573: dataIn1 = 32'd6613
; 
32'd180574: dataIn1 = 32'd8976
; 
32'd180575: dataIn1 = 32'd8977
; 
32'd180576: dataIn1 = 32'd8978
; 
32'd180577: dataIn1 = 32'd8979
; 
32'd180578: dataIn1 = 32'd8980
; 
32'd180579: dataIn1 = 32'd6611
; 
32'd180580: dataIn1 = 32'd6613
; 
32'd180581: dataIn1 = 32'd8976
; 
32'd180582: dataIn1 = 32'd8977
; 
32'd180583: dataIn1 = 32'd8978
; 
32'd180584: dataIn1 = 32'd8981
; 
32'd180585: dataIn1 = 32'd8982
; 
32'd180586: dataIn1 = 32'd6611
; 
32'd180587: dataIn1 = 32'd6612
; 
32'd180588: dataIn1 = 32'd8976
; 
32'd180589: dataIn1 = 32'd8977
; 
32'd180590: dataIn1 = 32'd8978
; 
32'd180591: dataIn1 = 32'd8983
; 
32'd180592: dataIn1 = 32'd8984
; 
32'd180593: dataIn1 = 32'd5279
; 
32'd180594: dataIn1 = 32'd6613
; 
32'd180595: dataIn1 = 32'd8976
; 
32'd180596: dataIn1 = 32'd8979
; 
32'd180597: dataIn1 = 32'd8980
; 
32'd180598: dataIn1 = 32'd8992
; 
32'd180599: dataIn1 = 32'd8995
; 
32'd180600: dataIn1 = 32'd5279
; 
32'd180601: dataIn1 = 32'd6612
; 
32'd180602: dataIn1 = 32'd8976
; 
32'd180603: dataIn1 = 32'd8979
; 
32'd180604: dataIn1 = 32'd8980
; 
32'd180605: dataIn1 = 32'd8985
; 
32'd180606: dataIn1 = 32'd8988
; 
32'd180607: dataIn1 = 32'd5280
; 
32'd180608: dataIn1 = 32'd6613
; 
32'd180609: dataIn1 = 32'd8977
; 
32'd180610: dataIn1 = 32'd8981
; 
32'd180611: dataIn1 = 32'd8982
; 
32'd180612: dataIn1 = 32'd8993
; 
32'd180613: dataIn1 = 32'd8996
; 
32'd180614: dataIn1 = 32'd5280
; 
32'd180615: dataIn1 = 32'd6611
; 
32'd180616: dataIn1 = 32'd6787
; 
32'd180617: dataIn1 = 32'd8977
; 
32'd180618: dataIn1 = 32'd8981
; 
32'd180619: dataIn1 = 32'd8982
; 
32'd180620: dataIn1 = 32'd5281
; 
32'd180621: dataIn1 = 32'd6612
; 
32'd180622: dataIn1 = 32'd8978
; 
32'd180623: dataIn1 = 32'd8983
; 
32'd180624: dataIn1 = 32'd8984
; 
32'd180625: dataIn1 = 32'd8987
; 
32'd180626: dataIn1 = 32'd8991
; 
32'd180627: dataIn1 = 32'd5281
; 
32'd180628: dataIn1 = 32'd6611
; 
32'd180629: dataIn1 = 32'd6786
; 
32'd180630: dataIn1 = 32'd8978
; 
32'd180631: dataIn1 = 32'd8983
; 
32'd180632: dataIn1 = 32'd8984
; 
32'd180633: dataIn1 = 32'd6612
; 
32'd180634: dataIn1 = 32'd6615
; 
32'd180635: dataIn1 = 32'd8980
; 
32'd180636: dataIn1 = 32'd8985
; 
32'd180637: dataIn1 = 32'd8986
; 
32'd180638: dataIn1 = 32'd8987
; 
32'd180639: dataIn1 = 32'd8988
; 
32'd180640: dataIn1 = 32'd6614
; 
32'd180641: dataIn1 = 32'd6615
; 
32'd180642: dataIn1 = 32'd8985
; 
32'd180643: dataIn1 = 32'd8986
; 
32'd180644: dataIn1 = 32'd8987
; 
32'd180645: dataIn1 = 32'd8989
; 
32'd180646: dataIn1 = 32'd8990
; 
32'd180647: dataIn1 = 32'd6612
; 
32'd180648: dataIn1 = 32'd6614
; 
32'd180649: dataIn1 = 32'd8983
; 
32'd180650: dataIn1 = 32'd8985
; 
32'd180651: dataIn1 = 32'd8986
; 
32'd180652: dataIn1 = 32'd8987
; 
32'd180653: dataIn1 = 32'd8991
; 
32'd180654: dataIn1 = 32'd5279
; 
32'd180655: dataIn1 = 32'd6615
; 
32'd180656: dataIn1 = 32'd8980
; 
32'd180657: dataIn1 = 32'd8985
; 
32'd180658: dataIn1 = 32'd8988
; 
32'd180659: dataIn1 = 32'd9003
; 
32'd180660: dataIn1 = 32'd9011
; 
32'd180661: dataIn1 = 32'd2708
; 
32'd180662: dataIn1 = 32'd6615
; 
32'd180663: dataIn1 = 32'd7599
; 
32'd180664: dataIn1 = 32'd8986
; 
32'd180665: dataIn1 = 32'd8989
; 
32'd180666: dataIn1 = 32'd8990
; 
32'd180667: dataIn1 = 32'd9012
; 
32'd180668: dataIn1 = 32'd2708
; 
32'd180669: dataIn1 = 32'd6614
; 
32'd180670: dataIn1 = 32'd7554
; 
32'd180671: dataIn1 = 32'd8986
; 
32'd180672: dataIn1 = 32'd8989
; 
32'd180673: dataIn1 = 32'd8990
; 
32'd180674: dataIn1 = 32'd9023
; 
32'd180675: dataIn1 = 32'd5281
; 
32'd180676: dataIn1 = 32'd6614
; 
32'd180677: dataIn1 = 32'd8983
; 
32'd180678: dataIn1 = 32'd8987
; 
32'd180679: dataIn1 = 32'd8991
; 
32'd180680: dataIn1 = 32'd9024
; 
32'd180681: dataIn1 = 32'd9026
; 
32'd180682: dataIn1 = 32'd6613
; 
32'd180683: dataIn1 = 32'd6617
; 
32'd180684: dataIn1 = 32'd8979
; 
32'd180685: dataIn1 = 32'd8992
; 
32'd180686: dataIn1 = 32'd8993
; 
32'd180687: dataIn1 = 32'd8994
; 
32'd180688: dataIn1 = 32'd8995
; 
32'd180689: dataIn1 = 32'd6613
; 
32'd180690: dataIn1 = 32'd6616
; 
32'd180691: dataIn1 = 32'd8981
; 
32'd180692: dataIn1 = 32'd8992
; 
32'd180693: dataIn1 = 32'd8993
; 
32'd180694: dataIn1 = 32'd8994
; 
32'd180695: dataIn1 = 32'd8996
; 
32'd180696: dataIn1 = 32'd6616
; 
32'd180697: dataIn1 = 32'd6617
; 
32'd180698: dataIn1 = 32'd8992
; 
32'd180699: dataIn1 = 32'd8993
; 
32'd180700: dataIn1 = 32'd8994
; 
32'd180701: dataIn1 = 32'd8997
; 
32'd180702: dataIn1 = 32'd8998
; 
32'd180703: dataIn1 = 32'd5279
; 
32'd180704: dataIn1 = 32'd6617
; 
32'd180705: dataIn1 = 32'd8979
; 
32'd180706: dataIn1 = 32'd8992
; 
32'd180707: dataIn1 = 32'd8995
; 
32'd180708: dataIn1 = 32'd9002
; 
32'd180709: dataIn1 = 32'd9014
; 
32'd180710: dataIn1 = 32'd5280
; 
32'd180711: dataIn1 = 32'd6616
; 
32'd180712: dataIn1 = 32'd8981
; 
32'd180713: dataIn1 = 32'd8993
; 
32'd180714: dataIn1 = 32'd8996
; 
32'd180715: dataIn1 = 32'd9018
; 
32'd180716: dataIn1 = 32'd9021
; 
32'd180717: dataIn1 = 32'd2712
; 
32'd180718: dataIn1 = 32'd6617
; 
32'd180719: dataIn1 = 32'd7719
; 
32'd180720: dataIn1 = 32'd8994
; 
32'd180721: dataIn1 = 32'd8997
; 
32'd180722: dataIn1 = 32'd8998
; 
32'd180723: dataIn1 = 32'd9016
; 
32'd180724: dataIn1 = 32'd2712
; 
32'd180725: dataIn1 = 32'd6616
; 
32'd180726: dataIn1 = 32'd7764
; 
32'd180727: dataIn1 = 32'd8994
; 
32'd180728: dataIn1 = 32'd8997
; 
32'd180729: dataIn1 = 32'd8998
; 
32'd180730: dataIn1 = 32'd9019
; 
32'd180731: dataIn1 = 32'd6619
; 
32'd180732: dataIn1 = 32'd6620
; 
32'd180733: dataIn1 = 32'd8999
; 
32'd180734: dataIn1 = 32'd9000
; 
32'd180735: dataIn1 = 32'd9001
; 
32'd180736: dataIn1 = 32'd9002
; 
32'd180737: dataIn1 = 32'd9003
; 
32'd180738: dataIn1 = 32'd6618
; 
32'd180739: dataIn1 = 32'd6620
; 
32'd180740: dataIn1 = 32'd8999
; 
32'd180741: dataIn1 = 32'd9000
; 
32'd180742: dataIn1 = 32'd9001
; 
32'd180743: dataIn1 = 32'd9004
; 
32'd180744: dataIn1 = 32'd9005
; 
32'd180745: dataIn1 = 32'd6618
; 
32'd180746: dataIn1 = 32'd6619
; 
32'd180747: dataIn1 = 32'd8999
; 
32'd180748: dataIn1 = 32'd9000
; 
32'd180749: dataIn1 = 32'd9001
; 
32'd180750: dataIn1 = 32'd9006
; 
32'd180751: dataIn1 = 32'd9007
; 
32'd180752: dataIn1 = 32'd5279
; 
32'd180753: dataIn1 = 32'd6620
; 
32'd180754: dataIn1 = 32'd8995
; 
32'd180755: dataIn1 = 32'd8999
; 
32'd180756: dataIn1 = 32'd9002
; 
32'd180757: dataIn1 = 32'd9003
; 
32'd180758: dataIn1 = 32'd9014
; 
32'd180759: dataIn1 = 32'd5279
; 
32'd180760: dataIn1 = 32'd6619
; 
32'd180761: dataIn1 = 32'd8988
; 
32'd180762: dataIn1 = 32'd8999
; 
32'd180763: dataIn1 = 32'd9002
; 
32'd180764: dataIn1 = 32'd9003
; 
32'd180765: dataIn1 = 32'd9011
; 
32'd180766: dataIn1 = 32'd5181
; 
32'd180767: dataIn1 = 32'd6620
; 
32'd180768: dataIn1 = 32'd7720
; 
32'd180769: dataIn1 = 32'd9000
; 
32'd180770: dataIn1 = 32'd9004
; 
32'd180771: dataIn1 = 32'd9005
; 
32'd180772: dataIn1 = 32'd9015
; 
32'd180773: dataIn1 = 32'd5181
; 
32'd180774: dataIn1 = 32'd6618
; 
32'd180775: dataIn1 = 32'd7715
; 
32'd180776: dataIn1 = 32'd9000
; 
32'd180777: dataIn1 = 32'd9004
; 
32'd180778: dataIn1 = 32'd9005
; 
32'd180779: dataIn1 = 32'd9009
; 
32'd180780: dataIn1 = 32'd5168
; 
32'd180781: dataIn1 = 32'd6619
; 
32'd180782: dataIn1 = 32'd7598
; 
32'd180783: dataIn1 = 32'd9001
; 
32'd180784: dataIn1 = 32'd9006
; 
32'd180785: dataIn1 = 32'd9007
; 
32'd180786: dataIn1 = 32'd9013
; 
32'd180787: dataIn1 = 32'd5168
; 
32'd180788: dataIn1 = 32'd6618
; 
32'd180789: dataIn1 = 32'd7603
; 
32'd180790: dataIn1 = 32'd9001
; 
32'd180791: dataIn1 = 32'd9006
; 
32'd180792: dataIn1 = 32'd9007
; 
32'd180793: dataIn1 = 32'd9010
; 
32'd180794: dataIn1 = 32'd6248
; 
32'd180795: dataIn1 = 32'd6279
; 
32'd180796: dataIn1 = 32'd7605
; 
32'd180797: dataIn1 = 32'd7713
; 
32'd180798: dataIn1 = 32'd9008
; 
32'd180799: dataIn1 = 32'd9009
; 
32'd180800: dataIn1 = 32'd9010
; 
32'd180801: dataIn1 = 32'd6279
; 
32'd180802: dataIn1 = 32'd6618
; 
32'd180803: dataIn1 = 32'd7715
; 
32'd180804: dataIn1 = 32'd9005
; 
32'd180805: dataIn1 = 32'd9008
; 
32'd180806: dataIn1 = 32'd9009
; 
32'd180807: dataIn1 = 32'd9010
; 
32'd180808: dataIn1 = 32'd6248
; 
32'd180809: dataIn1 = 32'd6618
; 
32'd180810: dataIn1 = 32'd7603
; 
32'd180811: dataIn1 = 32'd9007
; 
32'd180812: dataIn1 = 32'd9008
; 
32'd180813: dataIn1 = 32'd9009
; 
32'd180814: dataIn1 = 32'd9010
; 
32'd180815: dataIn1 = 32'd6615
; 
32'd180816: dataIn1 = 32'd6619
; 
32'd180817: dataIn1 = 32'd8988
; 
32'd180818: dataIn1 = 32'd9003
; 
32'd180819: dataIn1 = 32'd9011
; 
32'd180820: dataIn1 = 32'd9012
; 
32'd180821: dataIn1 = 32'd9013
; 
32'd180822: dataIn1 = 32'd6247
; 
32'd180823: dataIn1 = 32'd6615
; 
32'd180824: dataIn1 = 32'd7599
; 
32'd180825: dataIn1 = 32'd8989
; 
32'd180826: dataIn1 = 32'd9011
; 
32'd180827: dataIn1 = 32'd9012
; 
32'd180828: dataIn1 = 32'd9013
; 
32'd180829: dataIn1 = 32'd6247
; 
32'd180830: dataIn1 = 32'd6619
; 
32'd180831: dataIn1 = 32'd7598
; 
32'd180832: dataIn1 = 32'd9006
; 
32'd180833: dataIn1 = 32'd9011
; 
32'd180834: dataIn1 = 32'd9012
; 
32'd180835: dataIn1 = 32'd9013
; 
32'd180836: dataIn1 = 32'd6617
; 
32'd180837: dataIn1 = 32'd6620
; 
32'd180838: dataIn1 = 32'd8995
; 
32'd180839: dataIn1 = 32'd9002
; 
32'd180840: dataIn1 = 32'd9014
; 
32'd180841: dataIn1 = 32'd9015
; 
32'd180842: dataIn1 = 32'd9016
; 
32'd180843: dataIn1 = 32'd6280
; 
32'd180844: dataIn1 = 32'd6620
; 
32'd180845: dataIn1 = 32'd7720
; 
32'd180846: dataIn1 = 32'd9004
; 
32'd180847: dataIn1 = 32'd9014
; 
32'd180848: dataIn1 = 32'd9015
; 
32'd180849: dataIn1 = 32'd9016
; 
32'd180850: dataIn1 = 32'd6280
; 
32'd180851: dataIn1 = 32'd6617
; 
32'd180852: dataIn1 = 32'd7719
; 
32'd180853: dataIn1 = 32'd8997
; 
32'd180854: dataIn1 = 32'd9014
; 
32'd180855: dataIn1 = 32'd9015
; 
32'd180856: dataIn1 = 32'd9016
; 
32'd180857: dataIn1 = 32'd6287
; 
32'd180858: dataIn1 = 32'd6621
; 
32'd180859: dataIn1 = 32'd7763
; 
32'd180860: dataIn1 = 32'd9017
; 
32'd180861: dataIn1 = 32'd9018
; 
32'd180862: dataIn1 = 32'd9019
; 
32'd180863: dataIn1 = 32'd9020
; 
32'd180864: dataIn1 = 32'd6616
; 
32'd180865: dataIn1 = 32'd6621
; 
32'd180866: dataIn1 = 32'd8996
; 
32'd180867: dataIn1 = 32'd9017
; 
32'd180868: dataIn1 = 32'd9018
; 
32'd180869: dataIn1 = 32'd9019
; 
32'd180870: dataIn1 = 32'd9021
; 
32'd180871: dataIn1 = 32'd6287
; 
32'd180872: dataIn1 = 32'd6616
; 
32'd180873: dataIn1 = 32'd7764
; 
32'd180874: dataIn1 = 32'd8998
; 
32'd180875: dataIn1 = 32'd9017
; 
32'd180876: dataIn1 = 32'd9018
; 
32'd180877: dataIn1 = 32'd9019
; 
32'd180878: dataIn1 = 32'd5182
; 
32'd180879: dataIn1 = 32'd6621
; 
32'd180880: dataIn1 = 32'd6789
; 
32'd180881: dataIn1 = 32'd7763
; 
32'd180882: dataIn1 = 32'd9017
; 
32'd180883: dataIn1 = 32'd9020
; 
32'd180884: dataIn1 = 32'd5280
; 
32'd180885: dataIn1 = 32'd6621
; 
32'd180886: dataIn1 = 32'd6788
; 
32'd180887: dataIn1 = 32'd8996
; 
32'd180888: dataIn1 = 32'd9018
; 
32'd180889: dataIn1 = 32'd9021
; 
32'd180890: dataIn1 = 32'd6240
; 
32'd180891: dataIn1 = 32'd6622
; 
32'd180892: dataIn1 = 32'd7555
; 
32'd180893: dataIn1 = 32'd9022
; 
32'd180894: dataIn1 = 32'd9023
; 
32'd180895: dataIn1 = 32'd9024
; 
32'd180896: dataIn1 = 32'd9025
; 
32'd180897: dataIn1 = 32'd6240
; 
32'd180898: dataIn1 = 32'd6614
; 
32'd180899: dataIn1 = 32'd7554
; 
32'd180900: dataIn1 = 32'd8990
; 
32'd180901: dataIn1 = 32'd9022
; 
32'd180902: dataIn1 = 32'd9023
; 
32'd180903: dataIn1 = 32'd9024
; 
32'd180904: dataIn1 = 32'd6614
; 
32'd180905: dataIn1 = 32'd6622
; 
32'd180906: dataIn1 = 32'd8991
; 
32'd180907: dataIn1 = 32'd9022
; 
32'd180908: dataIn1 = 32'd9023
; 
32'd180909: dataIn1 = 32'd9024
; 
32'd180910: dataIn1 = 32'd9026
; 
32'd180911: dataIn1 = 32'd5167
; 
32'd180912: dataIn1 = 32'd6622
; 
32'd180913: dataIn1 = 32'd6791
; 
32'd180914: dataIn1 = 32'd7555
; 
32'd180915: dataIn1 = 32'd9022
; 
32'd180916: dataIn1 = 32'd9025
; 
32'd180917: dataIn1 = 32'd5281
; 
32'd180918: dataIn1 = 32'd6622
; 
32'd180919: dataIn1 = 32'd6790
; 
32'd180920: dataIn1 = 32'd8991
; 
32'd180921: dataIn1 = 32'd9024
; 
32'd180922: dataIn1 = 32'd9026
; 
32'd180923: dataIn1 = 32'd6624
; 
32'd180924: dataIn1 = 32'd6625
; 
32'd180925: dataIn1 = 32'd9027
; 
32'd180926: dataIn1 = 32'd9028
; 
32'd180927: dataIn1 = 32'd9029
; 
32'd180928: dataIn1 = 32'd9030
; 
32'd180929: dataIn1 = 32'd9031
; 
32'd180930: dataIn1 = 32'd6623
; 
32'd180931: dataIn1 = 32'd6625
; 
32'd180932: dataIn1 = 32'd9027
; 
32'd180933: dataIn1 = 32'd9028
; 
32'd180934: dataIn1 = 32'd9029
; 
32'd180935: dataIn1 = 32'd9032
; 
32'd180936: dataIn1 = 32'd9033
; 
32'd180937: dataIn1 = 32'd6623
; 
32'd180938: dataIn1 = 32'd6624
; 
32'd180939: dataIn1 = 32'd9027
; 
32'd180940: dataIn1 = 32'd9028
; 
32'd180941: dataIn1 = 32'd9029
; 
32'd180942: dataIn1 = 32'd9034
; 
32'd180943: dataIn1 = 32'd9035
; 
32'd180944: dataIn1 = 32'd5284
; 
32'd180945: dataIn1 = 32'd6625
; 
32'd180946: dataIn1 = 32'd9027
; 
32'd180947: dataIn1 = 32'd9030
; 
32'd180948: dataIn1 = 32'd9031
; 
32'd180949: dataIn1 = 32'd9044
; 
32'd180950: dataIn1 = 32'd9047
; 
32'd180951: dataIn1 = 32'd5284
; 
32'd180952: dataIn1 = 32'd6624
; 
32'd180953: dataIn1 = 32'd9027
; 
32'd180954: dataIn1 = 32'd9030
; 
32'd180955: dataIn1 = 32'd9031
; 
32'd180956: dataIn1 = 32'd9037
; 
32'd180957: dataIn1 = 32'd9040
; 
32'd180958: dataIn1 = 32'd5285
; 
32'd180959: dataIn1 = 32'd6625
; 
32'd180960: dataIn1 = 32'd9028
; 
32'd180961: dataIn1 = 32'd9032
; 
32'd180962: dataIn1 = 32'd9033
; 
32'd180963: dataIn1 = 32'd9045
; 
32'd180964: dataIn1 = 32'd9048
; 
32'd180965: dataIn1 = 32'd5285
; 
32'd180966: dataIn1 = 32'd6623
; 
32'd180967: dataIn1 = 32'd6627
; 
32'd180968: dataIn1 = 32'd9028
; 
32'd180969: dataIn1 = 32'd9032
; 
32'd180970: dataIn1 = 32'd9033
; 
32'd180971: dataIn1 = 32'd5286
; 
32'd180972: dataIn1 = 32'd6624
; 
32'd180973: dataIn1 = 32'd9029
; 
32'd180974: dataIn1 = 32'd9034
; 
32'd180975: dataIn1 = 32'd9035
; 
32'd180976: dataIn1 = 32'd9039
; 
32'd180977: dataIn1 = 32'd9043
; 
32'd180978: dataIn1 = 32'd5286
; 
32'd180979: dataIn1 = 32'd6623
; 
32'd180980: dataIn1 = 32'd6626
; 
32'd180981: dataIn1 = 32'd9029
; 
32'd180982: dataIn1 = 32'd9034
; 
32'd180983: dataIn1 = 32'd9035
; 
32'd180984: dataIn1 = 32'd2749
; 
32'd180985: dataIn1 = 32'd5288
; 
32'd180986: dataIn1 = 32'd6626
; 
32'd180987: dataIn1 = 32'd6792
; 
32'd180988: dataIn1 = 32'd9036
; 
32'd180989: dataIn1 = 32'd9282
; 
32'd180990: dataIn1 = 32'd6624
; 
32'd180991: dataIn1 = 32'd6629
; 
32'd180992: dataIn1 = 32'd9031
; 
32'd180993: dataIn1 = 32'd9037
; 
32'd180994: dataIn1 = 32'd9038
; 
32'd180995: dataIn1 = 32'd9039
; 
32'd180996: dataIn1 = 32'd9040
; 
32'd180997: dataIn1 = 32'd6628
; 
32'd180998: dataIn1 = 32'd6629
; 
32'd180999: dataIn1 = 32'd9037
; 
32'd181000: dataIn1 = 32'd9038
; 
32'd181001: dataIn1 = 32'd9039
; 
32'd181002: dataIn1 = 32'd9041
; 
32'd181003: dataIn1 = 32'd9042
; 
32'd181004: dataIn1 = 32'd6624
; 
32'd181005: dataIn1 = 32'd6628
; 
32'd181006: dataIn1 = 32'd9034
; 
32'd181007: dataIn1 = 32'd9037
; 
32'd181008: dataIn1 = 32'd9038
; 
32'd181009: dataIn1 = 32'd9039
; 
32'd181010: dataIn1 = 32'd9043
; 
32'd181011: dataIn1 = 32'd5284
; 
32'd181012: dataIn1 = 32'd6629
; 
32'd181013: dataIn1 = 32'd9031
; 
32'd181014: dataIn1 = 32'd9037
; 
32'd181015: dataIn1 = 32'd9040
; 
32'd181016: dataIn1 = 32'd9055
; 
32'd181017: dataIn1 = 32'd9063
; 
32'd181018: dataIn1 = 32'd2713
; 
32'd181019: dataIn1 = 32'd6629
; 
32'd181020: dataIn1 = 32'd7852
; 
32'd181021: dataIn1 = 32'd9038
; 
32'd181022: dataIn1 = 32'd9041
; 
32'd181023: dataIn1 = 32'd9042
; 
32'd181024: dataIn1 = 32'd9064
; 
32'd181025: dataIn1 = 32'd2713
; 
32'd181026: dataIn1 = 32'd6628
; 
32'd181027: dataIn1 = 32'd7807
; 
32'd181028: dataIn1 = 32'd9038
; 
32'd181029: dataIn1 = 32'd9041
; 
32'd181030: dataIn1 = 32'd9042
; 
32'd181031: dataIn1 = 32'd9075
; 
32'd181032: dataIn1 = 32'd5286
; 
32'd181033: dataIn1 = 32'd6628
; 
32'd181034: dataIn1 = 32'd9034
; 
32'd181035: dataIn1 = 32'd9039
; 
32'd181036: dataIn1 = 32'd9043
; 
32'd181037: dataIn1 = 32'd9076
; 
32'd181038: dataIn1 = 32'd9078
; 
32'd181039: dataIn1 = 32'd6625
; 
32'd181040: dataIn1 = 32'd6631
; 
32'd181041: dataIn1 = 32'd9030
; 
32'd181042: dataIn1 = 32'd9044
; 
32'd181043: dataIn1 = 32'd9045
; 
32'd181044: dataIn1 = 32'd9046
; 
32'd181045: dataIn1 = 32'd9047
; 
32'd181046: dataIn1 = 32'd6625
; 
32'd181047: dataIn1 = 32'd6630
; 
32'd181048: dataIn1 = 32'd9032
; 
32'd181049: dataIn1 = 32'd9044
; 
32'd181050: dataIn1 = 32'd9045
; 
32'd181051: dataIn1 = 32'd9046
; 
32'd181052: dataIn1 = 32'd9048
; 
32'd181053: dataIn1 = 32'd6630
; 
32'd181054: dataIn1 = 32'd6631
; 
32'd181055: dataIn1 = 32'd9044
; 
32'd181056: dataIn1 = 32'd9045
; 
32'd181057: dataIn1 = 32'd9046
; 
32'd181058: dataIn1 = 32'd9049
; 
32'd181059: dataIn1 = 32'd9050
; 
32'd181060: dataIn1 = 32'd5284
; 
32'd181061: dataIn1 = 32'd6631
; 
32'd181062: dataIn1 = 32'd9030
; 
32'd181063: dataIn1 = 32'd9044
; 
32'd181064: dataIn1 = 32'd9047
; 
32'd181065: dataIn1 = 32'd9054
; 
32'd181066: dataIn1 = 32'd9066
; 
32'd181067: dataIn1 = 32'd5285
; 
32'd181068: dataIn1 = 32'd6630
; 
32'd181069: dataIn1 = 32'd9032
; 
32'd181070: dataIn1 = 32'd9045
; 
32'd181071: dataIn1 = 32'd9048
; 
32'd181072: dataIn1 = 32'd9070
; 
32'd181073: dataIn1 = 32'd9073
; 
32'd181074: dataIn1 = 32'd2717
; 
32'd181075: dataIn1 = 32'd6631
; 
32'd181076: dataIn1 = 32'd7972
; 
32'd181077: dataIn1 = 32'd9046
; 
32'd181078: dataIn1 = 32'd9049
; 
32'd181079: dataIn1 = 32'd9050
; 
32'd181080: dataIn1 = 32'd9068
; 
32'd181081: dataIn1 = 32'd2717
; 
32'd181082: dataIn1 = 32'd6630
; 
32'd181083: dataIn1 = 32'd8017
; 
32'd181084: dataIn1 = 32'd9046
; 
32'd181085: dataIn1 = 32'd9049
; 
32'd181086: dataIn1 = 32'd9050
; 
32'd181087: dataIn1 = 32'd9071
; 
32'd181088: dataIn1 = 32'd6633
; 
32'd181089: dataIn1 = 32'd6634
; 
32'd181090: dataIn1 = 32'd9051
; 
32'd181091: dataIn1 = 32'd9052
; 
32'd181092: dataIn1 = 32'd9053
; 
32'd181093: dataIn1 = 32'd9054
; 
32'd181094: dataIn1 = 32'd9055
; 
32'd181095: dataIn1 = 32'd6632
; 
32'd181096: dataIn1 = 32'd6634
; 
32'd181097: dataIn1 = 32'd9051
; 
32'd181098: dataIn1 = 32'd9052
; 
32'd181099: dataIn1 = 32'd9053
; 
32'd181100: dataIn1 = 32'd9056
; 
32'd181101: dataIn1 = 32'd9057
; 
32'd181102: dataIn1 = 32'd6632
; 
32'd181103: dataIn1 = 32'd6633
; 
32'd181104: dataIn1 = 32'd9051
; 
32'd181105: dataIn1 = 32'd9052
; 
32'd181106: dataIn1 = 32'd9053
; 
32'd181107: dataIn1 = 32'd9058
; 
32'd181108: dataIn1 = 32'd9059
; 
32'd181109: dataIn1 = 32'd5284
; 
32'd181110: dataIn1 = 32'd6634
; 
32'd181111: dataIn1 = 32'd9047
; 
32'd181112: dataIn1 = 32'd9051
; 
32'd181113: dataIn1 = 32'd9054
; 
32'd181114: dataIn1 = 32'd9055
; 
32'd181115: dataIn1 = 32'd9066
; 
32'd181116: dataIn1 = 32'd5284
; 
32'd181117: dataIn1 = 32'd6633
; 
32'd181118: dataIn1 = 32'd9040
; 
32'd181119: dataIn1 = 32'd9051
; 
32'd181120: dataIn1 = 32'd9054
; 
32'd181121: dataIn1 = 32'd9055
; 
32'd181122: dataIn1 = 32'd9063
; 
32'd181123: dataIn1 = 32'd5200
; 
32'd181124: dataIn1 = 32'd6634
; 
32'd181125: dataIn1 = 32'd7973
; 
32'd181126: dataIn1 = 32'd9052
; 
32'd181127: dataIn1 = 32'd9056
; 
32'd181128: dataIn1 = 32'd9057
; 
32'd181129: dataIn1 = 32'd9067
; 
32'd181130: dataIn1 = 32'd5200
; 
32'd181131: dataIn1 = 32'd6632
; 
32'd181132: dataIn1 = 32'd7968
; 
32'd181133: dataIn1 = 32'd9052
; 
32'd181134: dataIn1 = 32'd9056
; 
32'd181135: dataIn1 = 32'd9057
; 
32'd181136: dataIn1 = 32'd9061
; 
32'd181137: dataIn1 = 32'd5187
; 
32'd181138: dataIn1 = 32'd6633
; 
32'd181139: dataIn1 = 32'd7851
; 
32'd181140: dataIn1 = 32'd9053
; 
32'd181141: dataIn1 = 32'd9058
; 
32'd181142: dataIn1 = 32'd9059
; 
32'd181143: dataIn1 = 32'd9065
; 
32'd181144: dataIn1 = 32'd5187
; 
32'd181145: dataIn1 = 32'd6632
; 
32'd181146: dataIn1 = 32'd7856
; 
32'd181147: dataIn1 = 32'd9053
; 
32'd181148: dataIn1 = 32'd9058
; 
32'd181149: dataIn1 = 32'd9059
; 
32'd181150: dataIn1 = 32'd9062
; 
32'd181151: dataIn1 = 32'd6308
; 
32'd181152: dataIn1 = 32'd6351
; 
32'd181153: dataIn1 = 32'd7858
; 
32'd181154: dataIn1 = 32'd7966
; 
32'd181155: dataIn1 = 32'd9060
; 
32'd181156: dataIn1 = 32'd9061
; 
32'd181157: dataIn1 = 32'd9062
; 
32'd181158: dataIn1 = 32'd6351
; 
32'd181159: dataIn1 = 32'd6632
; 
32'd181160: dataIn1 = 32'd7968
; 
32'd181161: dataIn1 = 32'd9057
; 
32'd181162: dataIn1 = 32'd9060
; 
32'd181163: dataIn1 = 32'd9061
; 
32'd181164: dataIn1 = 32'd9062
; 
32'd181165: dataIn1 = 32'd6308
; 
32'd181166: dataIn1 = 32'd6632
; 
32'd181167: dataIn1 = 32'd7856
; 
32'd181168: dataIn1 = 32'd9059
; 
32'd181169: dataIn1 = 32'd9060
; 
32'd181170: dataIn1 = 32'd9061
; 
32'd181171: dataIn1 = 32'd9062
; 
32'd181172: dataIn1 = 32'd6629
; 
32'd181173: dataIn1 = 32'd6633
; 
32'd181174: dataIn1 = 32'd9040
; 
32'd181175: dataIn1 = 32'd9055
; 
32'd181176: dataIn1 = 32'd9063
; 
32'd181177: dataIn1 = 32'd9064
; 
32'd181178: dataIn1 = 32'd9065
; 
32'd181179: dataIn1 = 32'd6307
; 
32'd181180: dataIn1 = 32'd6629
; 
32'd181181: dataIn1 = 32'd7852
; 
32'd181182: dataIn1 = 32'd9041
; 
32'd181183: dataIn1 = 32'd9063
; 
32'd181184: dataIn1 = 32'd9064
; 
32'd181185: dataIn1 = 32'd9065
; 
32'd181186: dataIn1 = 32'd6307
; 
32'd181187: dataIn1 = 32'd6633
; 
32'd181188: dataIn1 = 32'd7851
; 
32'd181189: dataIn1 = 32'd9058
; 
32'd181190: dataIn1 = 32'd9063
; 
32'd181191: dataIn1 = 32'd9064
; 
32'd181192: dataIn1 = 32'd9065
; 
32'd181193: dataIn1 = 32'd6631
; 
32'd181194: dataIn1 = 32'd6634
; 
32'd181195: dataIn1 = 32'd9047
; 
32'd181196: dataIn1 = 32'd9054
; 
32'd181197: dataIn1 = 32'd9066
; 
32'd181198: dataIn1 = 32'd9067
; 
32'd181199: dataIn1 = 32'd9068
; 
32'd181200: dataIn1 = 32'd6352
; 
32'd181201: dataIn1 = 32'd6634
; 
32'd181202: dataIn1 = 32'd7973
; 
32'd181203: dataIn1 = 32'd9056
; 
32'd181204: dataIn1 = 32'd9066
; 
32'd181205: dataIn1 = 32'd9067
; 
32'd181206: dataIn1 = 32'd9068
; 
32'd181207: dataIn1 = 32'd6352
; 
32'd181208: dataIn1 = 32'd6631
; 
32'd181209: dataIn1 = 32'd7972
; 
32'd181210: dataIn1 = 32'd9049
; 
32'd181211: dataIn1 = 32'd9066
; 
32'd181212: dataIn1 = 32'd9067
; 
32'd181213: dataIn1 = 32'd9068
; 
32'd181214: dataIn1 = 32'd6359
; 
32'd181215: dataIn1 = 32'd6639
; 
32'd181216: dataIn1 = 32'd8016
; 
32'd181217: dataIn1 = 32'd9069
; 
32'd181218: dataIn1 = 32'd9070
; 
32'd181219: dataIn1 = 32'd9071
; 
32'd181220: dataIn1 = 32'd9072
; 
32'd181221: dataIn1 = 32'd6630
; 
32'd181222: dataIn1 = 32'd6639
; 
32'd181223: dataIn1 = 32'd9048
; 
32'd181224: dataIn1 = 32'd9069
; 
32'd181225: dataIn1 = 32'd9070
; 
32'd181226: dataIn1 = 32'd9071
; 
32'd181227: dataIn1 = 32'd9073
; 
32'd181228: dataIn1 = 32'd6359
; 
32'd181229: dataIn1 = 32'd6630
; 
32'd181230: dataIn1 = 32'd8017
; 
32'd181231: dataIn1 = 32'd9050
; 
32'd181232: dataIn1 = 32'd9069
; 
32'd181233: dataIn1 = 32'd9070
; 
32'd181234: dataIn1 = 32'd9071
; 
32'd181235: dataIn1 = 32'd5201
; 
32'd181236: dataIn1 = 32'd6638
; 
32'd181237: dataIn1 = 32'd6639
; 
32'd181238: dataIn1 = 32'd8016
; 
32'd181239: dataIn1 = 32'd9069
; 
32'd181240: dataIn1 = 32'd9072
; 
32'd181241: dataIn1 = 32'd5285
; 
32'd181242: dataIn1 = 32'd6635
; 
32'd181243: dataIn1 = 32'd6639
; 
32'd181244: dataIn1 = 32'd9048
; 
32'd181245: dataIn1 = 32'd9070
; 
32'd181246: dataIn1 = 32'd9073
; 
32'd181247: dataIn1 = 32'd6300
; 
32'd181248: dataIn1 = 32'd6640
; 
32'd181249: dataIn1 = 32'd7808
; 
32'd181250: dataIn1 = 32'd9074
; 
32'd181251: dataIn1 = 32'd9075
; 
32'd181252: dataIn1 = 32'd9076
; 
32'd181253: dataIn1 = 32'd9077
; 
32'd181254: dataIn1 = 32'd6300
; 
32'd181255: dataIn1 = 32'd6628
; 
32'd181256: dataIn1 = 32'd7807
; 
32'd181257: dataIn1 = 32'd9042
; 
32'd181258: dataIn1 = 32'd9074
; 
32'd181259: dataIn1 = 32'd9075
; 
32'd181260: dataIn1 = 32'd9076
; 
32'd181261: dataIn1 = 32'd6628
; 
32'd181262: dataIn1 = 32'd6640
; 
32'd181263: dataIn1 = 32'd9043
; 
32'd181264: dataIn1 = 32'd9074
; 
32'd181265: dataIn1 = 32'd9075
; 
32'd181266: dataIn1 = 32'd9076
; 
32'd181267: dataIn1 = 32'd9078
; 
32'd181268: dataIn1 = 32'd5186
; 
32'd181269: dataIn1 = 32'd6640
; 
32'd181270: dataIn1 = 32'd6793
; 
32'd181271: dataIn1 = 32'd7808
; 
32'd181272: dataIn1 = 32'd9074
; 
32'd181273: dataIn1 = 32'd9077
; 
32'd181274: dataIn1 = 32'd5286
; 
32'd181275: dataIn1 = 32'd6640
; 
32'd181276: dataIn1 = 32'd6792
; 
32'd181277: dataIn1 = 32'd9043
; 
32'd181278: dataIn1 = 32'd9076
; 
32'd181279: dataIn1 = 32'd9078
; 
32'd181280: dataIn1 = 32'd6642
; 
32'd181281: dataIn1 = 32'd6643
; 
32'd181282: dataIn1 = 32'd9079
; 
32'd181283: dataIn1 = 32'd9080
; 
32'd181284: dataIn1 = 32'd9081
; 
32'd181285: dataIn1 = 32'd9082
; 
32'd181286: dataIn1 = 32'd9083
; 
32'd181287: dataIn1 = 32'd6641
; 
32'd181288: dataIn1 = 32'd6643
; 
32'd181289: dataIn1 = 32'd9079
; 
32'd181290: dataIn1 = 32'd9080
; 
32'd181291: dataIn1 = 32'd9081
; 
32'd181292: dataIn1 = 32'd9084
; 
32'd181293: dataIn1 = 32'd9085
; 
32'd181294: dataIn1 = 32'd6641
; 
32'd181295: dataIn1 = 32'd6642
; 
32'd181296: dataIn1 = 32'd9079
; 
32'd181297: dataIn1 = 32'd9080
; 
32'd181298: dataIn1 = 32'd9081
; 
32'd181299: dataIn1 = 32'd9086
; 
32'd181300: dataIn1 = 32'd9087
; 
32'd181301: dataIn1 = 32'd5289
; 
32'd181302: dataIn1 = 32'd6643
; 
32'd181303: dataIn1 = 32'd9079
; 
32'd181304: dataIn1 = 32'd9082
; 
32'd181305: dataIn1 = 32'd9083
; 
32'd181306: dataIn1 = 32'd9095
; 
32'd181307: dataIn1 = 32'd9098
; 
32'd181308: dataIn1 = 32'd5289
; 
32'd181309: dataIn1 = 32'd6642
; 
32'd181310: dataIn1 = 32'd9079
; 
32'd181311: dataIn1 = 32'd9082
; 
32'd181312: dataIn1 = 32'd9083
; 
32'd181313: dataIn1 = 32'd9088
; 
32'd181314: dataIn1 = 32'd9091
; 
32'd181315: dataIn1 = 32'd5290
; 
32'd181316: dataIn1 = 32'd6643
; 
32'd181317: dataIn1 = 32'd9080
; 
32'd181318: dataIn1 = 32'd9084
; 
32'd181319: dataIn1 = 32'd9085
; 
32'd181320: dataIn1 = 32'd9096
; 
32'd181321: dataIn1 = 32'd9099
; 
32'd181322: dataIn1 = 32'd5290
; 
32'd181323: dataIn1 = 32'd6641
; 
32'd181324: dataIn1 = 32'd6645
; 
32'd181325: dataIn1 = 32'd9080
; 
32'd181326: dataIn1 = 32'd9084
; 
32'd181327: dataIn1 = 32'd9085
; 
32'd181328: dataIn1 = 32'd5291
; 
32'd181329: dataIn1 = 32'd6642
; 
32'd181330: dataIn1 = 32'd9081
; 
32'd181331: dataIn1 = 32'd9086
; 
32'd181332: dataIn1 = 32'd9087
; 
32'd181333: dataIn1 = 32'd9090
; 
32'd181334: dataIn1 = 32'd9094
; 
32'd181335: dataIn1 = 32'd5291
; 
32'd181336: dataIn1 = 32'd6641
; 
32'd181337: dataIn1 = 32'd6644
; 
32'd181338: dataIn1 = 32'd9081
; 
32'd181339: dataIn1 = 32'd9086
; 
32'd181340: dataIn1 = 32'd9087
; 
32'd181341: dataIn1 = 32'd6642
; 
32'd181342: dataIn1 = 32'd6647
; 
32'd181343: dataIn1 = 32'd9083
; 
32'd181344: dataIn1 = 32'd9088
; 
32'd181345: dataIn1 = 32'd9089
; 
32'd181346: dataIn1 = 32'd9090
; 
32'd181347: dataIn1 = 32'd9091
; 
32'd181348: dataIn1 = 32'd6646
; 
32'd181349: dataIn1 = 32'd6647
; 
32'd181350: dataIn1 = 32'd9088
; 
32'd181351: dataIn1 = 32'd9089
; 
32'd181352: dataIn1 = 32'd9090
; 
32'd181353: dataIn1 = 32'd9092
; 
32'd181354: dataIn1 = 32'd9093
; 
32'd181355: dataIn1 = 32'd6642
; 
32'd181356: dataIn1 = 32'd6646
; 
32'd181357: dataIn1 = 32'd9086
; 
32'd181358: dataIn1 = 32'd9088
; 
32'd181359: dataIn1 = 32'd9089
; 
32'd181360: dataIn1 = 32'd9090
; 
32'd181361: dataIn1 = 32'd9094
; 
32'd181362: dataIn1 = 32'd5289
; 
32'd181363: dataIn1 = 32'd6647
; 
32'd181364: dataIn1 = 32'd9083
; 
32'd181365: dataIn1 = 32'd9088
; 
32'd181366: dataIn1 = 32'd9091
; 
32'd181367: dataIn1 = 32'd9106
; 
32'd181368: dataIn1 = 32'd9114
; 
32'd181369: dataIn1 = 32'd2718
; 
32'd181370: dataIn1 = 32'd6647
; 
32'd181371: dataIn1 = 32'd8105
; 
32'd181372: dataIn1 = 32'd9089
; 
32'd181373: dataIn1 = 32'd9092
; 
32'd181374: dataIn1 = 32'd9093
; 
32'd181375: dataIn1 = 32'd9115
; 
32'd181376: dataIn1 = 32'd2718
; 
32'd181377: dataIn1 = 32'd6646
; 
32'd181378: dataIn1 = 32'd8060
; 
32'd181379: dataIn1 = 32'd9089
; 
32'd181380: dataIn1 = 32'd9092
; 
32'd181381: dataIn1 = 32'd9093
; 
32'd181382: dataIn1 = 32'd9126
; 
32'd181383: dataIn1 = 32'd5291
; 
32'd181384: dataIn1 = 32'd6646
; 
32'd181385: dataIn1 = 32'd9086
; 
32'd181386: dataIn1 = 32'd9090
; 
32'd181387: dataIn1 = 32'd9094
; 
32'd181388: dataIn1 = 32'd9127
; 
32'd181389: dataIn1 = 32'd9129
; 
32'd181390: dataIn1 = 32'd6643
; 
32'd181391: dataIn1 = 32'd6649
; 
32'd181392: dataIn1 = 32'd9082
; 
32'd181393: dataIn1 = 32'd9095
; 
32'd181394: dataIn1 = 32'd9096
; 
32'd181395: dataIn1 = 32'd9097
; 
32'd181396: dataIn1 = 32'd9098
; 
32'd181397: dataIn1 = 32'd6643
; 
32'd181398: dataIn1 = 32'd6648
; 
32'd181399: dataIn1 = 32'd9084
; 
32'd181400: dataIn1 = 32'd9095
; 
32'd181401: dataIn1 = 32'd9096
; 
32'd181402: dataIn1 = 32'd9097
; 
32'd181403: dataIn1 = 32'd9099
; 
32'd181404: dataIn1 = 32'd6648
; 
32'd181405: dataIn1 = 32'd6649
; 
32'd181406: dataIn1 = 32'd9095
; 
32'd181407: dataIn1 = 32'd9096
; 
32'd181408: dataIn1 = 32'd9097
; 
32'd181409: dataIn1 = 32'd9100
; 
32'd181410: dataIn1 = 32'd9101
; 
32'd181411: dataIn1 = 32'd5289
; 
32'd181412: dataIn1 = 32'd6649
; 
32'd181413: dataIn1 = 32'd9082
; 
32'd181414: dataIn1 = 32'd9095
; 
32'd181415: dataIn1 = 32'd9098
; 
32'd181416: dataIn1 = 32'd9105
; 
32'd181417: dataIn1 = 32'd9117
; 
32'd181418: dataIn1 = 32'd5290
; 
32'd181419: dataIn1 = 32'd6648
; 
32'd181420: dataIn1 = 32'd9084
; 
32'd181421: dataIn1 = 32'd9096
; 
32'd181422: dataIn1 = 32'd9099
; 
32'd181423: dataIn1 = 32'd9121
; 
32'd181424: dataIn1 = 32'd9124
; 
32'd181425: dataIn1 = 32'd2722
; 
32'd181426: dataIn1 = 32'd6649
; 
32'd181427: dataIn1 = 32'd8225
; 
32'd181428: dataIn1 = 32'd9097
; 
32'd181429: dataIn1 = 32'd9100
; 
32'd181430: dataIn1 = 32'd9101
; 
32'd181431: dataIn1 = 32'd9119
; 
32'd181432: dataIn1 = 32'd2722
; 
32'd181433: dataIn1 = 32'd6648
; 
32'd181434: dataIn1 = 32'd8270
; 
32'd181435: dataIn1 = 32'd9097
; 
32'd181436: dataIn1 = 32'd9100
; 
32'd181437: dataIn1 = 32'd9101
; 
32'd181438: dataIn1 = 32'd9122
; 
32'd181439: dataIn1 = 32'd6651
; 
32'd181440: dataIn1 = 32'd6652
; 
32'd181441: dataIn1 = 32'd9102
; 
32'd181442: dataIn1 = 32'd9103
; 
32'd181443: dataIn1 = 32'd9104
; 
32'd181444: dataIn1 = 32'd9105
; 
32'd181445: dataIn1 = 32'd9106
; 
32'd181446: dataIn1 = 32'd6650
; 
32'd181447: dataIn1 = 32'd6652
; 
32'd181448: dataIn1 = 32'd9102
; 
32'd181449: dataIn1 = 32'd9103
; 
32'd181450: dataIn1 = 32'd9104
; 
32'd181451: dataIn1 = 32'd9107
; 
32'd181452: dataIn1 = 32'd9108
; 
32'd181453: dataIn1 = 32'd6650
; 
32'd181454: dataIn1 = 32'd6651
; 
32'd181455: dataIn1 = 32'd9102
; 
32'd181456: dataIn1 = 32'd9103
; 
32'd181457: dataIn1 = 32'd9104
; 
32'd181458: dataIn1 = 32'd9109
; 
32'd181459: dataIn1 = 32'd9110
; 
32'd181460: dataIn1 = 32'd5289
; 
32'd181461: dataIn1 = 32'd6652
; 
32'd181462: dataIn1 = 32'd9098
; 
32'd181463: dataIn1 = 32'd9102
; 
32'd181464: dataIn1 = 32'd9105
; 
32'd181465: dataIn1 = 32'd9106
; 
32'd181466: dataIn1 = 32'd9117
; 
32'd181467: dataIn1 = 32'd5289
; 
32'd181468: dataIn1 = 32'd6651
; 
32'd181469: dataIn1 = 32'd9091
; 
32'd181470: dataIn1 = 32'd9102
; 
32'd181471: dataIn1 = 32'd9105
; 
32'd181472: dataIn1 = 32'd9106
; 
32'd181473: dataIn1 = 32'd9114
; 
32'd181474: dataIn1 = 32'd5219
; 
32'd181475: dataIn1 = 32'd6652
; 
32'd181476: dataIn1 = 32'd8226
; 
32'd181477: dataIn1 = 32'd9103
; 
32'd181478: dataIn1 = 32'd9107
; 
32'd181479: dataIn1 = 32'd9108
; 
32'd181480: dataIn1 = 32'd9118
; 
32'd181481: dataIn1 = 32'd5219
; 
32'd181482: dataIn1 = 32'd6650
; 
32'd181483: dataIn1 = 32'd8221
; 
32'd181484: dataIn1 = 32'd9103
; 
32'd181485: dataIn1 = 32'd9107
; 
32'd181486: dataIn1 = 32'd9108
; 
32'd181487: dataIn1 = 32'd9112
; 
32'd181488: dataIn1 = 32'd5206
; 
32'd181489: dataIn1 = 32'd6651
; 
32'd181490: dataIn1 = 32'd8104
; 
32'd181491: dataIn1 = 32'd9104
; 
32'd181492: dataIn1 = 32'd9109
; 
32'd181493: dataIn1 = 32'd9110
; 
32'd181494: dataIn1 = 32'd9116
; 
32'd181495: dataIn1 = 32'd5206
; 
32'd181496: dataIn1 = 32'd6650
; 
32'd181497: dataIn1 = 32'd8109
; 
32'd181498: dataIn1 = 32'd9104
; 
32'd181499: dataIn1 = 32'd9109
; 
32'd181500: dataIn1 = 32'd9110
; 
32'd181501: dataIn1 = 32'd9113
; 
32'd181502: dataIn1 = 32'd6382
; 
32'd181503: dataIn1 = 32'd6422
; 
32'd181504: dataIn1 = 32'd8111
; 
32'd181505: dataIn1 = 32'd8219
; 
32'd181506: dataIn1 = 32'd9111
; 
32'd181507: dataIn1 = 32'd9112
; 
32'd181508: dataIn1 = 32'd9113
; 
32'd181509: dataIn1 = 32'd6422
; 
32'd181510: dataIn1 = 32'd6650
; 
32'd181511: dataIn1 = 32'd8221
; 
32'd181512: dataIn1 = 32'd9108
; 
32'd181513: dataIn1 = 32'd9111
; 
32'd181514: dataIn1 = 32'd9112
; 
32'd181515: dataIn1 = 32'd9113
; 
32'd181516: dataIn1 = 32'd6382
; 
32'd181517: dataIn1 = 32'd6650
; 
32'd181518: dataIn1 = 32'd8109
; 
32'd181519: dataIn1 = 32'd9110
; 
32'd181520: dataIn1 = 32'd9111
; 
32'd181521: dataIn1 = 32'd9112
; 
32'd181522: dataIn1 = 32'd9113
; 
32'd181523: dataIn1 = 32'd6647
; 
32'd181524: dataIn1 = 32'd6651
; 
32'd181525: dataIn1 = 32'd9091
; 
32'd181526: dataIn1 = 32'd9106
; 
32'd181527: dataIn1 = 32'd9114
; 
32'd181528: dataIn1 = 32'd9115
; 
32'd181529: dataIn1 = 32'd9116
; 
32'd181530: dataIn1 = 32'd6381
; 
32'd181531: dataIn1 = 32'd6647
; 
32'd181532: dataIn1 = 32'd8105
; 
32'd181533: dataIn1 = 32'd9092
; 
32'd181534: dataIn1 = 32'd9114
; 
32'd181535: dataIn1 = 32'd9115
; 
32'd181536: dataIn1 = 32'd9116
; 
32'd181537: dataIn1 = 32'd6381
; 
32'd181538: dataIn1 = 32'd6651
; 
32'd181539: dataIn1 = 32'd8104
; 
32'd181540: dataIn1 = 32'd9109
; 
32'd181541: dataIn1 = 32'd9114
; 
32'd181542: dataIn1 = 32'd9115
; 
32'd181543: dataIn1 = 32'd9116
; 
32'd181544: dataIn1 = 32'd6649
; 
32'd181545: dataIn1 = 32'd6652
; 
32'd181546: dataIn1 = 32'd9098
; 
32'd181547: dataIn1 = 32'd9105
; 
32'd181548: dataIn1 = 32'd9117
; 
32'd181549: dataIn1 = 32'd9118
; 
32'd181550: dataIn1 = 32'd9119
; 
32'd181551: dataIn1 = 32'd6423
; 
32'd181552: dataIn1 = 32'd6652
; 
32'd181553: dataIn1 = 32'd8226
; 
32'd181554: dataIn1 = 32'd9107
; 
32'd181555: dataIn1 = 32'd9117
; 
32'd181556: dataIn1 = 32'd9118
; 
32'd181557: dataIn1 = 32'd9119
; 
32'd181558: dataIn1 = 32'd6423
; 
32'd181559: dataIn1 = 32'd6649
; 
32'd181560: dataIn1 = 32'd8225
; 
32'd181561: dataIn1 = 32'd9100
; 
32'd181562: dataIn1 = 32'd9117
; 
32'd181563: dataIn1 = 32'd9118
; 
32'd181564: dataIn1 = 32'd9119
; 
32'd181565: dataIn1 = 32'd6430
; 
32'd181566: dataIn1 = 32'd6655
; 
32'd181567: dataIn1 = 32'd8269
; 
32'd181568: dataIn1 = 32'd9120
; 
32'd181569: dataIn1 = 32'd9121
; 
32'd181570: dataIn1 = 32'd9122
; 
32'd181571: dataIn1 = 32'd9123
; 
32'd181572: dataIn1 = 32'd6648
; 
32'd181573: dataIn1 = 32'd6655
; 
32'd181574: dataIn1 = 32'd9099
; 
32'd181575: dataIn1 = 32'd9120
; 
32'd181576: dataIn1 = 32'd9121
; 
32'd181577: dataIn1 = 32'd9122
; 
32'd181578: dataIn1 = 32'd9124
; 
32'd181579: dataIn1 = 32'd6430
; 
32'd181580: dataIn1 = 32'd6648
; 
32'd181581: dataIn1 = 32'd8270
; 
32'd181582: dataIn1 = 32'd9101
; 
32'd181583: dataIn1 = 32'd9120
; 
32'd181584: dataIn1 = 32'd9121
; 
32'd181585: dataIn1 = 32'd9122
; 
32'd181586: dataIn1 = 32'd5220
; 
32'd181587: dataIn1 = 32'd6655
; 
32'd181588: dataIn1 = 32'd6725
; 
32'd181589: dataIn1 = 32'd8269
; 
32'd181590: dataIn1 = 32'd9120
; 
32'd181591: dataIn1 = 32'd9123
; 
32'd181592: dataIn1 = 32'd5290
; 
32'd181593: dataIn1 = 32'd6653
; 
32'd181594: dataIn1 = 32'd6655
; 
32'd181595: dataIn1 = 32'd9099
; 
32'd181596: dataIn1 = 32'd9121
; 
32'd181597: dataIn1 = 32'd9124
; 
32'd181598: dataIn1 = 32'd6374
; 
32'd181599: dataIn1 = 32'd6658
; 
32'd181600: dataIn1 = 32'd8061
; 
32'd181601: dataIn1 = 32'd9125
; 
32'd181602: dataIn1 = 32'd9126
; 
32'd181603: dataIn1 = 32'd9127
; 
32'd181604: dataIn1 = 32'd9128
; 
32'd181605: dataIn1 = 32'd6374
; 
32'd181606: dataIn1 = 32'd6646
; 
32'd181607: dataIn1 = 32'd8060
; 
32'd181608: dataIn1 = 32'd9093
; 
32'd181609: dataIn1 = 32'd9125
; 
32'd181610: dataIn1 = 32'd9126
; 
32'd181611: dataIn1 = 32'd9127
; 
32'd181612: dataIn1 = 32'd6646
; 
32'd181613: dataIn1 = 32'd6658
; 
32'd181614: dataIn1 = 32'd9094
; 
32'd181615: dataIn1 = 32'd9125
; 
32'd181616: dataIn1 = 32'd9126
; 
32'd181617: dataIn1 = 32'd9127
; 
32'd181618: dataIn1 = 32'd9129
; 
32'd181619: dataIn1 = 32'd5205
; 
32'd181620: dataIn1 = 32'd6658
; 
32'd181621: dataIn1 = 32'd6660
; 
32'd181622: dataIn1 = 32'd8061
; 
32'd181623: dataIn1 = 32'd9125
; 
32'd181624: dataIn1 = 32'd9128
; 
32'd181625: dataIn1 = 32'd5291
; 
32'd181626: dataIn1 = 32'd6656
; 
32'd181627: dataIn1 = 32'd6658
; 
32'd181628: dataIn1 = 32'd9094
; 
32'd181629: dataIn1 = 32'd9127
; 
32'd181630: dataIn1 = 32'd9129
; 
32'd181631: dataIn1 = 32'd6662
; 
32'd181632: dataIn1 = 32'd6663
; 
32'd181633: dataIn1 = 32'd9130
; 
32'd181634: dataIn1 = 32'd9131
; 
32'd181635: dataIn1 = 32'd9132
; 
32'd181636: dataIn1 = 32'd9133
; 
32'd181637: dataIn1 = 32'd9134
; 
32'd181638: dataIn1 = 32'd6661
; 
32'd181639: dataIn1 = 32'd6663
; 
32'd181640: dataIn1 = 32'd9130
; 
32'd181641: dataIn1 = 32'd9131
; 
32'd181642: dataIn1 = 32'd9132
; 
32'd181643: dataIn1 = 32'd9135
; 
32'd181644: dataIn1 = 32'd9136
; 
32'd181645: dataIn1 = 32'd6661
; 
32'd181646: dataIn1 = 32'd6662
; 
32'd181647: dataIn1 = 32'd9130
; 
32'd181648: dataIn1 = 32'd9131
; 
32'd181649: dataIn1 = 32'd9132
; 
32'd181650: dataIn1 = 32'd9137
; 
32'd181651: dataIn1 = 32'd9138
; 
32'd181652: dataIn1 = 32'd5294
; 
32'd181653: dataIn1 = 32'd6663
; 
32'd181654: dataIn1 = 32'd9130
; 
32'd181655: dataIn1 = 32'd9133
; 
32'd181656: dataIn1 = 32'd9134
; 
32'd181657: dataIn1 = 32'd9147
; 
32'd181658: dataIn1 = 32'd9150
; 
32'd181659: dataIn1 = 32'd5294
; 
32'd181660: dataIn1 = 32'd6662
; 
32'd181661: dataIn1 = 32'd9130
; 
32'd181662: dataIn1 = 32'd9133
; 
32'd181663: dataIn1 = 32'd9134
; 
32'd181664: dataIn1 = 32'd9140
; 
32'd181665: dataIn1 = 32'd9143
; 
32'd181666: dataIn1 = 32'd5295
; 
32'd181667: dataIn1 = 32'd6663
; 
32'd181668: dataIn1 = 32'd9131
; 
32'd181669: dataIn1 = 32'd9135
; 
32'd181670: dataIn1 = 32'd9136
; 
32'd181671: dataIn1 = 32'd9148
; 
32'd181672: dataIn1 = 32'd9151
; 
32'd181673: dataIn1 = 32'd5295
; 
32'd181674: dataIn1 = 32'd6661
; 
32'd181675: dataIn1 = 32'd6665
; 
32'd181676: dataIn1 = 32'd9131
; 
32'd181677: dataIn1 = 32'd9135
; 
32'd181678: dataIn1 = 32'd9136
; 
32'd181679: dataIn1 = 32'd5296
; 
32'd181680: dataIn1 = 32'd6662
; 
32'd181681: dataIn1 = 32'd9132
; 
32'd181682: dataIn1 = 32'd9137
; 
32'd181683: dataIn1 = 32'd9138
; 
32'd181684: dataIn1 = 32'd9142
; 
32'd181685: dataIn1 = 32'd9146
; 
32'd181686: dataIn1 = 32'd5296
; 
32'd181687: dataIn1 = 32'd6661
; 
32'd181688: dataIn1 = 32'd6664
; 
32'd181689: dataIn1 = 32'd9132
; 
32'd181690: dataIn1 = 32'd9137
; 
32'd181691: dataIn1 = 32'd9138
; 
32'd181692: dataIn1 = 32'd2751
; 
32'd181693: dataIn1 = 32'd5297
; 
32'd181694: dataIn1 = 32'd6665
; 
32'd181695: dataIn1 = 32'd6794
; 
32'd181696: dataIn1 = 32'd9139
; 
32'd181697: dataIn1 = 32'd9284
; 
32'd181698: dataIn1 = 32'd6662
; 
32'd181699: dataIn1 = 32'd6667
; 
32'd181700: dataIn1 = 32'd9134
; 
32'd181701: dataIn1 = 32'd9140
; 
32'd181702: dataIn1 = 32'd9141
; 
32'd181703: dataIn1 = 32'd9142
; 
32'd181704: dataIn1 = 32'd9143
; 
32'd181705: dataIn1 = 32'd6666
; 
32'd181706: dataIn1 = 32'd6667
; 
32'd181707: dataIn1 = 32'd9140
; 
32'd181708: dataIn1 = 32'd9141
; 
32'd181709: dataIn1 = 32'd9142
; 
32'd181710: dataIn1 = 32'd9144
; 
32'd181711: dataIn1 = 32'd9145
; 
32'd181712: dataIn1 = 32'd6662
; 
32'd181713: dataIn1 = 32'd6666
; 
32'd181714: dataIn1 = 32'd9137
; 
32'd181715: dataIn1 = 32'd9140
; 
32'd181716: dataIn1 = 32'd9141
; 
32'd181717: dataIn1 = 32'd9142
; 
32'd181718: dataIn1 = 32'd9146
; 
32'd181719: dataIn1 = 32'd5294
; 
32'd181720: dataIn1 = 32'd6667
; 
32'd181721: dataIn1 = 32'd9134
; 
32'd181722: dataIn1 = 32'd9140
; 
32'd181723: dataIn1 = 32'd9143
; 
32'd181724: dataIn1 = 32'd9158
; 
32'd181725: dataIn1 = 32'd9166
; 
32'd181726: dataIn1 = 32'd2723
; 
32'd181727: dataIn1 = 32'd6667
; 
32'd181728: dataIn1 = 32'd8357
; 
32'd181729: dataIn1 = 32'd9141
; 
32'd181730: dataIn1 = 32'd9144
; 
32'd181731: dataIn1 = 32'd9145
; 
32'd181732: dataIn1 = 32'd9167
; 
32'd181733: dataIn1 = 32'd2723
; 
32'd181734: dataIn1 = 32'd6666
; 
32'd181735: dataIn1 = 32'd8313
; 
32'd181736: dataIn1 = 32'd9141
; 
32'd181737: dataIn1 = 32'd9144
; 
32'd181738: dataIn1 = 32'd9145
; 
32'd181739: dataIn1 = 32'd9178
; 
32'd181740: dataIn1 = 32'd5296
; 
32'd181741: dataIn1 = 32'd6666
; 
32'd181742: dataIn1 = 32'd9137
; 
32'd181743: dataIn1 = 32'd9142
; 
32'd181744: dataIn1 = 32'd9146
; 
32'd181745: dataIn1 = 32'd9179
; 
32'd181746: dataIn1 = 32'd9180
; 
32'd181747: dataIn1 = 32'd6663
; 
32'd181748: dataIn1 = 32'd6669
; 
32'd181749: dataIn1 = 32'd9133
; 
32'd181750: dataIn1 = 32'd9147
; 
32'd181751: dataIn1 = 32'd9148
; 
32'd181752: dataIn1 = 32'd9149
; 
32'd181753: dataIn1 = 32'd9150
; 
32'd181754: dataIn1 = 32'd6663
; 
32'd181755: dataIn1 = 32'd6668
; 
32'd181756: dataIn1 = 32'd9135
; 
32'd181757: dataIn1 = 32'd9147
; 
32'd181758: dataIn1 = 32'd9148
; 
32'd181759: dataIn1 = 32'd9149
; 
32'd181760: dataIn1 = 32'd9151
; 
32'd181761: dataIn1 = 32'd6668
; 
32'd181762: dataIn1 = 32'd6669
; 
32'd181763: dataIn1 = 32'd9147
; 
32'd181764: dataIn1 = 32'd9148
; 
32'd181765: dataIn1 = 32'd9149
; 
32'd181766: dataIn1 = 32'd9152
; 
32'd181767: dataIn1 = 32'd9153
; 
32'd181768: dataIn1 = 32'd5294
; 
32'd181769: dataIn1 = 32'd6669
; 
32'd181770: dataIn1 = 32'd9133
; 
32'd181771: dataIn1 = 32'd9147
; 
32'd181772: dataIn1 = 32'd9150
; 
32'd181773: dataIn1 = 32'd9157
; 
32'd181774: dataIn1 = 32'd9169
; 
32'd181775: dataIn1 = 32'd5295
; 
32'd181776: dataIn1 = 32'd6668
; 
32'd181777: dataIn1 = 32'd9135
; 
32'd181778: dataIn1 = 32'd9148
; 
32'd181779: dataIn1 = 32'd9151
; 
32'd181780: dataIn1 = 32'd9173
; 
32'd181781: dataIn1 = 32'd9176
; 
32'd181782: dataIn1 = 32'd2727
; 
32'd181783: dataIn1 = 32'd6669
; 
32'd181784: dataIn1 = 32'd8477
; 
32'd181785: dataIn1 = 32'd9149
; 
32'd181786: dataIn1 = 32'd9152
; 
32'd181787: dataIn1 = 32'd9153
; 
32'd181788: dataIn1 = 32'd9171
; 
32'd181789: dataIn1 = 32'd2727
; 
32'd181790: dataIn1 = 32'd6668
; 
32'd181791: dataIn1 = 32'd8522
; 
32'd181792: dataIn1 = 32'd9149
; 
32'd181793: dataIn1 = 32'd9152
; 
32'd181794: dataIn1 = 32'd9153
; 
32'd181795: dataIn1 = 32'd9174
; 
32'd181796: dataIn1 = 32'd6671
; 
32'd181797: dataIn1 = 32'd6672
; 
32'd181798: dataIn1 = 32'd9154
; 
32'd181799: dataIn1 = 32'd9155
; 
32'd181800: dataIn1 = 32'd9156
; 
32'd181801: dataIn1 = 32'd9157
; 
32'd181802: dataIn1 = 32'd9158
; 
32'd181803: dataIn1 = 32'd6670
; 
32'd181804: dataIn1 = 32'd6672
; 
32'd181805: dataIn1 = 32'd9154
; 
32'd181806: dataIn1 = 32'd9155
; 
32'd181807: dataIn1 = 32'd9156
; 
32'd181808: dataIn1 = 32'd9159
; 
32'd181809: dataIn1 = 32'd9160
; 
32'd181810: dataIn1 = 32'd6670
; 
32'd181811: dataIn1 = 32'd6671
; 
32'd181812: dataIn1 = 32'd9154
; 
32'd181813: dataIn1 = 32'd9155
; 
32'd181814: dataIn1 = 32'd9156
; 
32'd181815: dataIn1 = 32'd9161
; 
32'd181816: dataIn1 = 32'd9162
; 
32'd181817: dataIn1 = 32'd5294
; 
32'd181818: dataIn1 = 32'd6672
; 
32'd181819: dataIn1 = 32'd9150
; 
32'd181820: dataIn1 = 32'd9154
; 
32'd181821: dataIn1 = 32'd9157
; 
32'd181822: dataIn1 = 32'd9158
; 
32'd181823: dataIn1 = 32'd9169
; 
32'd181824: dataIn1 = 32'd5294
; 
32'd181825: dataIn1 = 32'd6671
; 
32'd181826: dataIn1 = 32'd9143
; 
32'd181827: dataIn1 = 32'd9154
; 
32'd181828: dataIn1 = 32'd9157
; 
32'd181829: dataIn1 = 32'd9158
; 
32'd181830: dataIn1 = 32'd9166
; 
32'd181831: dataIn1 = 32'd5238
; 
32'd181832: dataIn1 = 32'd6672
; 
32'd181833: dataIn1 = 32'd8478
; 
32'd181834: dataIn1 = 32'd9155
; 
32'd181835: dataIn1 = 32'd9159
; 
32'd181836: dataIn1 = 32'd9160
; 
32'd181837: dataIn1 = 32'd9170
; 
32'd181838: dataIn1 = 32'd5238
; 
32'd181839: dataIn1 = 32'd6670
; 
32'd181840: dataIn1 = 32'd8473
; 
32'd181841: dataIn1 = 32'd9155
; 
32'd181842: dataIn1 = 32'd9159
; 
32'd181843: dataIn1 = 32'd9160
; 
32'd181844: dataIn1 = 32'd9164
; 
32'd181845: dataIn1 = 32'd5225
; 
32'd181846: dataIn1 = 32'd6671
; 
32'd181847: dataIn1 = 32'd8356
; 
32'd181848: dataIn1 = 32'd9156
; 
32'd181849: dataIn1 = 32'd9161
; 
32'd181850: dataIn1 = 32'd9162
; 
32'd181851: dataIn1 = 32'd9168
; 
32'd181852: dataIn1 = 32'd5225
; 
32'd181853: dataIn1 = 32'd6670
; 
32'd181854: dataIn1 = 32'd8361
; 
32'd181855: dataIn1 = 32'd9156
; 
32'd181856: dataIn1 = 32'd9161
; 
32'd181857: dataIn1 = 32'd9162
; 
32'd181858: dataIn1 = 32'd9165
; 
32'd181859: dataIn1 = 32'd6452
; 
32'd181860: dataIn1 = 32'd6483
; 
32'd181861: dataIn1 = 32'd8363
; 
32'd181862: dataIn1 = 32'd8471
; 
32'd181863: dataIn1 = 32'd9163
; 
32'd181864: dataIn1 = 32'd9164
; 
32'd181865: dataIn1 = 32'd9165
; 
32'd181866: dataIn1 = 32'd6483
; 
32'd181867: dataIn1 = 32'd6670
; 
32'd181868: dataIn1 = 32'd8473
; 
32'd181869: dataIn1 = 32'd9160
; 
32'd181870: dataIn1 = 32'd9163
; 
32'd181871: dataIn1 = 32'd9164
; 
32'd181872: dataIn1 = 32'd9165
; 
32'd181873: dataIn1 = 32'd6452
; 
32'd181874: dataIn1 = 32'd6670
; 
32'd181875: dataIn1 = 32'd8361
; 
32'd181876: dataIn1 = 32'd9162
; 
32'd181877: dataIn1 = 32'd9163
; 
32'd181878: dataIn1 = 32'd9164
; 
32'd181879: dataIn1 = 32'd9165
; 
32'd181880: dataIn1 = 32'd6667
; 
32'd181881: dataIn1 = 32'd6671
; 
32'd181882: dataIn1 = 32'd9143
; 
32'd181883: dataIn1 = 32'd9158
; 
32'd181884: dataIn1 = 32'd9166
; 
32'd181885: dataIn1 = 32'd9167
; 
32'd181886: dataIn1 = 32'd9168
; 
32'd181887: dataIn1 = 32'd6451
; 
32'd181888: dataIn1 = 32'd6667
; 
32'd181889: dataIn1 = 32'd8357
; 
32'd181890: dataIn1 = 32'd9144
; 
32'd181891: dataIn1 = 32'd9166
; 
32'd181892: dataIn1 = 32'd9167
; 
32'd181893: dataIn1 = 32'd9168
; 
32'd181894: dataIn1 = 32'd6451
; 
32'd181895: dataIn1 = 32'd6671
; 
32'd181896: dataIn1 = 32'd8356
; 
32'd181897: dataIn1 = 32'd9161
; 
32'd181898: dataIn1 = 32'd9166
; 
32'd181899: dataIn1 = 32'd9167
; 
32'd181900: dataIn1 = 32'd9168
; 
32'd181901: dataIn1 = 32'd6669
; 
32'd181902: dataIn1 = 32'd6672
; 
32'd181903: dataIn1 = 32'd9150
; 
32'd181904: dataIn1 = 32'd9157
; 
32'd181905: dataIn1 = 32'd9169
; 
32'd181906: dataIn1 = 32'd9170
; 
32'd181907: dataIn1 = 32'd9171
; 
32'd181908: dataIn1 = 32'd6484
; 
32'd181909: dataIn1 = 32'd6672
; 
32'd181910: dataIn1 = 32'd8478
; 
32'd181911: dataIn1 = 32'd9159
; 
32'd181912: dataIn1 = 32'd9169
; 
32'd181913: dataIn1 = 32'd9170
; 
32'd181914: dataIn1 = 32'd9171
; 
32'd181915: dataIn1 = 32'd6484
; 
32'd181916: dataIn1 = 32'd6669
; 
32'd181917: dataIn1 = 32'd8477
; 
32'd181918: dataIn1 = 32'd9152
; 
32'd181919: dataIn1 = 32'd9169
; 
32'd181920: dataIn1 = 32'd9170
; 
32'd181921: dataIn1 = 32'd9171
; 
32'd181922: dataIn1 = 32'd6491
; 
32'd181923: dataIn1 = 32'd6673
; 
32'd181924: dataIn1 = 32'd8521
; 
32'd181925: dataIn1 = 32'd9172
; 
32'd181926: dataIn1 = 32'd9173
; 
32'd181927: dataIn1 = 32'd9174
; 
32'd181928: dataIn1 = 32'd9175
; 
32'd181929: dataIn1 = 32'd6668
; 
32'd181930: dataIn1 = 32'd6673
; 
32'd181931: dataIn1 = 32'd9151
; 
32'd181932: dataIn1 = 32'd9172
; 
32'd181933: dataIn1 = 32'd9173
; 
32'd181934: dataIn1 = 32'd9174
; 
32'd181935: dataIn1 = 32'd9176
; 
32'd181936: dataIn1 = 32'd6491
; 
32'd181937: dataIn1 = 32'd6668
; 
32'd181938: dataIn1 = 32'd8522
; 
32'd181939: dataIn1 = 32'd9153
; 
32'd181940: dataIn1 = 32'd9172
; 
32'd181941: dataIn1 = 32'd9173
; 
32'd181942: dataIn1 = 32'd9174
; 
32'd181943: dataIn1 = 32'd5239
; 
32'd181944: dataIn1 = 32'd6673
; 
32'd181945: dataIn1 = 32'd6795
; 
32'd181946: dataIn1 = 32'd8521
; 
32'd181947: dataIn1 = 32'd9172
; 
32'd181948: dataIn1 = 32'd9175
; 
32'd181949: dataIn1 = 32'd5295
; 
32'd181950: dataIn1 = 32'd6673
; 
32'd181951: dataIn1 = 32'd6794
; 
32'd181952: dataIn1 = 32'd9151
; 
32'd181953: dataIn1 = 32'd9173
; 
32'd181954: dataIn1 = 32'd9176
; 
32'd181955: dataIn1 = 32'd6444
; 
32'd181956: dataIn1 = 32'd6675
; 
32'd181957: dataIn1 = 32'd9177
; 
32'd181958: dataIn1 = 32'd9178
; 
32'd181959: dataIn1 = 32'd9179
; 
32'd181960: dataIn1 = 32'd9275
; 
32'd181961: dataIn1 = 32'd9285
; 
32'd181962: dataIn1 = 32'd6444
; 
32'd181963: dataIn1 = 32'd6666
; 
32'd181964: dataIn1 = 32'd8313
; 
32'd181965: dataIn1 = 32'd9145
; 
32'd181966: dataIn1 = 32'd9177
; 
32'd181967: dataIn1 = 32'd9178
; 
32'd181968: dataIn1 = 32'd9179
; 
32'd181969: dataIn1 = 32'd6666
; 
32'd181970: dataIn1 = 32'd6675
; 
32'd181971: dataIn1 = 32'd9146
; 
32'd181972: dataIn1 = 32'd9177
; 
32'd181973: dataIn1 = 32'd9178
; 
32'd181974: dataIn1 = 32'd9179
; 
32'd181975: dataIn1 = 32'd9180
; 
32'd181976: dataIn1 = 32'd5296
; 
32'd181977: dataIn1 = 32'd6674
; 
32'd181978: dataIn1 = 32'd6675
; 
32'd181979: dataIn1 = 32'd9146
; 
32'd181980: dataIn1 = 32'd9179
; 
32'd181981: dataIn1 = 32'd9180
; 
32'd181982: dataIn1 = 32'd6680
; 
32'd181983: dataIn1 = 32'd6681
; 
32'd181984: dataIn1 = 32'd9181
; 
32'd181985: dataIn1 = 32'd9182
; 
32'd181986: dataIn1 = 32'd9183
; 
32'd181987: dataIn1 = 32'd9184
; 
32'd181988: dataIn1 = 32'd9185
; 
32'd181989: dataIn1 = 32'd6679
; 
32'd181990: dataIn1 = 32'd6681
; 
32'd181991: dataIn1 = 32'd9181
; 
32'd181992: dataIn1 = 32'd9182
; 
32'd181993: dataIn1 = 32'd9183
; 
32'd181994: dataIn1 = 32'd9186
; 
32'd181995: dataIn1 = 32'd9187
; 
32'd181996: dataIn1 = 32'd6679
; 
32'd181997: dataIn1 = 32'd6680
; 
32'd181998: dataIn1 = 32'd9181
; 
32'd181999: dataIn1 = 32'd9182
; 
32'd182000: dataIn1 = 32'd9183
; 
32'd182001: dataIn1 = 32'd9188
; 
32'd182002: dataIn1 = 32'd9189
; 
32'd182003: dataIn1 = 32'd5299
; 
32'd182004: dataIn1 = 32'd6681
; 
32'd182005: dataIn1 = 32'd9181
; 
32'd182006: dataIn1 = 32'd9184
; 
32'd182007: dataIn1 = 32'd9185
; 
32'd182008: dataIn1 = 32'd9197
; 
32'd182009: dataIn1 = 32'd9200
; 
32'd182010: dataIn1 = 32'd5299
; 
32'd182011: dataIn1 = 32'd6680
; 
32'd182012: dataIn1 = 32'd9181
; 
32'd182013: dataIn1 = 32'd9184
; 
32'd182014: dataIn1 = 32'd9185
; 
32'd182015: dataIn1 = 32'd9190
; 
32'd182016: dataIn1 = 32'd9193
; 
32'd182017: dataIn1 = 32'd5300
; 
32'd182018: dataIn1 = 32'd6681
; 
32'd182019: dataIn1 = 32'd9182
; 
32'd182020: dataIn1 = 32'd9186
; 
32'd182021: dataIn1 = 32'd9187
; 
32'd182022: dataIn1 = 32'd9198
; 
32'd182023: dataIn1 = 32'd9201
; 
32'd182024: dataIn1 = 32'd5300
; 
32'd182025: dataIn1 = 32'd6679
; 
32'd182026: dataIn1 = 32'd6797
; 
32'd182027: dataIn1 = 32'd9182
; 
32'd182028: dataIn1 = 32'd9186
; 
32'd182029: dataIn1 = 32'd9187
; 
32'd182030: dataIn1 = 32'd5301
; 
32'd182031: dataIn1 = 32'd6680
; 
32'd182032: dataIn1 = 32'd9183
; 
32'd182033: dataIn1 = 32'd9188
; 
32'd182034: dataIn1 = 32'd9189
; 
32'd182035: dataIn1 = 32'd9192
; 
32'd182036: dataIn1 = 32'd9196
; 
32'd182037: dataIn1 = 32'd5301
; 
32'd182038: dataIn1 = 32'd6679
; 
32'd182039: dataIn1 = 32'd6796
; 
32'd182040: dataIn1 = 32'd9183
; 
32'd182041: dataIn1 = 32'd9188
; 
32'd182042: dataIn1 = 32'd9189
; 
32'd182043: dataIn1 = 32'd6680
; 
32'd182044: dataIn1 = 32'd6683
; 
32'd182045: dataIn1 = 32'd9185
; 
32'd182046: dataIn1 = 32'd9190
; 
32'd182047: dataIn1 = 32'd9191
; 
32'd182048: dataIn1 = 32'd9192
; 
32'd182049: dataIn1 = 32'd9193
; 
32'd182050: dataIn1 = 32'd6682
; 
32'd182051: dataIn1 = 32'd6683
; 
32'd182052: dataIn1 = 32'd9190
; 
32'd182053: dataIn1 = 32'd9191
; 
32'd182054: dataIn1 = 32'd9192
; 
32'd182055: dataIn1 = 32'd9194
; 
32'd182056: dataIn1 = 32'd9195
; 
32'd182057: dataIn1 = 32'd6680
; 
32'd182058: dataIn1 = 32'd6682
; 
32'd182059: dataIn1 = 32'd9188
; 
32'd182060: dataIn1 = 32'd9190
; 
32'd182061: dataIn1 = 32'd9191
; 
32'd182062: dataIn1 = 32'd9192
; 
32'd182063: dataIn1 = 32'd9196
; 
32'd182064: dataIn1 = 32'd5299
; 
32'd182065: dataIn1 = 32'd6683
; 
32'd182066: dataIn1 = 32'd9185
; 
32'd182067: dataIn1 = 32'd9190
; 
32'd182068: dataIn1 = 32'd9193
; 
32'd182069: dataIn1 = 32'd9208
; 
32'd182070: dataIn1 = 32'd9216
; 
32'd182071: dataIn1 = 32'd2728
; 
32'd182072: dataIn1 = 32'd6683
; 
32'd182073: dataIn1 = 32'd8610
; 
32'd182074: dataIn1 = 32'd9191
; 
32'd182075: dataIn1 = 32'd9194
; 
32'd182076: dataIn1 = 32'd9195
; 
32'd182077: dataIn1 = 32'd9217
; 
32'd182078: dataIn1 = 32'd2728
; 
32'd182079: dataIn1 = 32'd6682
; 
32'd182080: dataIn1 = 32'd8565
; 
32'd182081: dataIn1 = 32'd9191
; 
32'd182082: dataIn1 = 32'd9194
; 
32'd182083: dataIn1 = 32'd9195
; 
32'd182084: dataIn1 = 32'd9228
; 
32'd182085: dataIn1 = 32'd5301
; 
32'd182086: dataIn1 = 32'd6682
; 
32'd182087: dataIn1 = 32'd9188
; 
32'd182088: dataIn1 = 32'd9192
; 
32'd182089: dataIn1 = 32'd9196
; 
32'd182090: dataIn1 = 32'd9229
; 
32'd182091: dataIn1 = 32'd9231
; 
32'd182092: dataIn1 = 32'd6681
; 
32'd182093: dataIn1 = 32'd6685
; 
32'd182094: dataIn1 = 32'd9184
; 
32'd182095: dataIn1 = 32'd9197
; 
32'd182096: dataIn1 = 32'd9198
; 
32'd182097: dataIn1 = 32'd9199
; 
32'd182098: dataIn1 = 32'd9200
; 
32'd182099: dataIn1 = 32'd6681
; 
32'd182100: dataIn1 = 32'd6684
; 
32'd182101: dataIn1 = 32'd9186
; 
32'd182102: dataIn1 = 32'd9197
; 
32'd182103: dataIn1 = 32'd9198
; 
32'd182104: dataIn1 = 32'd9199
; 
32'd182105: dataIn1 = 32'd9201
; 
32'd182106: dataIn1 = 32'd6684
; 
32'd182107: dataIn1 = 32'd6685
; 
32'd182108: dataIn1 = 32'd9197
; 
32'd182109: dataIn1 = 32'd9198
; 
32'd182110: dataIn1 = 32'd9199
; 
32'd182111: dataIn1 = 32'd9202
; 
32'd182112: dataIn1 = 32'd9203
; 
32'd182113: dataIn1 = 32'd5299
; 
32'd182114: dataIn1 = 32'd6685
; 
32'd182115: dataIn1 = 32'd9184
; 
32'd182116: dataIn1 = 32'd9197
; 
32'd182117: dataIn1 = 32'd9200
; 
32'd182118: dataIn1 = 32'd9207
; 
32'd182119: dataIn1 = 32'd9219
; 
32'd182120: dataIn1 = 32'd5300
; 
32'd182121: dataIn1 = 32'd6684
; 
32'd182122: dataIn1 = 32'd9186
; 
32'd182123: dataIn1 = 32'd9198
; 
32'd182124: dataIn1 = 32'd9201
; 
32'd182125: dataIn1 = 32'd9223
; 
32'd182126: dataIn1 = 32'd9226
; 
32'd182127: dataIn1 = 32'd2732
; 
32'd182128: dataIn1 = 32'd6685
; 
32'd182129: dataIn1 = 32'd8730
; 
32'd182130: dataIn1 = 32'd9199
; 
32'd182131: dataIn1 = 32'd9202
; 
32'd182132: dataIn1 = 32'd9203
; 
32'd182133: dataIn1 = 32'd9221
; 
32'd182134: dataIn1 = 32'd2732
; 
32'd182135: dataIn1 = 32'd6684
; 
32'd182136: dataIn1 = 32'd8775
; 
32'd182137: dataIn1 = 32'd9199
; 
32'd182138: dataIn1 = 32'd9202
; 
32'd182139: dataIn1 = 32'd9203
; 
32'd182140: dataIn1 = 32'd9224
; 
32'd182141: dataIn1 = 32'd6687
; 
32'd182142: dataIn1 = 32'd6688
; 
32'd182143: dataIn1 = 32'd9204
; 
32'd182144: dataIn1 = 32'd9205
; 
32'd182145: dataIn1 = 32'd9206
; 
32'd182146: dataIn1 = 32'd9207
; 
32'd182147: dataIn1 = 32'd9208
; 
32'd182148: dataIn1 = 32'd6686
; 
32'd182149: dataIn1 = 32'd6688
; 
32'd182150: dataIn1 = 32'd9204
; 
32'd182151: dataIn1 = 32'd9205
; 
32'd182152: dataIn1 = 32'd9206
; 
32'd182153: dataIn1 = 32'd9209
; 
32'd182154: dataIn1 = 32'd9210
; 
32'd182155: dataIn1 = 32'd6686
; 
32'd182156: dataIn1 = 32'd6687
; 
32'd182157: dataIn1 = 32'd9204
; 
32'd182158: dataIn1 = 32'd9205
; 
32'd182159: dataIn1 = 32'd9206
; 
32'd182160: dataIn1 = 32'd9211
; 
32'd182161: dataIn1 = 32'd9212
; 
32'd182162: dataIn1 = 32'd5299
; 
32'd182163: dataIn1 = 32'd6688
; 
32'd182164: dataIn1 = 32'd9200
; 
32'd182165: dataIn1 = 32'd9204
; 
32'd182166: dataIn1 = 32'd9207
; 
32'd182167: dataIn1 = 32'd9208
; 
32'd182168: dataIn1 = 32'd9219
; 
32'd182169: dataIn1 = 32'd5299
; 
32'd182170: dataIn1 = 32'd6687
; 
32'd182171: dataIn1 = 32'd9193
; 
32'd182172: dataIn1 = 32'd9204
; 
32'd182173: dataIn1 = 32'd9207
; 
32'd182174: dataIn1 = 32'd9208
; 
32'd182175: dataIn1 = 32'd9216
; 
32'd182176: dataIn1 = 32'd5257
; 
32'd182177: dataIn1 = 32'd6688
; 
32'd182178: dataIn1 = 32'd8731
; 
32'd182179: dataIn1 = 32'd9205
; 
32'd182180: dataIn1 = 32'd9209
; 
32'd182181: dataIn1 = 32'd9210
; 
32'd182182: dataIn1 = 32'd9220
; 
32'd182183: dataIn1 = 32'd5257
; 
32'd182184: dataIn1 = 32'd6686
; 
32'd182185: dataIn1 = 32'd8726
; 
32'd182186: dataIn1 = 32'd9205
; 
32'd182187: dataIn1 = 32'd9209
; 
32'd182188: dataIn1 = 32'd9210
; 
32'd182189: dataIn1 = 32'd9214
; 
32'd182190: dataIn1 = 32'd5244
; 
32'd182191: dataIn1 = 32'd6687
; 
32'd182192: dataIn1 = 32'd8609
; 
32'd182193: dataIn1 = 32'd9206
; 
32'd182194: dataIn1 = 32'd9211
; 
32'd182195: dataIn1 = 32'd9212
; 
32'd182196: dataIn1 = 32'd9218
; 
32'd182197: dataIn1 = 32'd5244
; 
32'd182198: dataIn1 = 32'd6686
; 
32'd182199: dataIn1 = 32'd8614
; 
32'd182200: dataIn1 = 32'd9206
; 
32'd182201: dataIn1 = 32'd9211
; 
32'd182202: dataIn1 = 32'd9212
; 
32'd182203: dataIn1 = 32'd9215
; 
32'd182204: dataIn1 = 32'd6512
; 
32'd182205: dataIn1 = 32'd6543
; 
32'd182206: dataIn1 = 32'd8616
; 
32'd182207: dataIn1 = 32'd8724
; 
32'd182208: dataIn1 = 32'd9213
; 
32'd182209: dataIn1 = 32'd9214
; 
32'd182210: dataIn1 = 32'd9215
; 
32'd182211: dataIn1 = 32'd6543
; 
32'd182212: dataIn1 = 32'd6686
; 
32'd182213: dataIn1 = 32'd8726
; 
32'd182214: dataIn1 = 32'd9210
; 
32'd182215: dataIn1 = 32'd9213
; 
32'd182216: dataIn1 = 32'd9214
; 
32'd182217: dataIn1 = 32'd9215
; 
32'd182218: dataIn1 = 32'd6512
; 
32'd182219: dataIn1 = 32'd6686
; 
32'd182220: dataIn1 = 32'd8614
; 
32'd182221: dataIn1 = 32'd9212
; 
32'd182222: dataIn1 = 32'd9213
; 
32'd182223: dataIn1 = 32'd9214
; 
32'd182224: dataIn1 = 32'd9215
; 
32'd182225: dataIn1 = 32'd6683
; 
32'd182226: dataIn1 = 32'd6687
; 
32'd182227: dataIn1 = 32'd9193
; 
32'd182228: dataIn1 = 32'd9208
; 
32'd182229: dataIn1 = 32'd9216
; 
32'd182230: dataIn1 = 32'd9217
; 
32'd182231: dataIn1 = 32'd9218
; 
32'd182232: dataIn1 = 32'd6511
; 
32'd182233: dataIn1 = 32'd6683
; 
32'd182234: dataIn1 = 32'd8610
; 
32'd182235: dataIn1 = 32'd9194
; 
32'd182236: dataIn1 = 32'd9216
; 
32'd182237: dataIn1 = 32'd9217
; 
32'd182238: dataIn1 = 32'd9218
; 
32'd182239: dataIn1 = 32'd6511
; 
32'd182240: dataIn1 = 32'd6687
; 
32'd182241: dataIn1 = 32'd8609
; 
32'd182242: dataIn1 = 32'd9211
; 
32'd182243: dataIn1 = 32'd9216
; 
32'd182244: dataIn1 = 32'd9217
; 
32'd182245: dataIn1 = 32'd9218
; 
32'd182246: dataIn1 = 32'd6685
; 
32'd182247: dataIn1 = 32'd6688
; 
32'd182248: dataIn1 = 32'd9200
; 
32'd182249: dataIn1 = 32'd9207
; 
32'd182250: dataIn1 = 32'd9219
; 
32'd182251: dataIn1 = 32'd9220
; 
32'd182252: dataIn1 = 32'd9221
; 
32'd182253: dataIn1 = 32'd6544
; 
32'd182254: dataIn1 = 32'd6688
; 
32'd182255: dataIn1 = 32'd8731
; 
32'd182256: dataIn1 = 32'd9209
; 
32'd182257: dataIn1 = 32'd9219
; 
32'd182258: dataIn1 = 32'd9220
; 
32'd182259: dataIn1 = 32'd9221
; 
32'd182260: dataIn1 = 32'd6544
; 
32'd182261: dataIn1 = 32'd6685
; 
32'd182262: dataIn1 = 32'd8730
; 
32'd182263: dataIn1 = 32'd9202
; 
32'd182264: dataIn1 = 32'd9219
; 
32'd182265: dataIn1 = 32'd9220
; 
32'd182266: dataIn1 = 32'd9221
; 
32'd182267: dataIn1 = 32'd6551
; 
32'd182268: dataIn1 = 32'd6689
; 
32'd182269: dataIn1 = 32'd8774
; 
32'd182270: dataIn1 = 32'd9222
; 
32'd182271: dataIn1 = 32'd9223
; 
32'd182272: dataIn1 = 32'd9224
; 
32'd182273: dataIn1 = 32'd9225
; 
32'd182274: dataIn1 = 32'd6684
; 
32'd182275: dataIn1 = 32'd6689
; 
32'd182276: dataIn1 = 32'd9201
; 
32'd182277: dataIn1 = 32'd9222
; 
32'd182278: dataIn1 = 32'd9223
; 
32'd182279: dataIn1 = 32'd9224
; 
32'd182280: dataIn1 = 32'd9226
; 
32'd182281: dataIn1 = 32'd6551
; 
32'd182282: dataIn1 = 32'd6684
; 
32'd182283: dataIn1 = 32'd8775
; 
32'd182284: dataIn1 = 32'd9203
; 
32'd182285: dataIn1 = 32'd9222
; 
32'd182286: dataIn1 = 32'd9223
; 
32'd182287: dataIn1 = 32'd9224
; 
32'd182288: dataIn1 = 32'd5258
; 
32'd182289: dataIn1 = 32'd6689
; 
32'd182290: dataIn1 = 32'd6799
; 
32'd182291: dataIn1 = 32'd8774
; 
32'd182292: dataIn1 = 32'd9222
; 
32'd182293: dataIn1 = 32'd9225
; 
32'd182294: dataIn1 = 32'd5300
; 
32'd182295: dataIn1 = 32'd6689
; 
32'd182296: dataIn1 = 32'd6798
; 
32'd182297: dataIn1 = 32'd9201
; 
32'd182298: dataIn1 = 32'd9223
; 
32'd182299: dataIn1 = 32'd9226
; 
32'd182300: dataIn1 = 32'd6504
; 
32'd182301: dataIn1 = 32'd6690
; 
32'd182302: dataIn1 = 32'd8566
; 
32'd182303: dataIn1 = 32'd9227
; 
32'd182304: dataIn1 = 32'd9228
; 
32'd182305: dataIn1 = 32'd9229
; 
32'd182306: dataIn1 = 32'd9230
; 
32'd182307: dataIn1 = 32'd6504
; 
32'd182308: dataIn1 = 32'd6682
; 
32'd182309: dataIn1 = 32'd8565
; 
32'd182310: dataIn1 = 32'd9195
; 
32'd182311: dataIn1 = 32'd9227
; 
32'd182312: dataIn1 = 32'd9228
; 
32'd182313: dataIn1 = 32'd9229
; 
32'd182314: dataIn1 = 32'd6682
; 
32'd182315: dataIn1 = 32'd6690
; 
32'd182316: dataIn1 = 32'd9196
; 
32'd182317: dataIn1 = 32'd9227
; 
32'd182318: dataIn1 = 32'd9228
; 
32'd182319: dataIn1 = 32'd9229
; 
32'd182320: dataIn1 = 32'd9231
; 
32'd182321: dataIn1 = 32'd5243
; 
32'd182322: dataIn1 = 32'd6690
; 
32'd182323: dataIn1 = 32'd6801
; 
32'd182324: dataIn1 = 32'd8566
; 
32'd182325: dataIn1 = 32'd9227
; 
32'd182326: dataIn1 = 32'd9230
; 
32'd182327: dataIn1 = 32'd5301
; 
32'd182328: dataIn1 = 32'd6690
; 
32'd182329: dataIn1 = 32'd6800
; 
32'd182330: dataIn1 = 32'd9196
; 
32'd182331: dataIn1 = 32'd9229
; 
32'd182332: dataIn1 = 32'd9231
; 
32'd182333: dataIn1 = 32'd2631
; 
32'd182334: dataIn1 = 32'd6161
; 
32'd182335: dataIn1 = 32'd6703
; 
32'd182336: dataIn1 = 32'd7257
; 
32'd182337: dataIn1 = 32'd9232
; 
32'd182338: dataIn1 = 32'd9274
; 
32'd182339: dataIn1 = 32'd9286
; 
32'd182340: dataIn1 = 32'd1130
; 
32'd182341: dataIn1 = 32'd5214
; 
32'd182342: dataIn1 = 32'd6714
; 
32'd182343: dataIn1 = 32'd6715
; 
32'd182344: dataIn1 = 32'd6764
; 
32'd182345: dataIn1 = 32'd9233
; 
32'd182346: dataIn1 = 32'd1130
; 
32'd182347: dataIn1 = 32'd5292
; 
32'd182348: dataIn1 = 32'd6723
; 
32'd182349: dataIn1 = 32'd6725
; 
32'd182350: dataIn1 = 32'd6765
; 
32'd182351: dataIn1 = 32'd9234
; 
32'd182352: dataIn1 = 32'd2705
; 
32'd182353: dataIn1 = 32'd5154
; 
32'd182354: dataIn1 = 32'd6745
; 
32'd182355: dataIn1 = 32'd6747
; 
32'd182356: dataIn1 = 32'd9235
; 
32'd182357: dataIn1 = 32'd9287
; 
32'd182358: dataIn1 = 32'd2705
; 
32'd182359: dataIn1 = 32'd5157
; 
32'd182360: dataIn1 = 32'd6744
; 
32'd182361: dataIn1 = 32'd6748
; 
32'd182362: dataIn1 = 32'd9236
; 
32'd182363: dataIn1 = 32'd9290
; 
32'd182364: dataIn1 = 32'd1123
; 
32'd182365: dataIn1 = 32'd5154
; 
32'd182366: dataIn1 = 32'd6746
; 
32'd182367: dataIn1 = 32'd6753
; 
32'd182368: dataIn1 = 32'd9237
; 
32'd182369: dataIn1 = 32'd9288
; 
32'd182370: dataIn1 = 32'd1124
; 
32'd182371: dataIn1 = 32'd5157
; 
32'd182372: dataIn1 = 32'd6749
; 
32'd182373: dataIn1 = 32'd6750
; 
32'd182374: dataIn1 = 32'd9238
; 
32'd182375: dataIn1 = 32'd9289
; 
32'd182376: dataIn1 = 32'd1123
; 
32'd182377: dataIn1 = 32'd5283
; 
32'd182378: dataIn1 = 32'd6752
; 
32'd182379: dataIn1 = 32'd6791
; 
32'd182380: dataIn1 = 32'd9239
; 
32'd182381: dataIn1 = 32'd9291
; 
32'd182382: dataIn1 = 32'd2710
; 
32'd182383: dataIn1 = 32'd5173
; 
32'd182384: dataIn1 = 32'd6755
; 
32'd182385: dataIn1 = 32'd6757
; 
32'd182386: dataIn1 = 32'd9240
; 
32'd182387: dataIn1 = 32'd9293
; 
32'd182388: dataIn1 = 32'd2710
; 
32'd182389: dataIn1 = 32'd5176
; 
32'd182390: dataIn1 = 32'd6754
; 
32'd182391: dataIn1 = 32'd6758
; 
32'd182392: dataIn1 = 32'd9241
; 
32'd182393: dataIn1 = 32'd9296
; 
32'd182394: dataIn1 = 32'd1125
; 
32'd182395: dataIn1 = 32'd5173
; 
32'd182396: dataIn1 = 32'd6756
; 
32'd182397: dataIn1 = 32'd6763
; 
32'd182398: dataIn1 = 32'd9242
; 
32'd182399: dataIn1 = 32'd9294
; 
32'd182400: dataIn1 = 32'd1126
; 
32'd182401: dataIn1 = 32'd5176
; 
32'd182402: dataIn1 = 32'd6759
; 
32'd182403: dataIn1 = 32'd6760
; 
32'd182404: dataIn1 = 32'd9243
; 
32'd182405: dataIn1 = 32'd9295
; 
32'd182406: dataIn1 = 32'd1126
; 
32'd182407: dataIn1 = 32'd5282
; 
32'd182408: dataIn1 = 32'd6761
; 
32'd182409: dataIn1 = 32'd6789
; 
32'd182410: dataIn1 = 32'd9244
; 
32'd182411: dataIn1 = 32'd9297
; 
32'd182412: dataIn1 = 32'd1125
; 
32'd182413: dataIn1 = 32'd5288
; 
32'd182414: dataIn1 = 32'd6762
; 
32'd182415: dataIn1 = 32'd6793
; 
32'd182416: dataIn1 = 32'd9245
; 
32'd182417: dataIn1 = 32'd9281
; 
32'd182418: dataIn1 = 32'd2725
; 
32'd182419: dataIn1 = 32'd5230
; 
32'd182420: dataIn1 = 32'd6767
; 
32'd182421: dataIn1 = 32'd6769
; 
32'd182422: dataIn1 = 32'd9246
; 
32'd182423: dataIn1 = 32'd9299
; 
32'd182424: dataIn1 = 32'd2725
; 
32'd182425: dataIn1 = 32'd5233
; 
32'd182426: dataIn1 = 32'd6766
; 
32'd182427: dataIn1 = 32'd6770
; 
32'd182428: dataIn1 = 32'd9247
; 
32'd182429: dataIn1 = 32'd9302
; 
32'd182430: dataIn1 = 32'd1131
; 
32'd182431: dataIn1 = 32'd5230
; 
32'd182432: dataIn1 = 32'd6768
; 
32'd182433: dataIn1 = 32'd6775
; 
32'd182434: dataIn1 = 32'd9248
; 
32'd182435: dataIn1 = 32'd9300
; 
32'd182436: dataIn1 = 32'd1132
; 
32'd182437: dataIn1 = 32'd5233
; 
32'd182438: dataIn1 = 32'd6771
; 
32'd182439: dataIn1 = 32'd6772
; 
32'd182440: dataIn1 = 32'd9249
; 
32'd182441: dataIn1 = 32'd9301
; 
32'd182442: dataIn1 = 32'd1132
; 
32'd182443: dataIn1 = 32'd5297
; 
32'd182444: dataIn1 = 32'd6773
; 
32'd182445: dataIn1 = 32'd6795
; 
32'd182446: dataIn1 = 32'd9250
; 
32'd182447: dataIn1 = 32'd9283
; 
32'd182448: dataIn1 = 32'd1131
; 
32'd182449: dataIn1 = 32'd5303
; 
32'd182450: dataIn1 = 32'd6774
; 
32'd182451: dataIn1 = 32'd6801
; 
32'd182452: dataIn1 = 32'd9251
; 
32'd182453: dataIn1 = 32'd9303
; 
32'd182454: dataIn1 = 32'd2730
; 
32'd182455: dataIn1 = 32'd5249
; 
32'd182456: dataIn1 = 32'd6777
; 
32'd182457: dataIn1 = 32'd6779
; 
32'd182458: dataIn1 = 32'd9252
; 
32'd182459: dataIn1 = 32'd9305
; 
32'd182460: dataIn1 = 32'd2730
; 
32'd182461: dataIn1 = 32'd5252
; 
32'd182462: dataIn1 = 32'd6776
; 
32'd182463: dataIn1 = 32'd6780
; 
32'd182464: dataIn1 = 32'd9253
; 
32'd182465: dataIn1 = 32'd9308
; 
32'd182466: dataIn1 = 32'd1133
; 
32'd182467: dataIn1 = 32'd5249
; 
32'd182468: dataIn1 = 32'd6778
; 
32'd182469: dataIn1 = 32'd6785
; 
32'd182470: dataIn1 = 32'd9254
; 
32'd182471: dataIn1 = 32'd9306
; 
32'd182472: dataIn1 = 32'd1134
; 
32'd182473: dataIn1 = 32'd5252
; 
32'd182474: dataIn1 = 32'd6781
; 
32'd182475: dataIn1 = 32'd6782
; 
32'd182476: dataIn1 = 32'd9255
; 
32'd182477: dataIn1 = 32'd9307
; 
32'd182478: dataIn1 = 32'd1134
; 
32'd182479: dataIn1 = 32'd5302
; 
32'd182480: dataIn1 = 32'd6783
; 
32'd182481: dataIn1 = 32'd6799
; 
32'd182482: dataIn1 = 32'd9256
; 
32'd182483: dataIn1 = 32'd9309
; 
32'd182484: dataIn1 = 32'd1133
; 
32'd182485: dataIn1 = 32'd5648
; 
32'd182486: dataIn1 = 32'd6784
; 
32'd182487: dataIn1 = 32'd6849
; 
32'd182488: dataIn1 = 32'd9257
; 
32'd182489: dataIn1 = 32'd9268
; 
32'd182490: dataIn1 = 32'd9269
; 
32'd182491: dataIn1 = 32'd2747
; 
32'd182492: dataIn1 = 32'd5282
; 
32'd182493: dataIn1 = 32'd6787
; 
32'd182494: dataIn1 = 32'd6788
; 
32'd182495: dataIn1 = 32'd9258
; 
32'd182496: dataIn1 = 32'd9298
; 
32'd182497: dataIn1 = 32'd2747
; 
32'd182498: dataIn1 = 32'd5283
; 
32'd182499: dataIn1 = 32'd6786
; 
32'd182500: dataIn1 = 32'd6790
; 
32'd182501: dataIn1 = 32'd9259
; 
32'd182502: dataIn1 = 32'd9292
; 
32'd182503: dataIn1 = 32'd2752
; 
32'd182504: dataIn1 = 32'd5302
; 
32'd182505: dataIn1 = 32'd6797
; 
32'd182506: dataIn1 = 32'd6798
; 
32'd182507: dataIn1 = 32'd9260
; 
32'd182508: dataIn1 = 32'd9310
; 
32'd182509: dataIn1 = 32'd2752
; 
32'd182510: dataIn1 = 32'd5303
; 
32'd182511: dataIn1 = 32'd6796
; 
32'd182512: dataIn1 = 32'd6800
; 
32'd182513: dataIn1 = 32'd9261
; 
32'd182514: dataIn1 = 32'd9304
; 
32'd182515: dataIn1 = 32'd1120
; 
32'd182516: dataIn1 = 32'd6693
; 
32'd182517: dataIn1 = 32'd6706
; 
32'd182518: dataIn1 = 32'd6820
; 
32'd182519: dataIn1 = 32'd9262
; 
32'd182520: dataIn1 = 32'd9263
; 
32'd182521: dataIn1 = 32'd9312
; 
32'd182522: dataIn1 = 32'd5639
; 
32'd182523: dataIn1 = 32'd6693
; 
32'd182524: dataIn1 = 32'd6819
; 
32'd182525: dataIn1 = 32'd6820
; 
32'd182526: dataIn1 = 32'd9262
; 
32'd182527: dataIn1 = 32'd9263
; 
32'd182528: dataIn1 = 32'd9265
; 
32'd182529: dataIn1 = 32'd9311
; 
32'd182530: dataIn1 = 32'd5641
; 
32'd182531: dataIn1 = 32'd6692
; 
32'd182532: dataIn1 = 32'd6824
; 
32'd182533: dataIn1 = 32'd6826
; 
32'd182534: dataIn1 = 32'd9264
; 
32'd182535: dataIn1 = 32'd9265
; 
32'd182536: dataIn1 = 32'd9313
; 
32'd182537: dataIn1 = 32'd10286
; 
32'd182538: dataIn1 = 32'd3583
; 
32'd182539: dataIn1 = 32'd6692
; 
32'd182540: dataIn1 = 32'd6819
; 
32'd182541: dataIn1 = 32'd6824
; 
32'd182542: dataIn1 = 32'd9263
; 
32'd182543: dataIn1 = 32'd9264
; 
32'd182544: dataIn1 = 32'd9265
; 
32'd182545: dataIn1 = 32'd9311
; 
32'd182546: dataIn1 = 32'd2105
; 
32'd182547: dataIn1 = 32'd5647
; 
32'd182548: dataIn1 = 32'd6695
; 
32'd182549: dataIn1 = 32'd6845
; 
32'd182550: dataIn1 = 32'd9266
; 
32'd182551: dataIn1 = 32'd9267
; 
32'd182552: dataIn1 = 32'd9316
; 
32'd182553: dataIn1 = 32'd10290
; 
32'd182554: dataIn1 = 32'd3585
; 
32'd182555: dataIn1 = 32'd6695
; 
32'd182556: dataIn1 = 32'd6845
; 
32'd182557: dataIn1 = 32'd6850
; 
32'd182558: dataIn1 = 32'd9266
; 
32'd182559: dataIn1 = 32'd9267
; 
32'd182560: dataIn1 = 32'd9269
; 
32'd182561: dataIn1 = 32'd9315
; 
32'd182562: dataIn1 = 32'd1133
; 
32'd182563: dataIn1 = 32'd6694
; 
32'd182564: dataIn1 = 32'd9257
; 
32'd182565: dataIn1 = 32'd9268
; 
32'd182566: dataIn1 = 32'd9269
; 
32'd182567: dataIn1 = 32'd9306
; 
32'd182568: dataIn1 = 32'd9318
; 
32'd182569: dataIn1 = 32'd5648
; 
32'd182570: dataIn1 = 32'd6694
; 
32'd182571: dataIn1 = 32'd6850
; 
32'd182572: dataIn1 = 32'd9257
; 
32'd182573: dataIn1 = 32'd9267
; 
32'd182574: dataIn1 = 32'd9268
; 
32'd182575: dataIn1 = 32'd9269
; 
32'd182576: dataIn1 = 32'd9315
; 
32'd182577: dataIn1 = 32'd2320
; 
32'd182578: dataIn1 = 32'd3965
; 
32'd182579: dataIn1 = 32'd5828
; 
32'd182580: dataIn1 = 32'd5844
; 
32'd182581: dataIn1 = 32'd6858
; 
32'd182582: dataIn1 = 32'd9270
; 
32'd182583: dataIn1 = 32'd9271
; 
32'd182584: dataIn1 = 32'd9319
; 
32'd182585: dataIn1 = 32'd2320
; 
32'd182586: dataIn1 = 32'd3963
; 
32'd182587: dataIn1 = 32'd3967
; 
32'd182588: dataIn1 = 32'd5828
; 
32'd182589: dataIn1 = 32'd6855
; 
32'd182590: dataIn1 = 32'd9270
; 
32'd182591: dataIn1 = 32'd9271
; 
32'd182592: dataIn1 = 32'd2325
; 
32'd182593: dataIn1 = 32'd3984
; 
32'd182594: dataIn1 = 32'd5271
; 
32'd182595: dataIn1 = 32'd5877
; 
32'd182596: dataIn1 = 32'd9272
; 
32'd182597: dataIn1 = 32'd9273
; 
32'd182598: dataIn1 = 32'd3981
; 
32'd182599: dataIn1 = 32'd3984
; 
32'd182600: dataIn1 = 32'd5877
; 
32'd182601: dataIn1 = 32'd5880
; 
32'd182602: dataIn1 = 32'd7008
; 
32'd182603: dataIn1 = 32'd9272
; 
32'd182604: dataIn1 = 32'd9273
; 
32'd182605: dataIn1 = 32'd9320
; 
32'd182606: dataIn1 = 32'd2631
; 
32'd182607: dataIn1 = 32'd6059
; 
32'd182608: dataIn1 = 32'd6163
; 
32'd182609: dataIn1 = 32'd7260
; 
32'd182610: dataIn1 = 32'd9232
; 
32'd182611: dataIn1 = 32'd9274
; 
32'd182612: dataIn1 = 32'd9286
; 
32'd182613: dataIn1 = 32'd5224
; 
32'd182614: dataIn1 = 32'd6444
; 
32'd182615: dataIn1 = 32'd8308
; 
32'd182616: dataIn1 = 32'd8312
; 
32'd182617: dataIn1 = 32'd9177
; 
32'd182618: dataIn1 = 32'd9275
; 
32'd182619: dataIn1 = 32'd9285
; 
32'd182620: dataIn1 = 32'd2733
; 
32'd182621: dataIn1 = 32'd6564
; 
32'd182622: dataIn1 = 32'd8796
; 
32'd182623: dataIn1 = 32'd8816
; 
32'd182624: dataIn1 = 32'd9276
; 
32'd182625: dataIn1 = 32'd9405
; 
32'd182626: dataIn1 = 32'd9443
; 
32'd182627: dataIn1 = 32'd2743
; 
32'd182628: dataIn1 = 32'd5276
; 
32'd182629: dataIn1 = 32'd5278
; 
32'd182630: dataIn1 = 32'd6599
; 
32'd182631: dataIn1 = 32'd8935
; 
32'd182632: dataIn1 = 32'd9277
; 
32'd182633: dataIn1 = 32'd9278
; 
32'd182634: dataIn1 = 32'd2743
; 
32'd182635: dataIn1 = 32'd5275
; 
32'd182636: dataIn1 = 32'd6599
; 
32'd182637: dataIn1 = 32'd8933
; 
32'd182638: dataIn1 = 32'd9277
; 
32'd182639: dataIn1 = 32'd9278
; 
32'd182640: dataIn1 = 32'd9279
; 
32'd182641: dataIn1 = 32'd9321
; 
32'd182642: dataIn1 = 32'd5275
; 
32'd182643: dataIn1 = 32'd5277
; 
32'd182644: dataIn1 = 32'd6609
; 
32'd182645: dataIn1 = 32'd8974
; 
32'd182646: dataIn1 = 32'd9278
; 
32'd182647: dataIn1 = 32'd9279
; 
32'd182648: dataIn1 = 32'd9280
; 
32'd182649: dataIn1 = 32'd9321
; 
32'd182650: dataIn1 = 32'd5163
; 
32'd182651: dataIn1 = 32'd5277
; 
32'd182652: dataIn1 = 32'd6609
; 
32'd182653: dataIn1 = 32'd6751
; 
32'd182654: dataIn1 = 32'd8973
; 
32'd182655: dataIn1 = 32'd9279
; 
32'd182656: dataIn1 = 32'd9280
; 
32'd182657: dataIn1 = 32'd9322
; 
32'd182658: dataIn1 = 32'd1125
; 
32'd182659: dataIn1 = 32'd5288
; 
32'd182660: dataIn1 = 32'd5447
; 
32'd182661: dataIn1 = 32'd9245
; 
32'd182662: dataIn1 = 32'd9281
; 
32'd182663: dataIn1 = 32'd9282
; 
32'd182664: dataIn1 = 32'd9294
; 
32'd182665: dataIn1 = 32'd9324
; 
32'd182666: dataIn1 = 32'd2749
; 
32'd182667: dataIn1 = 32'd5288
; 
32'd182668: dataIn1 = 32'd5447
; 
32'd182669: dataIn1 = 32'd6722
; 
32'd182670: dataIn1 = 32'd9036
; 
32'd182671: dataIn1 = 32'd9281
; 
32'd182672: dataIn1 = 32'd9282
; 
32'd182673: dataIn1 = 32'd9323
; 
32'd182674: dataIn1 = 32'd1132
; 
32'd182675: dataIn1 = 32'd5297
; 
32'd182676: dataIn1 = 32'd5452
; 
32'd182677: dataIn1 = 32'd9250
; 
32'd182678: dataIn1 = 32'd9283
; 
32'd182679: dataIn1 = 32'd9284
; 
32'd182680: dataIn1 = 32'd9301
; 
32'd182681: dataIn1 = 32'd9326
; 
32'd182682: dataIn1 = 32'd2751
; 
32'd182683: dataIn1 = 32'd5297
; 
32'd182684: dataIn1 = 32'd5452
; 
32'd182685: dataIn1 = 32'd6729
; 
32'd182686: dataIn1 = 32'd9139
; 
32'd182687: dataIn1 = 32'd9283
; 
32'd182688: dataIn1 = 32'd9284
; 
32'd182689: dataIn1 = 32'd9325
; 
32'd182690: dataIn1 = 32'd5224
; 
32'd182691: dataIn1 = 32'd6675
; 
32'd182692: dataIn1 = 32'd6676
; 
32'd182693: dataIn1 = 32'd9177
; 
32'd182694: dataIn1 = 32'd9275
; 
32'd182695: dataIn1 = 32'd9285
; 
32'd182696: dataIn1 = 32'd6161
; 
32'd182697: dataIn1 = 32'd6163
; 
32'd182698: dataIn1 = 32'd9232
; 
32'd182699: dataIn1 = 32'd9274
; 
32'd182700: dataIn1 = 32'd9286
; 
32'd182701: dataIn1 = 32'd10151
; 
32'd182702: dataIn1 = 32'd10220
; 
32'd182703: dataIn1 = 32'd2705
; 
32'd182704: dataIn1 = 32'd5154
; 
32'd182705: dataIn1 = 32'd5434
; 
32'd182706: dataIn1 = 32'd9235
; 
32'd182707: dataIn1 = 32'd9287
; 
32'd182708: dataIn1 = 32'd9288
; 
32'd182709: dataIn1 = 32'd9290
; 
32'd182710: dataIn1 = 32'd9328
; 
32'd182711: dataIn1 = 32'd1123
; 
32'd182712: dataIn1 = 32'd5154
; 
32'd182713: dataIn1 = 32'd5434
; 
32'd182714: dataIn1 = 32'd9237
; 
32'd182715: dataIn1 = 32'd9287
; 
32'd182716: dataIn1 = 32'd9288
; 
32'd182717: dataIn1 = 32'd9291
; 
32'd182718: dataIn1 = 32'd9327
; 
32'd182719: dataIn1 = 32'd1124
; 
32'd182720: dataIn1 = 32'd5157
; 
32'd182721: dataIn1 = 32'd5433
; 
32'd182722: dataIn1 = 32'd9238
; 
32'd182723: dataIn1 = 32'd9289
; 
32'd182724: dataIn1 = 32'd9290
; 
32'd182725: dataIn1 = 32'd9337
; 
32'd182726: dataIn1 = 32'd9339
; 
32'd182727: dataIn1 = 32'd2705
; 
32'd182728: dataIn1 = 32'd5157
; 
32'd182729: dataIn1 = 32'd5433
; 
32'd182730: dataIn1 = 32'd9236
; 
32'd182731: dataIn1 = 32'd9287
; 
32'd182732: dataIn1 = 32'd9289
; 
32'd182733: dataIn1 = 32'd9290
; 
32'd182734: dataIn1 = 32'd9328
; 
32'd182735: dataIn1 = 32'd1123
; 
32'd182736: dataIn1 = 32'd5283
; 
32'd182737: dataIn1 = 32'd5445
; 
32'd182738: dataIn1 = 32'd9239
; 
32'd182739: dataIn1 = 32'd9288
; 
32'd182740: dataIn1 = 32'd9291
; 
32'd182741: dataIn1 = 32'd9292
; 
32'd182742: dataIn1 = 32'd9327
; 
32'd182743: dataIn1 = 32'd2747
; 
32'd182744: dataIn1 = 32'd5283
; 
32'd182745: dataIn1 = 32'd5445
; 
32'd182746: dataIn1 = 32'd9259
; 
32'd182747: dataIn1 = 32'd9291
; 
32'd182748: dataIn1 = 32'd9292
; 
32'd182749: dataIn1 = 32'd9298
; 
32'd182750: dataIn1 = 32'd9329
; 
32'd182751: dataIn1 = 32'd2710
; 
32'd182752: dataIn1 = 32'd5173
; 
32'd182753: dataIn1 = 32'd5436
; 
32'd182754: dataIn1 = 32'd9240
; 
32'd182755: dataIn1 = 32'd9293
; 
32'd182756: dataIn1 = 32'd9294
; 
32'd182757: dataIn1 = 32'd9296
; 
32'd182758: dataIn1 = 32'd9330
; 
32'd182759: dataIn1 = 32'd1125
; 
32'd182760: dataIn1 = 32'd5173
; 
32'd182761: dataIn1 = 32'd5436
; 
32'd182762: dataIn1 = 32'd9242
; 
32'd182763: dataIn1 = 32'd9281
; 
32'd182764: dataIn1 = 32'd9293
; 
32'd182765: dataIn1 = 32'd9294
; 
32'd182766: dataIn1 = 32'd9324
; 
32'd182767: dataIn1 = 32'd1126
; 
32'd182768: dataIn1 = 32'd5176
; 
32'd182769: dataIn1 = 32'd5435
; 
32'd182770: dataIn1 = 32'd9243
; 
32'd182771: dataIn1 = 32'd9295
; 
32'd182772: dataIn1 = 32'd9296
; 
32'd182773: dataIn1 = 32'd9297
; 
32'd182774: dataIn1 = 32'd9331
; 
32'd182775: dataIn1 = 32'd2710
; 
32'd182776: dataIn1 = 32'd5176
; 
32'd182777: dataIn1 = 32'd5435
; 
32'd182778: dataIn1 = 32'd9241
; 
32'd182779: dataIn1 = 32'd9293
; 
32'd182780: dataIn1 = 32'd9295
; 
32'd182781: dataIn1 = 32'd9296
; 
32'd182782: dataIn1 = 32'd9330
; 
32'd182783: dataIn1 = 32'd1126
; 
32'd182784: dataIn1 = 32'd5282
; 
32'd182785: dataIn1 = 32'd5446
; 
32'd182786: dataIn1 = 32'd9244
; 
32'd182787: dataIn1 = 32'd9295
; 
32'd182788: dataIn1 = 32'd9297
; 
32'd182789: dataIn1 = 32'd9298
; 
32'd182790: dataIn1 = 32'd9331
; 
32'd182791: dataIn1 = 32'd2747
; 
32'd182792: dataIn1 = 32'd5282
; 
32'd182793: dataIn1 = 32'd5446
; 
32'd182794: dataIn1 = 32'd9258
; 
32'd182795: dataIn1 = 32'd9292
; 
32'd182796: dataIn1 = 32'd9297
; 
32'd182797: dataIn1 = 32'd9298
; 
32'd182798: dataIn1 = 32'd9329
; 
32'd182799: dataIn1 = 32'd2725
; 
32'd182800: dataIn1 = 32'd5230
; 
32'd182801: dataIn1 = 32'd5442
; 
32'd182802: dataIn1 = 32'd9246
; 
32'd182803: dataIn1 = 32'd9299
; 
32'd182804: dataIn1 = 32'd9300
; 
32'd182805: dataIn1 = 32'd9302
; 
32'd182806: dataIn1 = 32'd9333
; 
32'd182807: dataIn1 = 32'd1131
; 
32'd182808: dataIn1 = 32'd5230
; 
32'd182809: dataIn1 = 32'd5442
; 
32'd182810: dataIn1 = 32'd9248
; 
32'd182811: dataIn1 = 32'd9299
; 
32'd182812: dataIn1 = 32'd9300
; 
32'd182813: dataIn1 = 32'd9303
; 
32'd182814: dataIn1 = 32'd9332
; 
32'd182815: dataIn1 = 32'd1132
; 
32'd182816: dataIn1 = 32'd5233
; 
32'd182817: dataIn1 = 32'd5441
; 
32'd182818: dataIn1 = 32'd9249
; 
32'd182819: dataIn1 = 32'd9283
; 
32'd182820: dataIn1 = 32'd9301
; 
32'd182821: dataIn1 = 32'd9302
; 
32'd182822: dataIn1 = 32'd9326
; 
32'd182823: dataIn1 = 32'd2725
; 
32'd182824: dataIn1 = 32'd5233
; 
32'd182825: dataIn1 = 32'd5441
; 
32'd182826: dataIn1 = 32'd9247
; 
32'd182827: dataIn1 = 32'd9299
; 
32'd182828: dataIn1 = 32'd9301
; 
32'd182829: dataIn1 = 32'd9302
; 
32'd182830: dataIn1 = 32'd9333
; 
32'd182831: dataIn1 = 32'd1131
; 
32'd182832: dataIn1 = 32'd5303
; 
32'd182833: dataIn1 = 32'd5453
; 
32'd182834: dataIn1 = 32'd9251
; 
32'd182835: dataIn1 = 32'd9300
; 
32'd182836: dataIn1 = 32'd9303
; 
32'd182837: dataIn1 = 32'd9304
; 
32'd182838: dataIn1 = 32'd9332
; 
32'd182839: dataIn1 = 32'd2752
; 
32'd182840: dataIn1 = 32'd5303
; 
32'd182841: dataIn1 = 32'd5453
; 
32'd182842: dataIn1 = 32'd9261
; 
32'd182843: dataIn1 = 32'd9303
; 
32'd182844: dataIn1 = 32'd9304
; 
32'd182845: dataIn1 = 32'd9310
; 
32'd182846: dataIn1 = 32'd9334
; 
32'd182847: dataIn1 = 32'd2730
; 
32'd182848: dataIn1 = 32'd5249
; 
32'd182849: dataIn1 = 32'd5444
; 
32'd182850: dataIn1 = 32'd9252
; 
32'd182851: dataIn1 = 32'd9305
; 
32'd182852: dataIn1 = 32'd9306
; 
32'd182853: dataIn1 = 32'd9308
; 
32'd182854: dataIn1 = 32'd9335
; 
32'd182855: dataIn1 = 32'd1133
; 
32'd182856: dataIn1 = 32'd5249
; 
32'd182857: dataIn1 = 32'd5444
; 
32'd182858: dataIn1 = 32'd9254
; 
32'd182859: dataIn1 = 32'd9268
; 
32'd182860: dataIn1 = 32'd9305
; 
32'd182861: dataIn1 = 32'd9306
; 
32'd182862: dataIn1 = 32'd9318
; 
32'd182863: dataIn1 = 32'd1134
; 
32'd182864: dataIn1 = 32'd5252
; 
32'd182865: dataIn1 = 32'd5443
; 
32'd182866: dataIn1 = 32'd9255
; 
32'd182867: dataIn1 = 32'd9307
; 
32'd182868: dataIn1 = 32'd9308
; 
32'd182869: dataIn1 = 32'd9309
; 
32'd182870: dataIn1 = 32'd9336
; 
32'd182871: dataIn1 = 32'd2730
; 
32'd182872: dataIn1 = 32'd5252
; 
32'd182873: dataIn1 = 32'd5443
; 
32'd182874: dataIn1 = 32'd9253
; 
32'd182875: dataIn1 = 32'd9305
; 
32'd182876: dataIn1 = 32'd9307
; 
32'd182877: dataIn1 = 32'd9308
; 
32'd182878: dataIn1 = 32'd9335
; 
32'd182879: dataIn1 = 32'd1134
; 
32'd182880: dataIn1 = 32'd5302
; 
32'd182881: dataIn1 = 32'd5454
; 
32'd182882: dataIn1 = 32'd9256
; 
32'd182883: dataIn1 = 32'd9307
; 
32'd182884: dataIn1 = 32'd9309
; 
32'd182885: dataIn1 = 32'd9310
; 
32'd182886: dataIn1 = 32'd9336
; 
32'd182887: dataIn1 = 32'd2752
; 
32'd182888: dataIn1 = 32'd5302
; 
32'd182889: dataIn1 = 32'd5454
; 
32'd182890: dataIn1 = 32'd9260
; 
32'd182891: dataIn1 = 32'd9304
; 
32'd182892: dataIn1 = 32'd9309
; 
32'd182893: dataIn1 = 32'd9310
; 
32'd182894: dataIn1 = 32'd9334
; 
32'd182895: dataIn1 = 32'd2102
; 
32'd182896: dataIn1 = 32'd6692
; 
32'd182897: dataIn1 = 32'd6693
; 
32'd182898: dataIn1 = 32'd9263
; 
32'd182899: dataIn1 = 32'd9265
; 
32'd182900: dataIn1 = 32'd9311
; 
32'd182901: dataIn1 = 32'd9314
; 
32'd182902: dataIn1 = 32'd2102
; 
32'd182903: dataIn1 = 32'd5431
; 
32'd182904: dataIn1 = 32'd6693
; 
32'd182905: dataIn1 = 32'd6706
; 
32'd182906: dataIn1 = 32'd6730
; 
32'd182907: dataIn1 = 32'd9262
; 
32'd182908: dataIn1 = 32'd9312
; 
32'd182909: dataIn1 = 32'd13
; 
32'd182910: dataIn1 = 32'd6692
; 
32'd182911: dataIn1 = 32'd9264
; 
32'd182912: dataIn1 = 32'd9313
; 
32'd182913: dataIn1 = 32'd9314
; 
32'd182914: dataIn1 = 32'd10286
; 
32'd182915: dataIn1 = 32'd13
; 
32'd182916: dataIn1 = 32'd2102
; 
32'd182917: dataIn1 = 32'd3457
; 
32'd182918: dataIn1 = 32'd3467
; 
32'd182919: dataIn1 = 32'd6692
; 
32'd182920: dataIn1 = 32'd9311
; 
32'd182921: dataIn1 = 32'd9313
; 
32'd182922: dataIn1 = 32'd9314
; 
32'd182923: dataIn1 = 32'd2104
; 
32'd182924: dataIn1 = 32'd6694
; 
32'd182925: dataIn1 = 32'd6695
; 
32'd182926: dataIn1 = 32'd9267
; 
32'd182927: dataIn1 = 32'd9269
; 
32'd182928: dataIn1 = 32'd9315
; 
32'd182929: dataIn1 = 32'd9317
; 
32'd182930: dataIn1 = 32'd23
; 
32'd182931: dataIn1 = 32'd6695
; 
32'd182932: dataIn1 = 32'd9266
; 
32'd182933: dataIn1 = 32'd9316
; 
32'd182934: dataIn1 = 32'd9317
; 
32'd182935: dataIn1 = 32'd10290
; 
32'd182936: dataIn1 = 32'd23
; 
32'd182937: dataIn1 = 32'd2104
; 
32'd182938: dataIn1 = 32'd2120
; 
32'd182939: dataIn1 = 32'd2121
; 
32'd182940: dataIn1 = 32'd6695
; 
32'd182941: dataIn1 = 32'd9315
; 
32'd182942: dataIn1 = 32'd9316
; 
32'd182943: dataIn1 = 32'd9317
; 
32'd182944: dataIn1 = 32'd2104
; 
32'd182945: dataIn1 = 32'd5444
; 
32'd182946: dataIn1 = 32'd6694
; 
32'd182947: dataIn1 = 32'd6731
; 
32'd182948: dataIn1 = 32'd9268
; 
32'd182949: dataIn1 = 32'd9306
; 
32'd182950: dataIn1 = 32'd9318
; 
32'd182951: dataIn1 = 32'd2320
; 
32'd182952: dataIn1 = 32'd3970
; 
32'd182953: dataIn1 = 32'd3979
; 
32'd182954: dataIn1 = 32'd5844
; 
32'd182955: dataIn1 = 32'd9270
; 
32'd182956: dataIn1 = 32'd9319
; 
32'd182957: dataIn1 = 32'd451
; 
32'd182958: dataIn1 = 32'd3966
; 
32'd182959: dataIn1 = 32'd3984
; 
32'd182960: dataIn1 = 32'd5880
; 
32'd182961: dataIn1 = 32'd9273
; 
32'd182962: dataIn1 = 32'd9320
; 
32'd182963: dataIn1 = 32'd2743
; 
32'd182964: dataIn1 = 32'd5277
; 
32'd182965: dataIn1 = 32'd9278
; 
32'd182966: dataIn1 = 32'd9279
; 
32'd182967: dataIn1 = 32'd9321
; 
32'd182968: dataIn1 = 32'd9338
; 
32'd182969: dataIn1 = 32'd1124
; 
32'd182970: dataIn1 = 32'd5277
; 
32'd182971: dataIn1 = 32'd6751
; 
32'd182972: dataIn1 = 32'd9280
; 
32'd182973: dataIn1 = 32'd9322
; 
32'd182974: dataIn1 = 32'd9337
; 
32'd182975: dataIn1 = 32'd1139
; 
32'd182976: dataIn1 = 32'd5447
; 
32'd182977: dataIn1 = 32'd5448
; 
32'd182978: dataIn1 = 32'd6722
; 
32'd182979: dataIn1 = 32'd9282
; 
32'd182980: dataIn1 = 32'd9323
; 
32'd182981: dataIn1 = 32'd5436
; 
32'd182982: dataIn1 = 32'd5447
; 
32'd182983: dataIn1 = 32'd5516
; 
32'd182984: dataIn1 = 32'd9281
; 
32'd182985: dataIn1 = 32'd9294
; 
32'd182986: dataIn1 = 32'd9324
; 
32'd182987: dataIn1 = 32'd5451
; 
32'd182988: dataIn1 = 32'd5452
; 
32'd182989: dataIn1 = 32'd6729
; 
32'd182990: dataIn1 = 32'd9284
; 
32'd182991: dataIn1 = 32'd9325
; 
32'd182992: dataIn1 = 32'd10277
; 
32'd182993: dataIn1 = 32'd10281
; 
32'd182994: dataIn1 = 32'd5441
; 
32'd182995: dataIn1 = 32'd5452
; 
32'd182996: dataIn1 = 32'd5523
; 
32'd182997: dataIn1 = 32'd9283
; 
32'd182998: dataIn1 = 32'd9301
; 
32'd182999: dataIn1 = 32'd9326
; 
32'd183000: dataIn1 = 32'd5434
; 
32'd183001: dataIn1 = 32'd5445
; 
32'd183002: dataIn1 = 32'd5514
; 
32'd183003: dataIn1 = 32'd9288
; 
32'd183004: dataIn1 = 32'd9291
; 
32'd183005: dataIn1 = 32'd9327
; 
32'd183006: dataIn1 = 32'd17
; 
32'd183007: dataIn1 = 32'd5433
; 
32'd183008: dataIn1 = 32'd5434
; 
32'd183009: dataIn1 = 32'd9287
; 
32'd183010: dataIn1 = 32'd9290
; 
32'd183011: dataIn1 = 32'd9328
; 
32'd183012: dataIn1 = 32'd1138
; 
32'd183013: dataIn1 = 32'd5445
; 
32'd183014: dataIn1 = 32'd5446
; 
32'd183015: dataIn1 = 32'd9292
; 
32'd183016: dataIn1 = 32'd9298
; 
32'd183017: dataIn1 = 32'd9329
; 
32'd183018: dataIn1 = 32'd18
; 
32'd183019: dataIn1 = 32'd5435
; 
32'd183020: dataIn1 = 32'd5436
; 
32'd183021: dataIn1 = 32'd9293
; 
32'd183022: dataIn1 = 32'd9296
; 
32'd183023: dataIn1 = 32'd9330
; 
32'd183024: dataIn1 = 32'd5435
; 
32'd183025: dataIn1 = 32'd5446
; 
32'd183026: dataIn1 = 32'd5517
; 
32'd183027: dataIn1 = 32'd9295
; 
32'd183028: dataIn1 = 32'd9297
; 
32'd183029: dataIn1 = 32'd9331
; 
32'd183030: dataIn1 = 32'd5442
; 
32'd183031: dataIn1 = 32'd5453
; 
32'd183032: dataIn1 = 32'd5522
; 
32'd183033: dataIn1 = 32'd9300
; 
32'd183034: dataIn1 = 32'd9303
; 
32'd183035: dataIn1 = 32'd9332
; 
32'd183036: dataIn1 = 32'd21
; 
32'd183037: dataIn1 = 32'd5441
; 
32'd183038: dataIn1 = 32'd5442
; 
32'd183039: dataIn1 = 32'd9299
; 
32'd183040: dataIn1 = 32'd9302
; 
32'd183041: dataIn1 = 32'd9333
; 
32'd183042: dataIn1 = 32'd1142
; 
32'd183043: dataIn1 = 32'd5453
; 
32'd183044: dataIn1 = 32'd5454
; 
32'd183045: dataIn1 = 32'd9304
; 
32'd183046: dataIn1 = 32'd9310
; 
32'd183047: dataIn1 = 32'd9334
; 
32'd183048: dataIn1 = 32'd22
; 
32'd183049: dataIn1 = 32'd5443
; 
32'd183050: dataIn1 = 32'd5444
; 
32'd183051: dataIn1 = 32'd9305
; 
32'd183052: dataIn1 = 32'd9308
; 
32'd183053: dataIn1 = 32'd9335
; 
32'd183054: dataIn1 = 32'd5443
; 
32'd183055: dataIn1 = 32'd5454
; 
32'd183056: dataIn1 = 32'd5524
; 
32'd183057: dataIn1 = 32'd9307
; 
32'd183058: dataIn1 = 32'd9309
; 
32'd183059: dataIn1 = 32'd9336
; 
32'd183060: dataIn1 = 32'd1124
; 
32'd183061: dataIn1 = 32'd2745
; 
32'd183062: dataIn1 = 32'd5277
; 
32'd183063: dataIn1 = 32'd9289
; 
32'd183064: dataIn1 = 32'd9322
; 
32'd183065: dataIn1 = 32'd9337
; 
32'd183066: dataIn1 = 32'd9338
; 
32'd183067: dataIn1 = 32'd9339
; 
32'd183068: dataIn1 = 32'd2743
; 
32'd183069: dataIn1 = 32'd2744
; 
32'd183070: dataIn1 = 32'd2745
; 
32'd183071: dataIn1 = 32'd5277
; 
32'd183072: dataIn1 = 32'd9321
; 
32'd183073: dataIn1 = 32'd9337
; 
32'd183074: dataIn1 = 32'd9338
; 
32'd183075: dataIn1 = 32'd2745
; 
32'd183076: dataIn1 = 32'd5433
; 
32'd183077: dataIn1 = 32'd5515
; 
32'd183078: dataIn1 = 32'd9289
; 
32'd183079: dataIn1 = 32'd9337
; 
32'd183080: dataIn1 = 32'd9339
; 
32'd183081: dataIn1 = 32'd6803
; 
32'd183082: dataIn1 = 32'd6804
; 
32'd183083: dataIn1 = 32'd9340
; 
32'd183084: dataIn1 = 32'd9341
; 
32'd183085: dataIn1 = 32'd9342
; 
32'd183086: dataIn1 = 32'd9343
; 
32'd183087: dataIn1 = 32'd9344
; 
32'd183088: dataIn1 = 32'd6802
; 
32'd183089: dataIn1 = 32'd6804
; 
32'd183090: dataIn1 = 32'd9340
; 
32'd183091: dataIn1 = 32'd9341
; 
32'd183092: dataIn1 = 32'd9342
; 
32'd183093: dataIn1 = 32'd9345
; 
32'd183094: dataIn1 = 32'd9346
; 
32'd183095: dataIn1 = 32'd6802
; 
32'd183096: dataIn1 = 32'd6803
; 
32'd183097: dataIn1 = 32'd9340
; 
32'd183098: dataIn1 = 32'd9341
; 
32'd183099: dataIn1 = 32'd9342
; 
32'd183100: dataIn1 = 32'd9347
; 
32'd183101: dataIn1 = 32'd9348
; 
32'd183102: dataIn1 = 32'd5635
; 
32'd183103: dataIn1 = 32'd6804
; 
32'd183104: dataIn1 = 32'd9340
; 
32'd183105: dataIn1 = 32'd9343
; 
32'd183106: dataIn1 = 32'd9344
; 
32'd183107: dataIn1 = 32'd9356
; 
32'd183108: dataIn1 = 32'd9359
; 
32'd183109: dataIn1 = 32'd5635
; 
32'd183110: dataIn1 = 32'd6803
; 
32'd183111: dataIn1 = 32'd9340
; 
32'd183112: dataIn1 = 32'd9343
; 
32'd183113: dataIn1 = 32'd9344
; 
32'd183114: dataIn1 = 32'd9349
; 
32'd183115: dataIn1 = 32'd9352
; 
32'd183116: dataIn1 = 32'd5636
; 
32'd183117: dataIn1 = 32'd6804
; 
32'd183118: dataIn1 = 32'd9341
; 
32'd183119: dataIn1 = 32'd9345
; 
32'd183120: dataIn1 = 32'd9346
; 
32'd183121: dataIn1 = 32'd9357
; 
32'd183122: dataIn1 = 32'd9360
; 
32'd183123: dataIn1 = 32'd5636
; 
32'd183124: dataIn1 = 32'd6802
; 
32'd183125: dataIn1 = 32'd6805
; 
32'd183126: dataIn1 = 32'd6806
; 
32'd183127: dataIn1 = 32'd9341
; 
32'd183128: dataIn1 = 32'd9345
; 
32'd183129: dataIn1 = 32'd9346
; 
32'd183130: dataIn1 = 32'd5637
; 
32'd183131: dataIn1 = 32'd6803
; 
32'd183132: dataIn1 = 32'd9342
; 
32'd183133: dataIn1 = 32'd9347
; 
32'd183134: dataIn1 = 32'd9348
; 
32'd183135: dataIn1 = 32'd9351
; 
32'd183136: dataIn1 = 32'd9355
; 
32'd183137: dataIn1 = 32'd5637
; 
32'd183138: dataIn1 = 32'd6802
; 
32'd183139: dataIn1 = 32'd6805
; 
32'd183140: dataIn1 = 32'd6821
; 
32'd183141: dataIn1 = 32'd9342
; 
32'd183142: dataIn1 = 32'd9347
; 
32'd183143: dataIn1 = 32'd9348
; 
32'd183144: dataIn1 = 32'd6803
; 
32'd183145: dataIn1 = 32'd6808
; 
32'd183146: dataIn1 = 32'd9344
; 
32'd183147: dataIn1 = 32'd9349
; 
32'd183148: dataIn1 = 32'd9350
; 
32'd183149: dataIn1 = 32'd9351
; 
32'd183150: dataIn1 = 32'd9352
; 
32'd183151: dataIn1 = 32'd6807
; 
32'd183152: dataIn1 = 32'd6808
; 
32'd183153: dataIn1 = 32'd9349
; 
32'd183154: dataIn1 = 32'd9350
; 
32'd183155: dataIn1 = 32'd9351
; 
32'd183156: dataIn1 = 32'd9353
; 
32'd183157: dataIn1 = 32'd9354
; 
32'd183158: dataIn1 = 32'd6803
; 
32'd183159: dataIn1 = 32'd6807
; 
32'd183160: dataIn1 = 32'd9347
; 
32'd183161: dataIn1 = 32'd9349
; 
32'd183162: dataIn1 = 32'd9350
; 
32'd183163: dataIn1 = 32'd9351
; 
32'd183164: dataIn1 = 32'd9355
; 
32'd183165: dataIn1 = 32'd5635
; 
32'd183166: dataIn1 = 32'd6808
; 
32'd183167: dataIn1 = 32'd9344
; 
32'd183168: dataIn1 = 32'd9349
; 
32'd183169: dataIn1 = 32'd9352
; 
32'd183170: dataIn1 = 32'd9367
; 
32'd183171: dataIn1 = 32'd9372
; 
32'd183172: dataIn1 = 32'd3584
; 
32'd183173: dataIn1 = 32'd6808
; 
32'd183174: dataIn1 = 32'd9350
; 
32'd183175: dataIn1 = 32'd9353
; 
32'd183176: dataIn1 = 32'd9354
; 
32'd183177: dataIn1 = 32'd9373
; 
32'd183178: dataIn1 = 32'd9375
; 
32'd183179: dataIn1 = 32'd3584
; 
32'd183180: dataIn1 = 32'd6807
; 
32'd183181: dataIn1 = 32'd9350
; 
32'd183182: dataIn1 = 32'd9353
; 
32'd183183: dataIn1 = 32'd9354
; 
32'd183184: dataIn1 = 32'd9385
; 
32'd183185: dataIn1 = 32'd9389
; 
32'd183186: dataIn1 = 32'd5637
; 
32'd183187: dataIn1 = 32'd6807
; 
32'd183188: dataIn1 = 32'd9347
; 
32'd183189: dataIn1 = 32'd9351
; 
32'd183190: dataIn1 = 32'd9355
; 
32'd183191: dataIn1 = 32'd9386
; 
32'd183192: dataIn1 = 32'd9390
; 
32'd183193: dataIn1 = 32'd6804
; 
32'd183194: dataIn1 = 32'd6810
; 
32'd183195: dataIn1 = 32'd9343
; 
32'd183196: dataIn1 = 32'd9356
; 
32'd183197: dataIn1 = 32'd9357
; 
32'd183198: dataIn1 = 32'd9358
; 
32'd183199: dataIn1 = 32'd9359
; 
32'd183200: dataIn1 = 32'd6804
; 
32'd183201: dataIn1 = 32'd6809
; 
32'd183202: dataIn1 = 32'd9345
; 
32'd183203: dataIn1 = 32'd9356
; 
32'd183204: dataIn1 = 32'd9357
; 
32'd183205: dataIn1 = 32'd9358
; 
32'd183206: dataIn1 = 32'd9360
; 
32'd183207: dataIn1 = 32'd6809
; 
32'd183208: dataIn1 = 32'd6810
; 
32'd183209: dataIn1 = 32'd9356
; 
32'd183210: dataIn1 = 32'd9357
; 
32'd183211: dataIn1 = 32'd9358
; 
32'd183212: dataIn1 = 32'd9361
; 
32'd183213: dataIn1 = 32'd9362
; 
32'd183214: dataIn1 = 32'd5635
; 
32'd183215: dataIn1 = 32'd6810
; 
32'd183216: dataIn1 = 32'd9343
; 
32'd183217: dataIn1 = 32'd9356
; 
32'd183218: dataIn1 = 32'd9359
; 
32'd183219: dataIn1 = 32'd9366
; 
32'd183220: dataIn1 = 32'd9377
; 
32'd183221: dataIn1 = 32'd5636
; 
32'd183222: dataIn1 = 32'd6809
; 
32'd183223: dataIn1 = 32'd9345
; 
32'd183224: dataIn1 = 32'd9357
; 
32'd183225: dataIn1 = 32'd9360
; 
32'd183226: dataIn1 = 32'd9381
; 
32'd183227: dataIn1 = 32'd9383
; 
32'd183228: dataIn1 = 32'd2695
; 
32'd183229: dataIn1 = 32'd6810
; 
32'd183230: dataIn1 = 32'd7138
; 
32'd183231: dataIn1 = 32'd9358
; 
32'd183232: dataIn1 = 32'd9361
; 
32'd183233: dataIn1 = 32'd9362
; 
32'd183234: dataIn1 = 32'd9379
; 
32'd183235: dataIn1 = 32'd2695
; 
32'd183236: dataIn1 = 32'd6809
; 
32'd183237: dataIn1 = 32'd7162
; 
32'd183238: dataIn1 = 32'd9358
; 
32'd183239: dataIn1 = 32'd9361
; 
32'd183240: dataIn1 = 32'd9362
; 
32'd183241: dataIn1 = 32'd9382
; 
32'd183242: dataIn1 = 32'd6812
; 
32'd183243: dataIn1 = 32'd6813
; 
32'd183244: dataIn1 = 32'd9363
; 
32'd183245: dataIn1 = 32'd9364
; 
32'd183246: dataIn1 = 32'd9365
; 
32'd183247: dataIn1 = 32'd9366
; 
32'd183248: dataIn1 = 32'd9367
; 
32'd183249: dataIn1 = 32'd6811
; 
32'd183250: dataIn1 = 32'd6813
; 
32'd183251: dataIn1 = 32'd9363
; 
32'd183252: dataIn1 = 32'd9364
; 
32'd183253: dataIn1 = 32'd9365
; 
32'd183254: dataIn1 = 32'd9368
; 
32'd183255: dataIn1 = 32'd9369
; 
32'd183256: dataIn1 = 32'd6811
; 
32'd183257: dataIn1 = 32'd6812
; 
32'd183258: dataIn1 = 32'd9363
; 
32'd183259: dataIn1 = 32'd9364
; 
32'd183260: dataIn1 = 32'd9365
; 
32'd183261: dataIn1 = 32'd9370
; 
32'd183262: dataIn1 = 32'd9371
; 
32'd183263: dataIn1 = 32'd5635
; 
32'd183264: dataIn1 = 32'd6813
; 
32'd183265: dataIn1 = 32'd9359
; 
32'd183266: dataIn1 = 32'd9363
; 
32'd183267: dataIn1 = 32'd9366
; 
32'd183268: dataIn1 = 32'd9367
; 
32'd183269: dataIn1 = 32'd9377
; 
32'd183270: dataIn1 = 32'd5635
; 
32'd183271: dataIn1 = 32'd6812
; 
32'd183272: dataIn1 = 32'd9352
; 
32'd183273: dataIn1 = 32'd9363
; 
32'd183274: dataIn1 = 32'd9366
; 
32'd183275: dataIn1 = 32'd9367
; 
32'd183276: dataIn1 = 32'd9372
; 
32'd183277: dataIn1 = 32'd5124
; 
32'd183278: dataIn1 = 32'd6813
; 
32'd183279: dataIn1 = 32'd7140
; 
32'd183280: dataIn1 = 32'd9364
; 
32'd183281: dataIn1 = 32'd9368
; 
32'd183282: dataIn1 = 32'd9369
; 
32'd183283: dataIn1 = 32'd9378
; 
32'd183284: dataIn1 = 32'd5124
; 
32'd183285: dataIn1 = 32'd6811
; 
32'd183286: dataIn1 = 32'd9364
; 
32'd183287: dataIn1 = 32'd9368
; 
32'd183288: dataIn1 = 32'd9369
; 
32'd183289: dataIn1 = 32'd9807
; 
32'd183290: dataIn1 = 32'd9808
; 
32'd183291: dataIn1 = 32'd5638
; 
32'd183292: dataIn1 = 32'd6812
; 
32'd183293: dataIn1 = 32'd9365
; 
32'd183294: dataIn1 = 32'd9370
; 
32'd183295: dataIn1 = 32'd9371
; 
32'd183296: dataIn1 = 32'd9374
; 
32'd183297: dataIn1 = 32'd9376
; 
32'd183298: dataIn1 = 32'd5638
; 
32'd183299: dataIn1 = 32'd6811
; 
32'd183300: dataIn1 = 32'd9365
; 
32'd183301: dataIn1 = 32'd9370
; 
32'd183302: dataIn1 = 32'd9371
; 
32'd183303: dataIn1 = 32'd9809
; 
32'd183304: dataIn1 = 32'd9810
; 
32'd183305: dataIn1 = 32'd6808
; 
32'd183306: dataIn1 = 32'd6812
; 
32'd183307: dataIn1 = 32'd9352
; 
32'd183308: dataIn1 = 32'd9367
; 
32'd183309: dataIn1 = 32'd9372
; 
32'd183310: dataIn1 = 32'd9373
; 
32'd183311: dataIn1 = 32'd9374
; 
32'd183312: dataIn1 = 32'd6808
; 
32'd183313: dataIn1 = 32'd6815
; 
32'd183314: dataIn1 = 32'd9353
; 
32'd183315: dataIn1 = 32'd9372
; 
32'd183316: dataIn1 = 32'd9373
; 
32'd183317: dataIn1 = 32'd9374
; 
32'd183318: dataIn1 = 32'd9375
; 
32'd183319: dataIn1 = 32'd6812
; 
32'd183320: dataIn1 = 32'd6815
; 
32'd183321: dataIn1 = 32'd9370
; 
32'd183322: dataIn1 = 32'd9372
; 
32'd183323: dataIn1 = 32'd9373
; 
32'd183324: dataIn1 = 32'd9374
; 
32'd183325: dataIn1 = 32'd9376
; 
32'd183326: dataIn1 = 32'd3584
; 
32'd183327: dataIn1 = 32'd6815
; 
32'd183328: dataIn1 = 32'd9353
; 
32'd183329: dataIn1 = 32'd9373
; 
32'd183330: dataIn1 = 32'd9375
; 
32'd183331: dataIn1 = 32'd5638
; 
32'd183332: dataIn1 = 32'd6815
; 
32'd183333: dataIn1 = 32'd9370
; 
32'd183334: dataIn1 = 32'd9374
; 
32'd183335: dataIn1 = 32'd9376
; 
32'd183336: dataIn1 = 32'd6810
; 
32'd183337: dataIn1 = 32'd6813
; 
32'd183338: dataIn1 = 32'd9359
; 
32'd183339: dataIn1 = 32'd9366
; 
32'd183340: dataIn1 = 32'd9377
; 
32'd183341: dataIn1 = 32'd9378
; 
32'd183342: dataIn1 = 32'd9379
; 
32'd183343: dataIn1 = 32'd6110
; 
32'd183344: dataIn1 = 32'd6813
; 
32'd183345: dataIn1 = 32'd7140
; 
32'd183346: dataIn1 = 32'd9368
; 
32'd183347: dataIn1 = 32'd9377
; 
32'd183348: dataIn1 = 32'd9378
; 
32'd183349: dataIn1 = 32'd9379
; 
32'd183350: dataIn1 = 32'd6110
; 
32'd183351: dataIn1 = 32'd6810
; 
32'd183352: dataIn1 = 32'd7138
; 
32'd183353: dataIn1 = 32'd9361
; 
32'd183354: dataIn1 = 32'd9377
; 
32'd183355: dataIn1 = 32'd9378
; 
32'd183356: dataIn1 = 32'd9379
; 
32'd183357: dataIn1 = 32'd6117
; 
32'd183358: dataIn1 = 32'd6818
; 
32'd183359: dataIn1 = 32'd7161
; 
32'd183360: dataIn1 = 32'd9380
; 
32'd183361: dataIn1 = 32'd9381
; 
32'd183362: dataIn1 = 32'd9382
; 
32'd183363: dataIn1 = 32'd9446
; 
32'd183364: dataIn1 = 32'd6809
; 
32'd183365: dataIn1 = 32'd6818
; 
32'd183366: dataIn1 = 32'd9360
; 
32'd183367: dataIn1 = 32'd9380
; 
32'd183368: dataIn1 = 32'd9381
; 
32'd183369: dataIn1 = 32'd9382
; 
32'd183370: dataIn1 = 32'd9383
; 
32'd183371: dataIn1 = 32'd6117
; 
32'd183372: dataIn1 = 32'd6809
; 
32'd183373: dataIn1 = 32'd7162
; 
32'd183374: dataIn1 = 32'd9362
; 
32'd183375: dataIn1 = 32'd9380
; 
32'd183376: dataIn1 = 32'd9381
; 
32'd183377: dataIn1 = 32'd9382
; 
32'd183378: dataIn1 = 32'd5636
; 
32'd183379: dataIn1 = 32'd6806
; 
32'd183380: dataIn1 = 32'd6816
; 
32'd183381: dataIn1 = 32'd6818
; 
32'd183382: dataIn1 = 32'd9360
; 
32'd183383: dataIn1 = 32'd9381
; 
32'd183384: dataIn1 = 32'd9383
; 
32'd183385: dataIn1 = 32'd6822
; 
32'd183386: dataIn1 = 32'd6825
; 
32'd183387: dataIn1 = 32'd9384
; 
32'd183388: dataIn1 = 32'd9385
; 
32'd183389: dataIn1 = 32'd9386
; 
32'd183390: dataIn1 = 32'd9387
; 
32'd183391: dataIn1 = 32'd9388
; 
32'd183392: dataIn1 = 32'd6807
; 
32'd183393: dataIn1 = 32'd6825
; 
32'd183394: dataIn1 = 32'd9354
; 
32'd183395: dataIn1 = 32'd9384
; 
32'd183396: dataIn1 = 32'd9385
; 
32'd183397: dataIn1 = 32'd9386
; 
32'd183398: dataIn1 = 32'd9389
; 
32'd183399: dataIn1 = 32'd6807
; 
32'd183400: dataIn1 = 32'd6822
; 
32'd183401: dataIn1 = 32'd9355
; 
32'd183402: dataIn1 = 32'd9384
; 
32'd183403: dataIn1 = 32'd9385
; 
32'd183404: dataIn1 = 32'd9386
; 
32'd183405: dataIn1 = 32'd9390
; 
32'd183406: dataIn1 = 32'd5640
; 
32'd183407: dataIn1 = 32'd6825
; 
32'd183408: dataIn1 = 32'd9384
; 
32'd183409: dataIn1 = 32'd9387
; 
32'd183410: dataIn1 = 32'd9388
; 
32'd183411: dataIn1 = 32'd5640
; 
32'd183412: dataIn1 = 32'd6822
; 
32'd183413: dataIn1 = 32'd6823
; 
32'd183414: dataIn1 = 32'd6827
; 
32'd183415: dataIn1 = 32'd9384
; 
32'd183416: dataIn1 = 32'd9387
; 
32'd183417: dataIn1 = 32'd9388
; 
32'd183418: dataIn1 = 32'd3584
; 
32'd183419: dataIn1 = 32'd6825
; 
32'd183420: dataIn1 = 32'd9354
; 
32'd183421: dataIn1 = 32'd9385
; 
32'd183422: dataIn1 = 32'd9389
; 
32'd183423: dataIn1 = 32'd5637
; 
32'd183424: dataIn1 = 32'd6821
; 
32'd183425: dataIn1 = 32'd6822
; 
32'd183426: dataIn1 = 32'd6823
; 
32'd183427: dataIn1 = 32'd9355
; 
32'd183428: dataIn1 = 32'd9386
; 
32'd183429: dataIn1 = 32'd9390
; 
32'd183430: dataIn1 = 32'd6829
; 
32'd183431: dataIn1 = 32'd6830
; 
32'd183432: dataIn1 = 32'd9391
; 
32'd183433: dataIn1 = 32'd9392
; 
32'd183434: dataIn1 = 32'd9393
; 
32'd183435: dataIn1 = 32'd9394
; 
32'd183436: dataIn1 = 32'd9395
; 
32'd183437: dataIn1 = 32'd6828
; 
32'd183438: dataIn1 = 32'd6830
; 
32'd183439: dataIn1 = 32'd9391
; 
32'd183440: dataIn1 = 32'd9392
; 
32'd183441: dataIn1 = 32'd9393
; 
32'd183442: dataIn1 = 32'd9396
; 
32'd183443: dataIn1 = 32'd9397
; 
32'd183444: dataIn1 = 32'd6828
; 
32'd183445: dataIn1 = 32'd6829
; 
32'd183446: dataIn1 = 32'd9391
; 
32'd183447: dataIn1 = 32'd9392
; 
32'd183448: dataIn1 = 32'd9393
; 
32'd183449: dataIn1 = 32'd9398
; 
32'd183450: dataIn1 = 32'd9399
; 
32'd183451: dataIn1 = 32'd5642
; 
32'd183452: dataIn1 = 32'd6830
; 
32'd183453: dataIn1 = 32'd9391
; 
32'd183454: dataIn1 = 32'd9394
; 
32'd183455: dataIn1 = 32'd9395
; 
32'd183456: dataIn1 = 32'd9407
; 
32'd183457: dataIn1 = 32'd9410
; 
32'd183458: dataIn1 = 32'd5642
; 
32'd183459: dataIn1 = 32'd6829
; 
32'd183460: dataIn1 = 32'd9391
; 
32'd183461: dataIn1 = 32'd9394
; 
32'd183462: dataIn1 = 32'd9395
; 
32'd183463: dataIn1 = 32'd9400
; 
32'd183464: dataIn1 = 32'd9403
; 
32'd183465: dataIn1 = 32'd5643
; 
32'd183466: dataIn1 = 32'd6830
; 
32'd183467: dataIn1 = 32'd9392
; 
32'd183468: dataIn1 = 32'd9396
; 
32'd183469: dataIn1 = 32'd9397
; 
32'd183470: dataIn1 = 32'd9408
; 
32'd183471: dataIn1 = 32'd9411
; 
32'd183472: dataIn1 = 32'd5643
; 
32'd183473: dataIn1 = 32'd6828
; 
32'd183474: dataIn1 = 32'd6832
; 
32'd183475: dataIn1 = 32'd6842
; 
32'd183476: dataIn1 = 32'd9392
; 
32'd183477: dataIn1 = 32'd9396
; 
32'd183478: dataIn1 = 32'd9397
; 
32'd183479: dataIn1 = 32'd5644
; 
32'd183480: dataIn1 = 32'd6829
; 
32'd183481: dataIn1 = 32'd9393
; 
32'd183482: dataIn1 = 32'd9398
; 
32'd183483: dataIn1 = 32'd9399
; 
32'd183484: dataIn1 = 32'd9402
; 
32'd183485: dataIn1 = 32'd9406
; 
32'd183486: dataIn1 = 32'd5644
; 
32'd183487: dataIn1 = 32'd6828
; 
32'd183488: dataIn1 = 32'd6831
; 
32'd183489: dataIn1 = 32'd6832
; 
32'd183490: dataIn1 = 32'd9393
; 
32'd183491: dataIn1 = 32'd9398
; 
32'd183492: dataIn1 = 32'd9399
; 
32'd183493: dataIn1 = 32'd6829
; 
32'd183494: dataIn1 = 32'd6834
; 
32'd183495: dataIn1 = 32'd9395
; 
32'd183496: dataIn1 = 32'd9400
; 
32'd183497: dataIn1 = 32'd9401
; 
32'd183498: dataIn1 = 32'd9402
; 
32'd183499: dataIn1 = 32'd9403
; 
32'd183500: dataIn1 = 32'd6833
; 
32'd183501: dataIn1 = 32'd6834
; 
32'd183502: dataIn1 = 32'd9400
; 
32'd183503: dataIn1 = 32'd9401
; 
32'd183504: dataIn1 = 32'd9402
; 
32'd183505: dataIn1 = 32'd9404
; 
32'd183506: dataIn1 = 32'd9405
; 
32'd183507: dataIn1 = 32'd6829
; 
32'd183508: dataIn1 = 32'd6833
; 
32'd183509: dataIn1 = 32'd9398
; 
32'd183510: dataIn1 = 32'd9400
; 
32'd183511: dataIn1 = 32'd9401
; 
32'd183512: dataIn1 = 32'd9402
; 
32'd183513: dataIn1 = 32'd9406
; 
32'd183514: dataIn1 = 32'd5642
; 
32'd183515: dataIn1 = 32'd6834
; 
32'd183516: dataIn1 = 32'd9395
; 
32'd183517: dataIn1 = 32'd9400
; 
32'd183518: dataIn1 = 32'd9403
; 
32'd183519: dataIn1 = 32'd9418
; 
32'd183520: dataIn1 = 32'd9427
; 
32'd183521: dataIn1 = 32'd2733
; 
32'd183522: dataIn1 = 32'd6834
; 
32'd183523: dataIn1 = 32'd8862
; 
32'd183524: dataIn1 = 32'd9401
; 
32'd183525: dataIn1 = 32'd9404
; 
32'd183526: dataIn1 = 32'd9405
; 
32'd183527: dataIn1 = 32'd9428
; 
32'd183528: dataIn1 = 32'd2733
; 
32'd183529: dataIn1 = 32'd6833
; 
32'd183530: dataIn1 = 32'd9276
; 
32'd183531: dataIn1 = 32'd9401
; 
32'd183532: dataIn1 = 32'd9404
; 
32'd183533: dataIn1 = 32'd9405
; 
32'd183534: dataIn1 = 32'd9443
; 
32'd183535: dataIn1 = 32'd5644
; 
32'd183536: dataIn1 = 32'd6833
; 
32'd183537: dataIn1 = 32'd9398
; 
32'd183538: dataIn1 = 32'd9402
; 
32'd183539: dataIn1 = 32'd9406
; 
32'd183540: dataIn1 = 32'd9444
; 
32'd183541: dataIn1 = 32'd9445
; 
32'd183542: dataIn1 = 32'd6830
; 
32'd183543: dataIn1 = 32'd6836
; 
32'd183544: dataIn1 = 32'd9394
; 
32'd183545: dataIn1 = 32'd9407
; 
32'd183546: dataIn1 = 32'd9408
; 
32'd183547: dataIn1 = 32'd9409
; 
32'd183548: dataIn1 = 32'd9410
; 
32'd183549: dataIn1 = 32'd6830
; 
32'd183550: dataIn1 = 32'd6835
; 
32'd183551: dataIn1 = 32'd9396
; 
32'd183552: dataIn1 = 32'd9407
; 
32'd183553: dataIn1 = 32'd9408
; 
32'd183554: dataIn1 = 32'd9409
; 
32'd183555: dataIn1 = 32'd9411
; 
32'd183556: dataIn1 = 32'd6835
; 
32'd183557: dataIn1 = 32'd6836
; 
32'd183558: dataIn1 = 32'd9407
; 
32'd183559: dataIn1 = 32'd9408
; 
32'd183560: dataIn1 = 32'd9409
; 
32'd183561: dataIn1 = 32'd9412
; 
32'd183562: dataIn1 = 32'd9413
; 
32'd183563: dataIn1 = 32'd5642
; 
32'd183564: dataIn1 = 32'd6836
; 
32'd183565: dataIn1 = 32'd9394
; 
32'd183566: dataIn1 = 32'd9407
; 
32'd183567: dataIn1 = 32'd9410
; 
32'd183568: dataIn1 = 32'd9417
; 
32'd183569: dataIn1 = 32'd9430
; 
32'd183570: dataIn1 = 32'd5643
; 
32'd183571: dataIn1 = 32'd6835
; 
32'd183572: dataIn1 = 32'd9396
; 
32'd183573: dataIn1 = 32'd9408
; 
32'd183574: dataIn1 = 32'd9411
; 
32'd183575: dataIn1 = 32'd9436
; 
32'd183576: dataIn1 = 32'd9440
; 
32'd183577: dataIn1 = 32'd3586
; 
32'd183578: dataIn1 = 32'd6836
; 
32'd183579: dataIn1 = 32'd9409
; 
32'd183580: dataIn1 = 32'd9412
; 
32'd183581: dataIn1 = 32'd9413
; 
32'd183582: dataIn1 = 32'd9432
; 
32'd183583: dataIn1 = 32'd9434
; 
32'd183584: dataIn1 = 32'd3586
; 
32'd183585: dataIn1 = 32'd6835
; 
32'd183586: dataIn1 = 32'd9409
; 
32'd183587: dataIn1 = 32'd9412
; 
32'd183588: dataIn1 = 32'd9413
; 
32'd183589: dataIn1 = 32'd9437
; 
32'd183590: dataIn1 = 32'd9441
; 
32'd183591: dataIn1 = 32'd6838
; 
32'd183592: dataIn1 = 32'd6839
; 
32'd183593: dataIn1 = 32'd9414
; 
32'd183594: dataIn1 = 32'd9415
; 
32'd183595: dataIn1 = 32'd9416
; 
32'd183596: dataIn1 = 32'd9417
; 
32'd183597: dataIn1 = 32'd9418
; 
32'd183598: dataIn1 = 32'd6837
; 
32'd183599: dataIn1 = 32'd6839
; 
32'd183600: dataIn1 = 32'd9414
; 
32'd183601: dataIn1 = 32'd9415
; 
32'd183602: dataIn1 = 32'd9416
; 
32'd183603: dataIn1 = 32'd9419
; 
32'd183604: dataIn1 = 32'd9420
; 
32'd183605: dataIn1 = 32'd6837
; 
32'd183606: dataIn1 = 32'd6838
; 
32'd183607: dataIn1 = 32'd9414
; 
32'd183608: dataIn1 = 32'd9415
; 
32'd183609: dataIn1 = 32'd9416
; 
32'd183610: dataIn1 = 32'd9421
; 
32'd183611: dataIn1 = 32'd9422
; 
32'd183612: dataIn1 = 32'd5642
; 
32'd183613: dataIn1 = 32'd6839
; 
32'd183614: dataIn1 = 32'd9410
; 
32'd183615: dataIn1 = 32'd9414
; 
32'd183616: dataIn1 = 32'd9417
; 
32'd183617: dataIn1 = 32'd9418
; 
32'd183618: dataIn1 = 32'd9430
; 
32'd183619: dataIn1 = 32'd5642
; 
32'd183620: dataIn1 = 32'd6838
; 
32'd183621: dataIn1 = 32'd9403
; 
32'd183622: dataIn1 = 32'd9414
; 
32'd183623: dataIn1 = 32'd9417
; 
32'd183624: dataIn1 = 32'd9418
; 
32'd183625: dataIn1 = 32'd9427
; 
32'd183626: dataIn1 = 32'd5645
; 
32'd183627: dataIn1 = 32'd6839
; 
32'd183628: dataIn1 = 32'd9415
; 
32'd183629: dataIn1 = 32'd9419
; 
32'd183630: dataIn1 = 32'd9420
; 
32'd183631: dataIn1 = 32'd9431
; 
32'd183632: dataIn1 = 32'd9433
; 
32'd183633: dataIn1 = 32'd5645
; 
32'd183634: dataIn1 = 32'd6837
; 
32'd183635: dataIn1 = 32'd9415
; 
32'd183636: dataIn1 = 32'd9419
; 
32'd183637: dataIn1 = 32'd9420
; 
32'd183638: dataIn1 = 32'd9424
; 
32'd183639: dataIn1 = 32'd9426
; 
32'd183640: dataIn1 = 32'd5263
; 
32'd183641: dataIn1 = 32'd6838
; 
32'd183642: dataIn1 = 32'd8861
; 
32'd183643: dataIn1 = 32'd9416
; 
32'd183644: dataIn1 = 32'd9421
; 
32'd183645: dataIn1 = 32'd9422
; 
32'd183646: dataIn1 = 32'd9429
; 
32'd183647: dataIn1 = 32'd5263
; 
32'd183648: dataIn1 = 32'd6837
; 
32'd183649: dataIn1 = 32'd8866
; 
32'd183650: dataIn1 = 32'd9416
; 
32'd183651: dataIn1 = 32'd9421
; 
32'd183652: dataIn1 = 32'd9422
; 
32'd183653: dataIn1 = 32'd9425
; 
32'd183654: dataIn1 = 32'd6572
; 
32'd183655: dataIn1 = 32'd6840
; 
32'd183656: dataIn1 = 32'd8868
; 
32'd183657: dataIn1 = 32'd9423
; 
32'd183658: dataIn1 = 32'd9424
; 
32'd183659: dataIn1 = 32'd9425
; 
32'd183660: dataIn1 = 32'd9448
; 
32'd183661: dataIn1 = 32'd6837
; 
32'd183662: dataIn1 = 32'd6840
; 
32'd183663: dataIn1 = 32'd9420
; 
32'd183664: dataIn1 = 32'd9423
; 
32'd183665: dataIn1 = 32'd9424
; 
32'd183666: dataIn1 = 32'd9425
; 
32'd183667: dataIn1 = 32'd9426
; 
32'd183668: dataIn1 = 32'd6572
; 
32'd183669: dataIn1 = 32'd6837
; 
32'd183670: dataIn1 = 32'd8866
; 
32'd183671: dataIn1 = 32'd9422
; 
32'd183672: dataIn1 = 32'd9423
; 
32'd183673: dataIn1 = 32'd9424
; 
32'd183674: dataIn1 = 32'd9425
; 
32'd183675: dataIn1 = 32'd5645
; 
32'd183676: dataIn1 = 32'd6840
; 
32'd183677: dataIn1 = 32'd9420
; 
32'd183678: dataIn1 = 32'd9424
; 
32'd183679: dataIn1 = 32'd9426
; 
32'd183680: dataIn1 = 32'd6834
; 
32'd183681: dataIn1 = 32'd6838
; 
32'd183682: dataIn1 = 32'd9403
; 
32'd183683: dataIn1 = 32'd9418
; 
32'd183684: dataIn1 = 32'd9427
; 
32'd183685: dataIn1 = 32'd9428
; 
32'd183686: dataIn1 = 32'd9429
; 
32'd183687: dataIn1 = 32'd6571
; 
32'd183688: dataIn1 = 32'd6834
; 
32'd183689: dataIn1 = 32'd8862
; 
32'd183690: dataIn1 = 32'd9404
; 
32'd183691: dataIn1 = 32'd9427
; 
32'd183692: dataIn1 = 32'd9428
; 
32'd183693: dataIn1 = 32'd9429
; 
32'd183694: dataIn1 = 32'd6571
; 
32'd183695: dataIn1 = 32'd6838
; 
32'd183696: dataIn1 = 32'd8861
; 
32'd183697: dataIn1 = 32'd9421
; 
32'd183698: dataIn1 = 32'd9427
; 
32'd183699: dataIn1 = 32'd9428
; 
32'd183700: dataIn1 = 32'd9429
; 
32'd183701: dataIn1 = 32'd6836
; 
32'd183702: dataIn1 = 32'd6839
; 
32'd183703: dataIn1 = 32'd9410
; 
32'd183704: dataIn1 = 32'd9417
; 
32'd183705: dataIn1 = 32'd9430
; 
32'd183706: dataIn1 = 32'd9431
; 
32'd183707: dataIn1 = 32'd9432
; 
32'd183708: dataIn1 = 32'd6839
; 
32'd183709: dataIn1 = 32'd6841
; 
32'd183710: dataIn1 = 32'd9419
; 
32'd183711: dataIn1 = 32'd9430
; 
32'd183712: dataIn1 = 32'd9431
; 
32'd183713: dataIn1 = 32'd9432
; 
32'd183714: dataIn1 = 32'd9433
; 
32'd183715: dataIn1 = 32'd6836
; 
32'd183716: dataIn1 = 32'd6841
; 
32'd183717: dataIn1 = 32'd9412
; 
32'd183718: dataIn1 = 32'd9430
; 
32'd183719: dataIn1 = 32'd9431
; 
32'd183720: dataIn1 = 32'd9432
; 
32'd183721: dataIn1 = 32'd9434
; 
32'd183722: dataIn1 = 32'd5645
; 
32'd183723: dataIn1 = 32'd6841
; 
32'd183724: dataIn1 = 32'd9419
; 
32'd183725: dataIn1 = 32'd9431
; 
32'd183726: dataIn1 = 32'd9433
; 
32'd183727: dataIn1 = 32'd3586
; 
32'd183728: dataIn1 = 32'd6841
; 
32'd183729: dataIn1 = 32'd9412
; 
32'd183730: dataIn1 = 32'd9432
; 
32'd183731: dataIn1 = 32'd9434
; 
32'd183732: dataIn1 = 32'd6844
; 
32'd183733: dataIn1 = 32'd6846
; 
32'd183734: dataIn1 = 32'd9435
; 
32'd183735: dataIn1 = 32'd9436
; 
32'd183736: dataIn1 = 32'd9437
; 
32'd183737: dataIn1 = 32'd9438
; 
32'd183738: dataIn1 = 32'd9439
; 
32'd183739: dataIn1 = 32'd6835
; 
32'd183740: dataIn1 = 32'd6844
; 
32'd183741: dataIn1 = 32'd9411
; 
32'd183742: dataIn1 = 32'd9435
; 
32'd183743: dataIn1 = 32'd9436
; 
32'd183744: dataIn1 = 32'd9437
; 
32'd183745: dataIn1 = 32'd9440
; 
32'd183746: dataIn1 = 32'd6835
; 
32'd183747: dataIn1 = 32'd6846
; 
32'd183748: dataIn1 = 32'd9413
; 
32'd183749: dataIn1 = 32'd9435
; 
32'd183750: dataIn1 = 32'd9436
; 
32'd183751: dataIn1 = 32'd9437
; 
32'd183752: dataIn1 = 32'd9441
; 
32'd183753: dataIn1 = 32'd5646
; 
32'd183754: dataIn1 = 32'd6843
; 
32'd183755: dataIn1 = 32'd6844
; 
32'd183756: dataIn1 = 32'd9435
; 
32'd183757: dataIn1 = 32'd9438
; 
32'd183758: dataIn1 = 32'd9439
; 
32'd183759: dataIn1 = 32'd10291
; 
32'd183760: dataIn1 = 32'd5646
; 
32'd183761: dataIn1 = 32'd6846
; 
32'd183762: dataIn1 = 32'd9435
; 
32'd183763: dataIn1 = 32'd9438
; 
32'd183764: dataIn1 = 32'd9439
; 
32'd183765: dataIn1 = 32'd5643
; 
32'd183766: dataIn1 = 32'd6842
; 
32'd183767: dataIn1 = 32'd6843
; 
32'd183768: dataIn1 = 32'd6844
; 
32'd183769: dataIn1 = 32'd9411
; 
32'd183770: dataIn1 = 32'd9436
; 
32'd183771: dataIn1 = 32'd9440
; 
32'd183772: dataIn1 = 32'd3586
; 
32'd183773: dataIn1 = 32'd6846
; 
32'd183774: dataIn1 = 32'd9413
; 
32'd183775: dataIn1 = 32'd9437
; 
32'd183776: dataIn1 = 32'd9441
; 
32'd183777: dataIn1 = 32'd6564
; 
32'd183778: dataIn1 = 32'd6848
; 
32'd183779: dataIn1 = 32'd8818
; 
32'd183780: dataIn1 = 32'd9442
; 
32'd183781: dataIn1 = 32'd9443
; 
32'd183782: dataIn1 = 32'd9444
; 
32'd183783: dataIn1 = 32'd9447
; 
32'd183784: dataIn1 = 32'd6564
; 
32'd183785: dataIn1 = 32'd6833
; 
32'd183786: dataIn1 = 32'd9276
; 
32'd183787: dataIn1 = 32'd9405
; 
32'd183788: dataIn1 = 32'd9442
; 
32'd183789: dataIn1 = 32'd9443
; 
32'd183790: dataIn1 = 32'd9444
; 
32'd183791: dataIn1 = 32'd6833
; 
32'd183792: dataIn1 = 32'd6848
; 
32'd183793: dataIn1 = 32'd9406
; 
32'd183794: dataIn1 = 32'd9442
; 
32'd183795: dataIn1 = 32'd9443
; 
32'd183796: dataIn1 = 32'd9444
; 
32'd183797: dataIn1 = 32'd9445
; 
32'd183798: dataIn1 = 32'd5644
; 
32'd183799: dataIn1 = 32'd6831
; 
32'd183800: dataIn1 = 32'd6847
; 
32'd183801: dataIn1 = 32'd6848
; 
32'd183802: dataIn1 = 32'd9406
; 
32'd183803: dataIn1 = 32'd9444
; 
32'd183804: dataIn1 = 32'd9445
; 
32'd183805: dataIn1 = 32'd5125
; 
32'd183806: dataIn1 = 32'd6816
; 
32'd183807: dataIn1 = 32'd6817
; 
32'd183808: dataIn1 = 32'd6818
; 
32'd183809: dataIn1 = 32'd7161
; 
32'd183810: dataIn1 = 32'd9380
; 
32'd183811: dataIn1 = 32'd9446
; 
32'd183812: dataIn1 = 32'd5262
; 
32'd183813: dataIn1 = 32'd6847
; 
32'd183814: dataIn1 = 32'd6848
; 
32'd183815: dataIn1 = 32'd6849
; 
32'd183816: dataIn1 = 32'd8818
; 
32'd183817: dataIn1 = 32'd9442
; 
32'd183818: dataIn1 = 32'd9447
; 
32'd183819: dataIn1 = 32'd12
; 
32'd183820: dataIn1 = 32'd6840
; 
32'd183821: dataIn1 = 32'd8868
; 
32'd183822: dataIn1 = 32'd9423
; 
32'd183823: dataIn1 = 32'd9448
; 
32'd183824: dataIn1 = 32'd2112
; 
32'd183825: dataIn1 = 32'd9449
; 
32'd183826: dataIn1 = 32'd9450
; 
32'd183827: dataIn1 = 32'd9452
; 
32'd183828: dataIn1 = 32'd9812
; 
32'd183829: dataIn1 = 32'd9813
; 
32'd183830: dataIn1 = 32'd9815
; 
32'd183831: dataIn1 = 32'd30
; 
32'd183832: dataIn1 = 32'd2112
; 
32'd183833: dataIn1 = 32'd2113
; 
32'd183834: dataIn1 = 32'd9449
; 
32'd183835: dataIn1 = 32'd9450
; 
32'd183836: dataIn1 = 32'd9451
; 
32'd183837: dataIn1 = 32'd9812
; 
32'd183838: dataIn1 = 32'd9819
; 
32'd183839: dataIn1 = 32'd9450
; 
32'd183840: dataIn1 = 32'd9451
; 
32'd183841: dataIn1 = 32'd9811
; 
32'd183842: dataIn1 = 32'd9812
; 
32'd183843: dataIn1 = 32'd9816
; 
32'd183844: dataIn1 = 32'd9817
; 
32'd183845: dataIn1 = 32'd9819
; 
32'd183846: dataIn1 = 32'd20
; 
32'd183847: dataIn1 = 32'd2112
; 
32'd183848: dataIn1 = 32'd5521
; 
32'd183849: dataIn1 = 32'd9449
; 
32'd183850: dataIn1 = 32'd9452
; 
32'd183851: dataIn1 = 32'd9453
; 
32'd183852: dataIn1 = 32'd9676
; 
32'd183853: dataIn1 = 32'd9815
; 
32'd183854: dataIn1 = 32'd9825
; 
32'd183855: dataIn1 = 32'd9452
; 
32'd183856: dataIn1 = 32'd9453
; 
32'd183857: dataIn1 = 32'd9814
; 
32'd183858: dataIn1 = 32'd9815
; 
32'd183859: dataIn1 = 32'd9822
; 
32'd183860: dataIn1 = 32'd9824
; 
32'd183861: dataIn1 = 32'd9825
; 
32'd183862: dataIn1 = 32'd31
; 
32'd183863: dataIn1 = 32'd9454
; 
32'd183864: dataIn1 = 32'd9817
; 
32'd183865: dataIn1 = 32'd9818
; 
32'd183866: dataIn1 = 32'd9821
; 
32'd183867: dataIn1 = 32'd10152
; 
32'd183868: dataIn1 = 32'd10153
; 
32'd183869: dataIn1 = 32'd31
; 
32'd183870: dataIn1 = 32'd9455
; 
32'd183871: dataIn1 = 32'd9816
; 
32'd183872: dataIn1 = 32'd9818
; 
32'd183873: dataIn1 = 32'd9820
; 
32'd183874: dataIn1 = 32'd9828
; 
32'd183875: dataIn1 = 32'd9829
; 
32'd183876: dataIn1 = 32'd9456
; 
32'd183877: dataIn1 = 32'd9823
; 
32'd183878: dataIn1 = 32'd9824
; 
32'd183879: dataIn1 = 32'd9826
; 
32'd183880: dataIn1 = 32'd10152
; 
32'd183881: dataIn1 = 32'd10154
; 
32'd183882: dataIn1 = 32'd10283
; 
32'd183883: dataIn1 = 32'd31
; 
32'd183884: dataIn1 = 32'd9457
; 
32'd183885: dataIn1 = 32'd9462
; 
32'd183886: dataIn1 = 32'd9827
; 
32'd183887: dataIn1 = 32'd9829
; 
32'd183888: dataIn1 = 32'd9831
; 
32'd183889: dataIn1 = 32'd9836
; 
32'd183890: dataIn1 = 32'd9458
; 
32'd183891: dataIn1 = 32'd9827
; 
32'd183892: dataIn1 = 32'd9828
; 
32'd183893: dataIn1 = 32'd9830
; 
32'd183894: dataIn1 = 32'd9832
; 
32'd183895: dataIn1 = 32'd10155
; 
32'd183896: dataIn1 = 32'd10156
; 
32'd183897: dataIn1 = 32'd2149
; 
32'd183898: dataIn1 = 32'd9459
; 
32'd183899: dataIn1 = 32'd9461
; 
32'd183900: dataIn1 = 32'd9462
; 
32'd183901: dataIn1 = 32'd9834
; 
32'd183902: dataIn1 = 32'd9835
; 
32'd183903: dataIn1 = 32'd9836
; 
32'd183904: dataIn1 = 32'd9460
; 
32'd183905: dataIn1 = 32'd9461
; 
32'd183906: dataIn1 = 32'd9833
; 
32'd183907: dataIn1 = 32'd9835
; 
32'd183908: dataIn1 = 32'd9837
; 
32'd183909: dataIn1 = 32'd9839
; 
32'd183910: dataIn1 = 32'd9841
; 
32'd183911: dataIn1 = 32'd2148
; 
32'd183912: dataIn1 = 32'd2149
; 
32'd183913: dataIn1 = 32'd9459
; 
32'd183914: dataIn1 = 32'd9460
; 
32'd183915: dataIn1 = 32'd9461
; 
32'd183916: dataIn1 = 32'd9477
; 
32'd183917: dataIn1 = 32'd9769
; 
32'd183918: dataIn1 = 32'd9835
; 
32'd183919: dataIn1 = 32'd9841
; 
32'd183920: dataIn1 = 32'd31
; 
32'd183921: dataIn1 = 32'd2116
; 
32'd183922: dataIn1 = 32'd2149
; 
32'd183923: dataIn1 = 32'd9457
; 
32'd183924: dataIn1 = 32'd9459
; 
32'd183925: dataIn1 = 32'd9462
; 
32'd183926: dataIn1 = 32'd9836
; 
32'd183927: dataIn1 = 32'd41
; 
32'd183928: dataIn1 = 32'd9463
; 
32'd183929: dataIn1 = 32'd9838
; 
32'd183930: dataIn1 = 32'd9839
; 
32'd183931: dataIn1 = 32'd9842
; 
32'd183932: dataIn1 = 32'd10156
; 
32'd183933: dataIn1 = 32'd10157
; 
32'd183934: dataIn1 = 32'd41
; 
32'd183935: dataIn1 = 32'd9464
; 
32'd183936: dataIn1 = 32'd9837
; 
32'd183937: dataIn1 = 32'd9838
; 
32'd183938: dataIn1 = 32'd9840
; 
32'd183939: dataIn1 = 32'd9845
; 
32'd183940: dataIn1 = 32'd9846
; 
32'd183941: dataIn1 = 32'd9465
; 
32'd183942: dataIn1 = 32'd9466
; 
32'd183943: dataIn1 = 32'd9843
; 
32'd183944: dataIn1 = 32'd9844
; 
32'd183945: dataIn1 = 32'd9846
; 
32'd183946: dataIn1 = 32'd9847
; 
32'd183947: dataIn1 = 32'd9848
; 
32'd183948: dataIn1 = 32'd2148
; 
32'd183949: dataIn1 = 32'd2178
; 
32'd183950: dataIn1 = 32'd3590
; 
32'd183951: dataIn1 = 32'd3595
; 
32'd183952: dataIn1 = 32'd9465
; 
32'd183953: dataIn1 = 32'd9466
; 
32'd183954: dataIn1 = 32'd9477
; 
32'd183955: dataIn1 = 32'd9844
; 
32'd183956: dataIn1 = 32'd9848
; 
32'd183957: dataIn1 = 32'd41
; 
32'd183958: dataIn1 = 32'd9467
; 
32'd183959: dataIn1 = 32'd9781
; 
32'd183960: dataIn1 = 32'd9845
; 
32'd183961: dataIn1 = 32'd9847
; 
32'd183962: dataIn1 = 32'd9849
; 
32'd183963: dataIn1 = 32'd10227
; 
32'd183964: dataIn1 = 32'd9468
; 
32'd183965: dataIn1 = 32'd9471
; 
32'd183966: dataIn1 = 32'd9851
; 
32'd183967: dataIn1 = 32'd9852
; 
32'd183968: dataIn1 = 32'd9854
; 
32'd183969: dataIn1 = 32'd9856
; 
32'd183970: dataIn1 = 32'd9858
; 
32'd183971: dataIn1 = 32'd3587
; 
32'd183972: dataIn1 = 32'd9469
; 
32'd183973: dataIn1 = 32'd9850
; 
32'd183974: dataIn1 = 32'd9852
; 
32'd183975: dataIn1 = 32'd9855
; 
32'd183976: dataIn1 = 32'd9859
; 
32'd183977: dataIn1 = 32'd9861
; 
32'd183978: dataIn1 = 32'd3587
; 
32'd183979: dataIn1 = 32'd9470
; 
32'd183980: dataIn1 = 32'd9850
; 
32'd183981: dataIn1 = 32'd9851
; 
32'd183982: dataIn1 = 32'd9853
; 
32'd183983: dataIn1 = 32'd10158
; 
32'd183984: dataIn1 = 32'd10159
; 
32'd183985: dataIn1 = 32'd2176
; 
32'd183986: dataIn1 = 32'd3589
; 
32'd183987: dataIn1 = 32'd9468
; 
32'd183988: dataIn1 = 32'd9471
; 
32'd183989: dataIn1 = 32'd9472
; 
32'd183990: dataIn1 = 32'd9771
; 
32'd183991: dataIn1 = 32'd9856
; 
32'd183992: dataIn1 = 32'd9858
; 
32'd183993: dataIn1 = 32'd2176
; 
32'd183994: dataIn1 = 32'd9471
; 
32'd183995: dataIn1 = 32'd9472
; 
32'd183996: dataIn1 = 32'd9857
; 
32'd183997: dataIn1 = 32'd9858
; 
32'd183998: dataIn1 = 32'd9906
; 
32'd183999: dataIn1 = 32'd9907
; 
32'd184000: dataIn1 = 32'd9473
; 
32'd184001: dataIn1 = 32'd9860
; 
32'd184002: dataIn1 = 32'd9861
; 
32'd184003: dataIn1 = 32'd9863
; 
32'd184004: dataIn1 = 32'd9864
; 
32'd184005: dataIn1 = 32'd10160
; 
32'd184006: dataIn1 = 32'd10161
; 
32'd184007: dataIn1 = 32'd3587
; 
32'd184008: dataIn1 = 32'd9474
; 
32'd184009: dataIn1 = 32'd9476
; 
32'd184010: dataIn1 = 32'd9859
; 
32'd184011: dataIn1 = 32'd9860
; 
32'd184012: dataIn1 = 32'd9862
; 
32'd184013: dataIn1 = 32'd9866
; 
32'd184014: dataIn1 = 32'd3590
; 
32'd184015: dataIn1 = 32'd9475
; 
32'd184016: dataIn1 = 32'd9476
; 
32'd184017: dataIn1 = 32'd9843
; 
32'd184018: dataIn1 = 32'd9844
; 
32'd184019: dataIn1 = 32'd9865
; 
32'd184020: dataIn1 = 32'd9866
; 
32'd184021: dataIn1 = 32'd3587
; 
32'd184022: dataIn1 = 32'd3590
; 
32'd184023: dataIn1 = 32'd3591
; 
32'd184024: dataIn1 = 32'd9474
; 
32'd184025: dataIn1 = 32'd9475
; 
32'd184026: dataIn1 = 32'd9476
; 
32'd184027: dataIn1 = 32'd9866
; 
32'd184028: dataIn1 = 32'd42
; 
32'd184029: dataIn1 = 32'd2148
; 
32'd184030: dataIn1 = 32'd3595
; 
32'd184031: dataIn1 = 32'd9461
; 
32'd184032: dataIn1 = 32'd9466
; 
32'd184033: dataIn1 = 32'd9477
; 
32'd184034: dataIn1 = 32'd9769
; 
32'd184035: dataIn1 = 32'd9478
; 
32'd184036: dataIn1 = 32'd9480
; 
32'd184037: dataIn1 = 32'd9868
; 
32'd184038: dataIn1 = 32'd9869
; 
32'd184039: dataIn1 = 32'd9871
; 
32'd184040: dataIn1 = 32'd9872
; 
32'd184041: dataIn1 = 32'd9874
; 
32'd184042: dataIn1 = 32'd3620
; 
32'd184043: dataIn1 = 32'd9479
; 
32'd184044: dataIn1 = 32'd9480
; 
32'd184045: dataIn1 = 32'd9484
; 
32'd184046: dataIn1 = 32'd9867
; 
32'd184047: dataIn1 = 32'd9869
; 
32'd184048: dataIn1 = 32'd9877
; 
32'd184049: dataIn1 = 32'd2203
; 
32'd184050: dataIn1 = 32'd3620
; 
32'd184051: dataIn1 = 32'd3621
; 
32'd184052: dataIn1 = 32'd9478
; 
32'd184053: dataIn1 = 32'd9479
; 
32'd184054: dataIn1 = 32'd9480
; 
32'd184055: dataIn1 = 32'd9869
; 
32'd184056: dataIn1 = 32'd9874
; 
32'd184057: dataIn1 = 32'd2204
; 
32'd184058: dataIn1 = 32'd9481
; 
32'd184059: dataIn1 = 32'd9870
; 
32'd184060: dataIn1 = 32'd9872
; 
32'd184061: dataIn1 = 32'd9875
; 
32'd184062: dataIn1 = 32'd10162
; 
32'd184063: dataIn1 = 32'd10163
; 
32'd184064: dataIn1 = 32'd2204
; 
32'd184065: dataIn1 = 32'd9482
; 
32'd184066: dataIn1 = 32'd9870
; 
32'd184067: dataIn1 = 32'd9871
; 
32'd184068: dataIn1 = 32'd9873
; 
32'd184069: dataIn1 = 32'd9878
; 
32'd184070: dataIn1 = 32'd9879
; 
32'd184071: dataIn1 = 32'd9483
; 
32'd184072: dataIn1 = 32'd9484
; 
32'd184073: dataIn1 = 32'd9876
; 
32'd184074: dataIn1 = 32'd9877
; 
32'd184075: dataIn1 = 32'd9885
; 
32'd184076: dataIn1 = 32'd9886
; 
32'd184077: dataIn1 = 32'd9888
; 
32'd184078: dataIn1 = 32'd2205
; 
32'd184079: dataIn1 = 32'd3620
; 
32'd184080: dataIn1 = 32'd9479
; 
32'd184081: dataIn1 = 32'd9483
; 
32'd184082: dataIn1 = 32'd9484
; 
32'd184083: dataIn1 = 32'd9877
; 
32'd184084: dataIn1 = 32'd9888
; 
32'd184085: dataIn1 = 32'd10169
; 
32'd184086: dataIn1 = 32'd10229
; 
32'd184087: dataIn1 = 32'd9485
; 
32'd184088: dataIn1 = 32'd9879
; 
32'd184089: dataIn1 = 32'd9880
; 
32'd184090: dataIn1 = 32'd9881
; 
32'd184091: dataIn1 = 32'd9883
; 
32'd184092: dataIn1 = 32'd10164
; 
32'd184093: dataIn1 = 32'd10165
; 
32'd184094: dataIn1 = 32'd2204
; 
32'd184095: dataIn1 = 32'd9486
; 
32'd184096: dataIn1 = 32'd9557
; 
32'd184097: dataIn1 = 32'd9878
; 
32'd184098: dataIn1 = 32'd9880
; 
32'd184099: dataIn1 = 32'd9882
; 
32'd184100: dataIn1 = 32'd10026
; 
32'd184101: dataIn1 = 32'd3626
; 
32'd184102: dataIn1 = 32'd9487
; 
32'd184103: dataIn1 = 32'd9884
; 
32'd184104: dataIn1 = 32'd9886
; 
32'd184105: dataIn1 = 32'd9889
; 
32'd184106: dataIn1 = 32'd10162
; 
32'd184107: dataIn1 = 32'd10166
; 
32'd184108: dataIn1 = 32'd3626
; 
32'd184109: dataIn1 = 32'd9488
; 
32'd184110: dataIn1 = 32'd9496
; 
32'd184111: dataIn1 = 32'd9884
; 
32'd184112: dataIn1 = 32'd9885
; 
32'd184113: dataIn1 = 32'd9887
; 
32'd184114: dataIn1 = 32'd9905
; 
32'd184115: dataIn1 = 32'd3629
; 
32'd184116: dataIn1 = 32'd9489
; 
32'd184117: dataIn1 = 32'd9891
; 
32'd184118: dataIn1 = 32'd9892
; 
32'd184119: dataIn1 = 32'd9896
; 
32'd184120: dataIn1 = 32'd10167
; 
32'd184121: dataIn1 = 32'd10168
; 
32'd184122: dataIn1 = 32'd9490
; 
32'd184123: dataIn1 = 32'd9493
; 
32'd184124: dataIn1 = 32'd9890
; 
32'd184125: dataIn1 = 32'd9892
; 
32'd184126: dataIn1 = 32'd9894
; 
32'd184127: dataIn1 = 32'd9895
; 
32'd184128: dataIn1 = 32'd9898
; 
32'd184129: dataIn1 = 32'd3629
; 
32'd184130: dataIn1 = 32'd9491
; 
32'd184131: dataIn1 = 32'd9890
; 
32'd184132: dataIn1 = 32'd9891
; 
32'd184133: dataIn1 = 32'd9893
; 
32'd184134: dataIn1 = 32'd9899
; 
32'd184135: dataIn1 = 32'd9900
; 
32'd184136: dataIn1 = 32'd2176
; 
32'd184137: dataIn1 = 32'd9492
; 
32'd184138: dataIn1 = 32'd9493
; 
32'd184139: dataIn1 = 32'd9897
; 
32'd184140: dataIn1 = 32'd9898
; 
32'd184141: dataIn1 = 32'd9907
; 
32'd184142: dataIn1 = 32'd9908
; 
32'd184143: dataIn1 = 32'd2176
; 
32'd184144: dataIn1 = 32'd3628
; 
32'd184145: dataIn1 = 32'd3631
; 
32'd184146: dataIn1 = 32'd9490
; 
32'd184147: dataIn1 = 32'd9492
; 
32'd184148: dataIn1 = 32'd9493
; 
32'd184149: dataIn1 = 32'd9894
; 
32'd184150: dataIn1 = 32'd9898
; 
32'd184151: dataIn1 = 32'd3629
; 
32'd184152: dataIn1 = 32'd9494
; 
32'd184153: dataIn1 = 32'd9496
; 
32'd184154: dataIn1 = 32'd9900
; 
32'd184155: dataIn1 = 32'd9901
; 
32'd184156: dataIn1 = 32'd9904
; 
32'd184157: dataIn1 = 32'd9905
; 
32'd184158: dataIn1 = 32'd9495
; 
32'd184159: dataIn1 = 32'd9899
; 
32'd184160: dataIn1 = 32'd9901
; 
32'd184161: dataIn1 = 32'd9902
; 
32'd184162: dataIn1 = 32'd9903
; 
32'd184163: dataIn1 = 32'd10169
; 
32'd184164: dataIn1 = 32'd10170
; 
32'd184165: dataIn1 = 32'd3626
; 
32'd184166: dataIn1 = 32'd3629
; 
32'd184167: dataIn1 = 32'd3632
; 
32'd184168: dataIn1 = 32'd9488
; 
32'd184169: dataIn1 = 32'd9494
; 
32'd184170: dataIn1 = 32'd9496
; 
32'd184171: dataIn1 = 32'd9905
; 
32'd184172: dataIn1 = 32'd9497
; 
32'd184173: dataIn1 = 32'd9906
; 
32'd184174: dataIn1 = 32'd9908
; 
32'd184175: dataIn1 = 32'd9909
; 
32'd184176: dataIn1 = 32'd9910
; 
32'd184177: dataIn1 = 32'd10171
; 
32'd184178: dataIn1 = 32'd10172
; 
32'd184179: dataIn1 = 32'd3666
; 
32'd184180: dataIn1 = 32'd9498
; 
32'd184181: dataIn1 = 32'd9499
; 
32'd184182: dataIn1 = 32'd9501
; 
32'd184183: dataIn1 = 32'd9912
; 
32'd184184: dataIn1 = 32'd9913
; 
32'd184185: dataIn1 = 32'd9915
; 
32'd184186: dataIn1 = 32'd2224
; 
32'd184187: dataIn1 = 32'd3666
; 
32'd184188: dataIn1 = 32'd3668
; 
32'd184189: dataIn1 = 32'd9498
; 
32'd184190: dataIn1 = 32'd9499
; 
32'd184191: dataIn1 = 32'd9500
; 
32'd184192: dataIn1 = 32'd9912
; 
32'd184193: dataIn1 = 32'd3668
; 
32'd184194: dataIn1 = 32'd9499
; 
32'd184195: dataIn1 = 32'd9500
; 
32'd184196: dataIn1 = 32'd9911
; 
32'd184197: dataIn1 = 32'd9912
; 
32'd184198: dataIn1 = 32'd9916
; 
32'd184199: dataIn1 = 32'd9917
; 
32'd184200: dataIn1 = 32'd2223
; 
32'd184201: dataIn1 = 32'd3666
; 
32'd184202: dataIn1 = 32'd9498
; 
32'd184203: dataIn1 = 32'd9501
; 
32'd184204: dataIn1 = 32'd9502
; 
32'd184205: dataIn1 = 32'd9915
; 
32'd184206: dataIn1 = 32'd10118
; 
32'd184207: dataIn1 = 32'd10218
; 
32'd184208: dataIn1 = 32'd10245
; 
32'd184209: dataIn1 = 32'd9501
; 
32'd184210: dataIn1 = 32'd9502
; 
32'd184211: dataIn1 = 32'd9914
; 
32'd184212: dataIn1 = 32'd9915
; 
32'd184213: dataIn1 = 32'd10114
; 
32'd184214: dataIn1 = 32'd10115
; 
32'd184215: dataIn1 = 32'd10118
; 
32'd184216: dataIn1 = 32'd9503
; 
32'd184217: dataIn1 = 32'd9917
; 
32'd184218: dataIn1 = 32'd9918
; 
32'd184219: dataIn1 = 32'd9919
; 
32'd184220: dataIn1 = 32'd9921
; 
32'd184221: dataIn1 = 32'd10173
; 
32'd184222: dataIn1 = 32'd10174
; 
32'd184223: dataIn1 = 32'd3668
; 
32'd184224: dataIn1 = 32'd9504
; 
32'd184225: dataIn1 = 32'd9506
; 
32'd184226: dataIn1 = 32'd9916
; 
32'd184227: dataIn1 = 32'd9918
; 
32'd184228: dataIn1 = 32'd9920
; 
32'd184229: dataIn1 = 32'd9922
; 
32'd184230: dataIn1 = 32'd3671
; 
32'd184231: dataIn1 = 32'd9505
; 
32'd184232: dataIn1 = 32'd9506
; 
32'd184233: dataIn1 = 32'd9922
; 
32'd184234: dataIn1 = 32'd9923
; 
32'd184235: dataIn1 = 32'd9939
; 
32'd184236: dataIn1 = 32'd9940
; 
32'd184237: dataIn1 = 32'd3668
; 
32'd184238: dataIn1 = 32'd3670
; 
32'd184239: dataIn1 = 32'd3671
; 
32'd184240: dataIn1 = 32'd9504
; 
32'd184241: dataIn1 = 32'd9505
; 
32'd184242: dataIn1 = 32'd9506
; 
32'd184243: dataIn1 = 32'd9922
; 
32'd184244: dataIn1 = 32'd3673
; 
32'd184245: dataIn1 = 32'd9507
; 
32'd184246: dataIn1 = 32'd9925
; 
32'd184247: dataIn1 = 32'd9926
; 
32'd184248: dataIn1 = 32'd9930
; 
32'd184249: dataIn1 = 32'd10175
; 
32'd184250: dataIn1 = 32'd10176
; 
32'd184251: dataIn1 = 32'd9508
; 
32'd184252: dataIn1 = 32'd9518
; 
32'd184253: dataIn1 = 32'd9924
; 
32'd184254: dataIn1 = 32'd9926
; 
32'd184255: dataIn1 = 32'd9928
; 
32'd184256: dataIn1 = 32'd9929
; 
32'd184257: dataIn1 = 32'd9951
; 
32'd184258: dataIn1 = 32'd3673
; 
32'd184259: dataIn1 = 32'd9509
; 
32'd184260: dataIn1 = 32'd9924
; 
32'd184261: dataIn1 = 32'd9925
; 
32'd184262: dataIn1 = 32'd9927
; 
32'd184263: dataIn1 = 32'd9934
; 
32'd184264: dataIn1 = 32'd9935
; 
32'd184265: dataIn1 = 32'd3673
; 
32'd184266: dataIn1 = 32'd9510
; 
32'd184267: dataIn1 = 32'd9512
; 
32'd184268: dataIn1 = 32'd9932
; 
32'd184269: dataIn1 = 32'd9933
; 
32'd184270: dataIn1 = 32'd9935
; 
32'd184271: dataIn1 = 32'd9936
; 
32'd184272: dataIn1 = 32'd3671
; 
32'd184273: dataIn1 = 32'd9511
; 
32'd184274: dataIn1 = 32'd9512
; 
32'd184275: dataIn1 = 32'd9931
; 
32'd184276: dataIn1 = 32'd9933
; 
32'd184277: dataIn1 = 32'd9939
; 
32'd184278: dataIn1 = 32'd9941
; 
32'd184279: dataIn1 = 32'd2225
; 
32'd184280: dataIn1 = 32'd3671
; 
32'd184281: dataIn1 = 32'd3673
; 
32'd184282: dataIn1 = 32'd9510
; 
32'd184283: dataIn1 = 32'd9511
; 
32'd184284: dataIn1 = 32'd9512
; 
32'd184285: dataIn1 = 32'd9933
; 
32'd184286: dataIn1 = 32'd9513
; 
32'd184287: dataIn1 = 32'd9934
; 
32'd184288: dataIn1 = 32'd9936
; 
32'd184289: dataIn1 = 32'd9937
; 
32'd184290: dataIn1 = 32'd9938
; 
32'd184291: dataIn1 = 32'd10177
; 
32'd184292: dataIn1 = 32'd10178
; 
32'd184293: dataIn1 = 32'd9514
; 
32'd184294: dataIn1 = 32'd9940
; 
32'd184295: dataIn1 = 32'd9941
; 
32'd184296: dataIn1 = 32'd9942
; 
32'd184297: dataIn1 = 32'd9943
; 
32'd184298: dataIn1 = 32'd10179
; 
32'd184299: dataIn1 = 32'd10180
; 
32'd184300: dataIn1 = 32'd3679
; 
32'd184301: dataIn1 = 32'd9515
; 
32'd184302: dataIn1 = 32'd9518
; 
32'd184303: dataIn1 = 32'd9945
; 
32'd184304: dataIn1 = 32'd9946
; 
32'd184305: dataIn1 = 32'd9950
; 
32'd184306: dataIn1 = 32'd9951
; 
32'd184307: dataIn1 = 32'd9516
; 
32'd184308: dataIn1 = 32'd9944
; 
32'd184309: dataIn1 = 32'd9946
; 
32'd184310: dataIn1 = 32'd9948
; 
32'd184311: dataIn1 = 32'd9949
; 
32'd184312: dataIn1 = 32'd10181
; 
32'd184313: dataIn1 = 32'd10182
; 
32'd184314: dataIn1 = 32'd3679
; 
32'd184315: dataIn1 = 32'd9517
; 
32'd184316: dataIn1 = 32'd9519
; 
32'd184317: dataIn1 = 32'd9944
; 
32'd184318: dataIn1 = 32'd9945
; 
32'd184319: dataIn1 = 32'd9947
; 
32'd184320: dataIn1 = 32'd9952
; 
32'd184321: dataIn1 = 32'd2226
; 
32'd184322: dataIn1 = 32'd3679
; 
32'd184323: dataIn1 = 32'd3782
; 
32'd184324: dataIn1 = 32'd9508
; 
32'd184325: dataIn1 = 32'd9515
; 
32'd184326: dataIn1 = 32'd9518
; 
32'd184327: dataIn1 = 32'd9928
; 
32'd184328: dataIn1 = 32'd9951
; 
32'd184329: dataIn1 = 32'd70
; 
32'd184330: dataIn1 = 32'd3679
; 
32'd184331: dataIn1 = 32'd3784
; 
32'd184332: dataIn1 = 32'd9517
; 
32'd184333: dataIn1 = 32'd9519
; 
32'd184334: dataIn1 = 32'd9520
; 
32'd184335: dataIn1 = 32'd9952
; 
32'd184336: dataIn1 = 32'd70
; 
32'd184337: dataIn1 = 32'd9519
; 
32'd184338: dataIn1 = 32'd9520
; 
32'd184339: dataIn1 = 32'd9952
; 
32'd184340: dataIn1 = 32'd9953
; 
32'd184341: dataIn1 = 32'd9959
; 
32'd184342: dataIn1 = 32'd9960
; 
32'd184343: dataIn1 = 32'd3681
; 
32'd184344: dataIn1 = 32'd9521
; 
32'd184345: dataIn1 = 32'd9523
; 
32'd184346: dataIn1 = 32'd9525
; 
32'd184347: dataIn1 = 32'd9955
; 
32'd184348: dataIn1 = 32'd9956
; 
32'd184349: dataIn1 = 32'd9958
; 
32'd184350: dataIn1 = 32'd9522
; 
32'd184351: dataIn1 = 32'd9523
; 
32'd184352: dataIn1 = 32'd9954
; 
32'd184353: dataIn1 = 32'd9956
; 
32'd184354: dataIn1 = 32'd9959
; 
32'd184355: dataIn1 = 32'd9961
; 
32'd184356: dataIn1 = 32'd9962
; 
32'd184357: dataIn1 = 32'd3678
; 
32'd184358: dataIn1 = 32'd3681
; 
32'd184359: dataIn1 = 32'd9521
; 
32'd184360: dataIn1 = 32'd9522
; 
32'd184361: dataIn1 = 32'd9523
; 
32'd184362: dataIn1 = 32'd9956
; 
32'd184363: dataIn1 = 32'd9962
; 
32'd184364: dataIn1 = 32'd10182
; 
32'd184365: dataIn1 = 32'd10233
; 
32'd184366: dataIn1 = 32'd2228
; 
32'd184367: dataIn1 = 32'd9524
; 
32'd184368: dataIn1 = 32'd9525
; 
32'd184369: dataIn1 = 32'd9957
; 
32'd184370: dataIn1 = 32'd9958
; 
32'd184371: dataIn1 = 32'd9979
; 
32'd184372: dataIn1 = 32'd9981
; 
32'd184373: dataIn1 = 32'd2228
; 
32'd184374: dataIn1 = 32'd3681
; 
32'd184375: dataIn1 = 32'd3682
; 
32'd184376: dataIn1 = 32'd9521
; 
32'd184377: dataIn1 = 32'd9524
; 
32'd184378: dataIn1 = 32'd9525
; 
32'd184379: dataIn1 = 32'd9958
; 
32'd184380: dataIn1 = 32'd70
; 
32'd184381: dataIn1 = 32'd9526
; 
32'd184382: dataIn1 = 32'd9960
; 
32'd184383: dataIn1 = 32'd9961
; 
32'd184384: dataIn1 = 32'd9963
; 
32'd184385: dataIn1 = 32'd10183
; 
32'd184386: dataIn1 = 32'd10184
; 
32'd184387: dataIn1 = 32'd3689
; 
32'd184388: dataIn1 = 32'd9527
; 
32'd184389: dataIn1 = 32'd9965
; 
32'd184390: dataIn1 = 32'd9966
; 
32'd184391: dataIn1 = 32'd9970
; 
32'd184392: dataIn1 = 32'd10185
; 
32'd184393: dataIn1 = 32'd10186
; 
32'd184394: dataIn1 = 32'd3689
; 
32'd184395: dataIn1 = 32'd9528
; 
32'd184396: dataIn1 = 32'd9964
; 
32'd184397: dataIn1 = 32'd9966
; 
32'd184398: dataIn1 = 32'd9968
; 
32'd184399: dataIn1 = 32'd9971
; 
32'd184400: dataIn1 = 32'd9973
; 
32'd184401: dataIn1 = 32'd9529
; 
32'd184402: dataIn1 = 32'd9533
; 
32'd184403: dataIn1 = 32'd9964
; 
32'd184404: dataIn1 = 32'd9965
; 
32'd184405: dataIn1 = 32'd9967
; 
32'd184406: dataIn1 = 32'd9969
; 
32'd184407: dataIn1 = 32'd9977
; 
32'd184408: dataIn1 = 32'd3689
; 
32'd184409: dataIn1 = 32'd9530
; 
32'd184410: dataIn1 = 32'd9535
; 
32'd184411: dataIn1 = 32'd9972
; 
32'd184412: dataIn1 = 32'd9973
; 
32'd184413: dataIn1 = 32'd9976
; 
32'd184414: dataIn1 = 32'd9985
; 
32'd184415: dataIn1 = 32'd9531
; 
32'd184416: dataIn1 = 32'd9971
; 
32'd184417: dataIn1 = 32'd9972
; 
32'd184418: dataIn1 = 32'd9974
; 
32'd184419: dataIn1 = 32'd9975
; 
32'd184420: dataIn1 = 32'd10187
; 
32'd184421: dataIn1 = 32'd10188
; 
32'd184422: dataIn1 = 32'd2228
; 
32'd184423: dataIn1 = 32'd9532
; 
32'd184424: dataIn1 = 32'd9533
; 
32'd184425: dataIn1 = 32'd9977
; 
32'd184426: dataIn1 = 32'd9978
; 
32'd184427: dataIn1 = 32'd9980
; 
32'd184428: dataIn1 = 32'd9981
; 
32'd184429: dataIn1 = 32'd2228
; 
32'd184430: dataIn1 = 32'd3686
; 
32'd184431: dataIn1 = 32'd3687
; 
32'd184432: dataIn1 = 32'd9529
; 
32'd184433: dataIn1 = 32'd9532
; 
32'd184434: dataIn1 = 32'd9533
; 
32'd184435: dataIn1 = 32'd9967
; 
32'd184436: dataIn1 = 32'd9977
; 
32'd184437: dataIn1 = 32'd9534
; 
32'd184438: dataIn1 = 32'd9979
; 
32'd184439: dataIn1 = 32'd9980
; 
32'd184440: dataIn1 = 32'd9982
; 
32'd184441: dataIn1 = 32'd9983
; 
32'd184442: dataIn1 = 32'd10184
; 
32'd184443: dataIn1 = 32'd10189
; 
32'd184444: dataIn1 = 32'd3689
; 
32'd184445: dataIn1 = 32'd3692
; 
32'd184446: dataIn1 = 32'd3693
; 
32'd184447: dataIn1 = 32'd9530
; 
32'd184448: dataIn1 = 32'd9535
; 
32'd184449: dataIn1 = 32'd9536
; 
32'd184450: dataIn1 = 32'd9985
; 
32'd184451: dataIn1 = 32'd3692
; 
32'd184452: dataIn1 = 32'd9535
; 
32'd184453: dataIn1 = 32'd9536
; 
32'd184454: dataIn1 = 32'd9544
; 
32'd184455: dataIn1 = 32'd9984
; 
32'd184456: dataIn1 = 32'd9985
; 
32'd184457: dataIn1 = 32'd10001
; 
32'd184458: dataIn1 = 32'd9537
; 
32'd184459: dataIn1 = 32'd9538
; 
32'd184460: dataIn1 = 32'd9987
; 
32'd184461: dataIn1 = 32'd9988
; 
32'd184462: dataIn1 = 32'd9990
; 
32'd184463: dataIn1 = 32'd9991
; 
32'd184464: dataIn1 = 32'd9994
; 
32'd184465: dataIn1 = 32'd2201
; 
32'd184466: dataIn1 = 32'd3694
; 
32'd184467: dataIn1 = 32'd3696
; 
32'd184468: dataIn1 = 32'd9537
; 
32'd184469: dataIn1 = 32'd9538
; 
32'd184470: dataIn1 = 32'd9539
; 
32'd184471: dataIn1 = 32'd9987
; 
32'd184472: dataIn1 = 32'd9994
; 
32'd184473: dataIn1 = 32'd3694
; 
32'd184474: dataIn1 = 32'd9538
; 
32'd184475: dataIn1 = 32'd9539
; 
32'd184476: dataIn1 = 32'd9986
; 
32'd184477: dataIn1 = 32'd9987
; 
32'd184478: dataIn1 = 32'd9995
; 
32'd184479: dataIn1 = 32'd9996
; 
32'd184480: dataIn1 = 32'd2231
; 
32'd184481: dataIn1 = 32'd9540
; 
32'd184482: dataIn1 = 32'd9989
; 
32'd184483: dataIn1 = 32'd9991
; 
32'd184484: dataIn1 = 32'd9993
; 
32'd184485: dataIn1 = 32'd10005
; 
32'd184486: dataIn1 = 32'd10007
; 
32'd184487: dataIn1 = 32'd2231
; 
32'd184488: dataIn1 = 32'd9541
; 
32'd184489: dataIn1 = 32'd9989
; 
32'd184490: dataIn1 = 32'd9990
; 
32'd184491: dataIn1 = 32'd9992
; 
32'd184492: dataIn1 = 32'd10190
; 
32'd184493: dataIn1 = 32'd10191
; 
32'd184494: dataIn1 = 32'd9542
; 
32'd184495: dataIn1 = 32'd9544
; 
32'd184496: dataIn1 = 32'd9996
; 
32'd184497: dataIn1 = 32'd9997
; 
32'd184498: dataIn1 = 32'd9998
; 
32'd184499: dataIn1 = 32'd10000
; 
32'd184500: dataIn1 = 32'd10001
; 
32'd184501: dataIn1 = 32'd3694
; 
32'd184502: dataIn1 = 32'd9543
; 
32'd184503: dataIn1 = 32'd9995
; 
32'd184504: dataIn1 = 32'd9997
; 
32'd184505: dataIn1 = 32'd9999
; 
32'd184506: dataIn1 = 32'd10187
; 
32'd184507: dataIn1 = 32'd10192
; 
32'd184508: dataIn1 = 32'd3692
; 
32'd184509: dataIn1 = 32'd3695
; 
32'd184510: dataIn1 = 32'd9536
; 
32'd184511: dataIn1 = 32'd9542
; 
32'd184512: dataIn1 = 32'd9544
; 
32'd184513: dataIn1 = 32'd9998
; 
32'd184514: dataIn1 = 32'd10001
; 
32'd184515: dataIn1 = 32'd10190
; 
32'd184516: dataIn1 = 32'd10235
; 
32'd184517: dataIn1 = 32'd9545
; 
32'd184518: dataIn1 = 32'd9546
; 
32'd184519: dataIn1 = 32'd10003
; 
32'd184520: dataIn1 = 32'd10004
; 
32'd184521: dataIn1 = 32'd10006
; 
32'd184522: dataIn1 = 32'd10007
; 
32'd184523: dataIn1 = 32'd10009
; 
32'd184524: dataIn1 = 32'd2201
; 
32'd184525: dataIn1 = 32'd3617
; 
32'd184526: dataIn1 = 32'd3696
; 
32'd184527: dataIn1 = 32'd9545
; 
32'd184528: dataIn1 = 32'd9546
; 
32'd184529: dataIn1 = 32'd9547
; 
32'd184530: dataIn1 = 32'd10003
; 
32'd184531: dataIn1 = 32'd10009
; 
32'd184532: dataIn1 = 32'd3617
; 
32'd184533: dataIn1 = 32'd9546
; 
32'd184534: dataIn1 = 32'd9547
; 
32'd184535: dataIn1 = 32'd9550
; 
32'd184536: dataIn1 = 32'd10002
; 
32'd184537: dataIn1 = 32'd10003
; 
32'd184538: dataIn1 = 32'd10010
; 
32'd184539: dataIn1 = 32'd2231
; 
32'd184540: dataIn1 = 32'd9548
; 
32'd184541: dataIn1 = 32'd10005
; 
32'd184542: dataIn1 = 32'd10006
; 
32'd184543: dataIn1 = 32'd10008
; 
32'd184544: dataIn1 = 32'd10193
; 
32'd184545: dataIn1 = 32'd10194
; 
32'd184546: dataIn1 = 32'd61
; 
32'd184547: dataIn1 = 32'd9549
; 
32'd184548: dataIn1 = 32'd9550
; 
32'd184549: dataIn1 = 32'd10010
; 
32'd184550: dataIn1 = 32'd10011
; 
32'd184551: dataIn1 = 32'd10012
; 
32'd184552: dataIn1 = 32'd10013
; 
32'd184553: dataIn1 = 32'd61
; 
32'd184554: dataIn1 = 32'd3616
; 
32'd184555: dataIn1 = 32'd3617
; 
32'd184556: dataIn1 = 32'd9547
; 
32'd184557: dataIn1 = 32'd9549
; 
32'd184558: dataIn1 = 32'd9550
; 
32'd184559: dataIn1 = 32'd10010
; 
32'd184560: dataIn1 = 32'd9551
; 
32'd184561: dataIn1 = 32'd10013
; 
32'd184562: dataIn1 = 32'd10014
; 
32'd184563: dataIn1 = 32'd10015
; 
32'd184564: dataIn1 = 32'd10017
; 
32'd184565: dataIn1 = 32'd10194
; 
32'd184566: dataIn1 = 32'd10195
; 
32'd184567: dataIn1 = 32'd61
; 
32'd184568: dataIn1 = 32'd9552
; 
32'd184569: dataIn1 = 32'd10012
; 
32'd184570: dataIn1 = 32'd10014
; 
32'd184571: dataIn1 = 32'd10016
; 
32'd184572: dataIn1 = 32'd10021
; 
32'd184573: dataIn1 = 32'd10022
; 
32'd184574: dataIn1 = 32'd9553
; 
32'd184575: dataIn1 = 32'd9555
; 
32'd184576: dataIn1 = 32'd10019
; 
32'd184577: dataIn1 = 32'd10020
; 
32'd184578: dataIn1 = 32'd10022
; 
32'd184579: dataIn1 = 32'd10023
; 
32'd184580: dataIn1 = 32'd10024
; 
32'd184581: dataIn1 = 32'd3706
; 
32'd184582: dataIn1 = 32'd9554
; 
32'd184583: dataIn1 = 32'd9555
; 
32'd184584: dataIn1 = 32'd9557
; 
32'd184585: dataIn1 = 32'd10018
; 
32'd184586: dataIn1 = 32'd10020
; 
32'd184587: dataIn1 = 32'd10026
; 
32'd184588: dataIn1 = 32'd2233
; 
32'd184589: dataIn1 = 32'd3702
; 
32'd184590: dataIn1 = 32'd3706
; 
32'd184591: dataIn1 = 32'd9553
; 
32'd184592: dataIn1 = 32'd9554
; 
32'd184593: dataIn1 = 32'd9555
; 
32'd184594: dataIn1 = 32'd10020
; 
32'd184595: dataIn1 = 32'd10024
; 
32'd184596: dataIn1 = 32'd61
; 
32'd184597: dataIn1 = 32'd9556
; 
32'd184598: dataIn1 = 32'd10021
; 
32'd184599: dataIn1 = 32'd10023
; 
32'd184600: dataIn1 = 32'd10025
; 
32'd184601: dataIn1 = 32'd10164
; 
32'd184602: dataIn1 = 32'd10196
; 
32'd184603: dataIn1 = 32'd2204
; 
32'd184604: dataIn1 = 32'd3706
; 
32'd184605: dataIn1 = 32'd3708
; 
32'd184606: dataIn1 = 32'd9486
; 
32'd184607: dataIn1 = 32'd9554
; 
32'd184608: dataIn1 = 32'd9557
; 
32'd184609: dataIn1 = 32'd10026
; 
32'd184610: dataIn1 = 32'd9558
; 
32'd184611: dataIn1 = 32'd10028
; 
32'd184612: dataIn1 = 32'd10029
; 
32'd184613: dataIn1 = 32'd10031
; 
32'd184614: dataIn1 = 32'd10033
; 
32'd184615: dataIn1 = 32'd10198
; 
32'd184616: dataIn1 = 32'd66
; 
32'd184617: dataIn1 = 32'd9559
; 
32'd184618: dataIn1 = 32'd9567
; 
32'd184619: dataIn1 = 32'd10027
; 
32'd184620: dataIn1 = 32'd10029
; 
32'd184621: dataIn1 = 32'd10032
; 
32'd184622: dataIn1 = 32'd10048
; 
32'd184623: dataIn1 = 32'd66
; 
32'd184624: dataIn1 = 32'd9560
; 
32'd184625: dataIn1 = 32'd10027
; 
32'd184626: dataIn1 = 32'd10028
; 
32'd184627: dataIn1 = 32'd10030
; 
32'd184628: dataIn1 = 32'd3743
; 
32'd184629: dataIn1 = 32'd9561
; 
32'd184630: dataIn1 = 32'd10035
; 
32'd184631: dataIn1 = 32'd10036
; 
32'd184632: dataIn1 = 32'd10040
; 
32'd184633: dataIn1 = 32'd10054
; 
32'd184634: dataIn1 = 32'd10055
; 
32'd184635: dataIn1 = 32'd3743
; 
32'd184636: dataIn1 = 32'd9562
; 
32'd184637: dataIn1 = 32'd10034
; 
32'd184638: dataIn1 = 32'd10036
; 
32'd184639: dataIn1 = 32'd10038
; 
32'd184640: dataIn1 = 32'd10199
; 
32'd184641: dataIn1 = 32'd10200
; 
32'd184642: dataIn1 = 32'd9563
; 
32'd184643: dataIn1 = 32'd9568
; 
32'd184644: dataIn1 = 32'd10034
; 
32'd184645: dataIn1 = 32'd10035
; 
32'd184646: dataIn1 = 32'd10037
; 
32'd184647: dataIn1 = 32'd10039
; 
32'd184648: dataIn1 = 32'd10049
; 
32'd184649: dataIn1 = 32'd3744
; 
32'd184650: dataIn1 = 32'd9564
; 
32'd184651: dataIn1 = 32'd9567
; 
32'd184652: dataIn1 = 32'd10042
; 
32'd184653: dataIn1 = 32'd10043
; 
32'd184654: dataIn1 = 32'd10047
; 
32'd184655: dataIn1 = 32'd10048
; 
32'd184656: dataIn1 = 32'd3744
; 
32'd184657: dataIn1 = 32'd9565
; 
32'd184658: dataIn1 = 32'd9568
; 
32'd184659: dataIn1 = 32'd10041
; 
32'd184660: dataIn1 = 32'd10043
; 
32'd184661: dataIn1 = 32'd10045
; 
32'd184662: dataIn1 = 32'd10049
; 
32'd184663: dataIn1 = 32'd9566
; 
32'd184664: dataIn1 = 32'd10041
; 
32'd184665: dataIn1 = 32'd10042
; 
32'd184666: dataIn1 = 32'd10044
; 
32'd184667: dataIn1 = 32'd10046
; 
32'd184668: dataIn1 = 32'd10201
; 
32'd184669: dataIn1 = 32'd10202
; 
32'd184670: dataIn1 = 32'd66
; 
32'd184671: dataIn1 = 32'd3658
; 
32'd184672: dataIn1 = 32'd3744
; 
32'd184673: dataIn1 = 32'd9559
; 
32'd184674: dataIn1 = 32'd9564
; 
32'd184675: dataIn1 = 32'd9567
; 
32'd184676: dataIn1 = 32'd10048
; 
32'd184677: dataIn1 = 32'd2217
; 
32'd184678: dataIn1 = 32'd3744
; 
32'd184679: dataIn1 = 32'd5310
; 
32'd184680: dataIn1 = 32'd9563
; 
32'd184681: dataIn1 = 32'd9565
; 
32'd184682: dataIn1 = 32'd9568
; 
32'd184683: dataIn1 = 32'd10039
; 
32'd184684: dataIn1 = 32'd10049
; 
32'd184685: dataIn1 = 32'd2244
; 
32'd184686: dataIn1 = 32'd3743
; 
32'd184687: dataIn1 = 32'd3747
; 
32'd184688: dataIn1 = 32'd9569
; 
32'd184689: dataIn1 = 32'd9570
; 
32'd184690: dataIn1 = 32'd9571
; 
32'd184691: dataIn1 = 32'd10050
; 
32'd184692: dataIn1 = 32'd3743
; 
32'd184693: dataIn1 = 32'd9569
; 
32'd184694: dataIn1 = 32'd9570
; 
32'd184695: dataIn1 = 32'd10050
; 
32'd184696: dataIn1 = 32'd10052
; 
32'd184697: dataIn1 = 32'd10053
; 
32'd184698: dataIn1 = 32'd10055
; 
32'd184699: dataIn1 = 32'd3747
; 
32'd184700: dataIn1 = 32'd9569
; 
32'd184701: dataIn1 = 32'd9571
; 
32'd184702: dataIn1 = 32'd10050
; 
32'd184703: dataIn1 = 32'd10051
; 
32'd184704: dataIn1 = 32'd10058
; 
32'd184705: dataIn1 = 32'd10059
; 
32'd184706: dataIn1 = 32'd9572
; 
32'd184707: dataIn1 = 32'd10053
; 
32'd184708: dataIn1 = 32'd10054
; 
32'd184709: dataIn1 = 32'd10056
; 
32'd184710: dataIn1 = 32'd10057
; 
32'd184711: dataIn1 = 32'd10203
; 
32'd184712: dataIn1 = 32'd10204
; 
32'd184713: dataIn1 = 32'd3747
; 
32'd184714: dataIn1 = 32'd9573
; 
32'd184715: dataIn1 = 32'd9575
; 
32'd184716: dataIn1 = 32'd10059
; 
32'd184717: dataIn1 = 32'd10060
; 
32'd184718: dataIn1 = 32'd10063
; 
32'd184719: dataIn1 = 32'd10064
; 
32'd184720: dataIn1 = 32'd9574
; 
32'd184721: dataIn1 = 32'd10058
; 
32'd184722: dataIn1 = 32'd10060
; 
32'd184723: dataIn1 = 32'd10061
; 
32'd184724: dataIn1 = 32'd10062
; 
32'd184725: dataIn1 = 32'd10205
; 
32'd184726: dataIn1 = 32'd10206
; 
32'd184727: dataIn1 = 32'd3747
; 
32'd184728: dataIn1 = 32'd3748
; 
32'd184729: dataIn1 = 32'd3751
; 
32'd184730: dataIn1 = 32'd9573
; 
32'd184731: dataIn1 = 32'd9575
; 
32'd184732: dataIn1 = 32'd9576
; 
32'd184733: dataIn1 = 32'd10064
; 
32'd184734: dataIn1 = 32'd3751
; 
32'd184735: dataIn1 = 32'd9575
; 
32'd184736: dataIn1 = 32'd9576
; 
32'd184737: dataIn1 = 32'd10064
; 
32'd184738: dataIn1 = 32'd10065
; 
32'd184739: dataIn1 = 32'd10072
; 
32'd184740: dataIn1 = 32'd10073
; 
32'd184741: dataIn1 = 32'd3757
; 
32'd184742: dataIn1 = 32'd9577
; 
32'd184743: dataIn1 = 32'd9578
; 
32'd184744: dataIn1 = 32'd10067
; 
32'd184745: dataIn1 = 32'd10068
; 
32'd184746: dataIn1 = 32'd10086
; 
32'd184747: dataIn1 = 32'd10087
; 
32'd184748: dataIn1 = 32'd3755
; 
32'd184749: dataIn1 = 32'd3756
; 
32'd184750: dataIn1 = 32'd3757
; 
32'd184751: dataIn1 = 32'd9577
; 
32'd184752: dataIn1 = 32'd9578
; 
32'd184753: dataIn1 = 32'd9579
; 
32'd184754: dataIn1 = 32'd10067
; 
32'd184755: dataIn1 = 32'd3755
; 
32'd184756: dataIn1 = 32'd9578
; 
32'd184757: dataIn1 = 32'd9579
; 
32'd184758: dataIn1 = 32'd10066
; 
32'd184759: dataIn1 = 32'd10067
; 
32'd184760: dataIn1 = 32'd10077
; 
32'd184761: dataIn1 = 32'd10078
; 
32'd184762: dataIn1 = 32'd3751
; 
32'd184763: dataIn1 = 32'd9580
; 
32'd184764: dataIn1 = 32'd9582
; 
32'd184765: dataIn1 = 32'd10070
; 
32'd184766: dataIn1 = 32'd10071
; 
32'd184767: dataIn1 = 32'd10073
; 
32'd184768: dataIn1 = 32'd10074
; 
32'd184769: dataIn1 = 32'd3755
; 
32'd184770: dataIn1 = 32'd9581
; 
32'd184771: dataIn1 = 32'd9582
; 
32'd184772: dataIn1 = 32'd10069
; 
32'd184773: dataIn1 = 32'd10071
; 
32'd184774: dataIn1 = 32'd10077
; 
32'd184775: dataIn1 = 32'd10079
; 
32'd184776: dataIn1 = 32'd2246
; 
32'd184777: dataIn1 = 32'd3751
; 
32'd184778: dataIn1 = 32'd3755
; 
32'd184779: dataIn1 = 32'd9580
; 
32'd184780: dataIn1 = 32'd9581
; 
32'd184781: dataIn1 = 32'd9582
; 
32'd184782: dataIn1 = 32'd10071
; 
32'd184783: dataIn1 = 32'd9583
; 
32'd184784: dataIn1 = 32'd10072
; 
32'd184785: dataIn1 = 32'd10074
; 
32'd184786: dataIn1 = 32'd10075
; 
32'd184787: dataIn1 = 32'd10076
; 
32'd184788: dataIn1 = 32'd10207
; 
32'd184789: dataIn1 = 32'd10208
; 
32'd184790: dataIn1 = 32'd9584
; 
32'd184791: dataIn1 = 32'd10078
; 
32'd184792: dataIn1 = 32'd10079
; 
32'd184793: dataIn1 = 32'd10080
; 
32'd184794: dataIn1 = 32'd10081
; 
32'd184795: dataIn1 = 32'd10209
; 
32'd184796: dataIn1 = 32'd10210
; 
32'd184797: dataIn1 = 32'd2247
; 
32'd184798: dataIn1 = 32'd3757
; 
32'd184799: dataIn1 = 32'd3760
; 
32'd184800: dataIn1 = 32'd9585
; 
32'd184801: dataIn1 = 32'd9586
; 
32'd184802: dataIn1 = 32'd9587
; 
32'd184803: dataIn1 = 32'd10082
; 
32'd184804: dataIn1 = 32'd3757
; 
32'd184805: dataIn1 = 32'd9585
; 
32'd184806: dataIn1 = 32'd9586
; 
32'd184807: dataIn1 = 32'd10082
; 
32'd184808: dataIn1 = 32'd10084
; 
32'd184809: dataIn1 = 32'd10085
; 
32'd184810: dataIn1 = 32'd10087
; 
32'd184811: dataIn1 = 32'd3760
; 
32'd184812: dataIn1 = 32'd9585
; 
32'd184813: dataIn1 = 32'd9587
; 
32'd184814: dataIn1 = 32'd10082
; 
32'd184815: dataIn1 = 32'd10083
; 
32'd184816: dataIn1 = 32'd10090
; 
32'd184817: dataIn1 = 32'd10091
; 
32'd184818: dataIn1 = 32'd9588
; 
32'd184819: dataIn1 = 32'd10085
; 
32'd184820: dataIn1 = 32'd10086
; 
32'd184821: dataIn1 = 32'd10088
; 
32'd184822: dataIn1 = 32'd10089
; 
32'd184823: dataIn1 = 32'd10211
; 
32'd184824: dataIn1 = 32'd10212
; 
32'd184825: dataIn1 = 32'd3760
; 
32'd184826: dataIn1 = 32'd9589
; 
32'd184827: dataIn1 = 32'd9591
; 
32'd184828: dataIn1 = 32'd10091
; 
32'd184829: dataIn1 = 32'd10092
; 
32'd184830: dataIn1 = 32'd10095
; 
32'd184831: dataIn1 = 32'd10096
; 
32'd184832: dataIn1 = 32'd9590
; 
32'd184833: dataIn1 = 32'd10090
; 
32'd184834: dataIn1 = 32'd10092
; 
32'd184835: dataIn1 = 32'd10093
; 
32'd184836: dataIn1 = 32'd10094
; 
32'd184837: dataIn1 = 32'd10213
; 
32'd184838: dataIn1 = 32'd10214
; 
32'd184839: dataIn1 = 32'd3760
; 
32'd184840: dataIn1 = 32'd3761
; 
32'd184841: dataIn1 = 32'd3764
; 
32'd184842: dataIn1 = 32'd9589
; 
32'd184843: dataIn1 = 32'd9591
; 
32'd184844: dataIn1 = 32'd9592
; 
32'd184845: dataIn1 = 32'd10096
; 
32'd184846: dataIn1 = 32'd3764
; 
32'd184847: dataIn1 = 32'd9591
; 
32'd184848: dataIn1 = 32'd9592
; 
32'd184849: dataIn1 = 32'd10096
; 
32'd184850: dataIn1 = 32'd10097
; 
32'd184851: dataIn1 = 32'd10104
; 
32'd184852: dataIn1 = 32'd10105
; 
32'd184853: dataIn1 = 32'd3770
; 
32'd184854: dataIn1 = 32'd9593
; 
32'd184855: dataIn1 = 32'd9594
; 
32'd184856: dataIn1 = 32'd10099
; 
32'd184857: dataIn1 = 32'd10100
; 
32'd184858: dataIn1 = 32'd10115
; 
32'd184859: dataIn1 = 32'd10116
; 
32'd184860: dataIn1 = 32'd3768
; 
32'd184861: dataIn1 = 32'd3769
; 
32'd184862: dataIn1 = 32'd3770
; 
32'd184863: dataIn1 = 32'd9593
; 
32'd184864: dataIn1 = 32'd9594
; 
32'd184865: dataIn1 = 32'd9595
; 
32'd184866: dataIn1 = 32'd10099
; 
32'd184867: dataIn1 = 32'd3768
; 
32'd184868: dataIn1 = 32'd9594
; 
32'd184869: dataIn1 = 32'd9595
; 
32'd184870: dataIn1 = 32'd10098
; 
32'd184871: dataIn1 = 32'd10099
; 
32'd184872: dataIn1 = 32'd10109
; 
32'd184873: dataIn1 = 32'd10110
; 
32'd184874: dataIn1 = 32'd3764
; 
32'd184875: dataIn1 = 32'd9596
; 
32'd184876: dataIn1 = 32'd9598
; 
32'd184877: dataIn1 = 32'd10102
; 
32'd184878: dataIn1 = 32'd10103
; 
32'd184879: dataIn1 = 32'd10105
; 
32'd184880: dataIn1 = 32'd10106
; 
32'd184881: dataIn1 = 32'd3768
; 
32'd184882: dataIn1 = 32'd9597
; 
32'd184883: dataIn1 = 32'd9598
; 
32'd184884: dataIn1 = 32'd10101
; 
32'd184885: dataIn1 = 32'd10103
; 
32'd184886: dataIn1 = 32'd10109
; 
32'd184887: dataIn1 = 32'd10111
; 
32'd184888: dataIn1 = 32'd2249
; 
32'd184889: dataIn1 = 32'd3764
; 
32'd184890: dataIn1 = 32'd3768
; 
32'd184891: dataIn1 = 32'd9596
; 
32'd184892: dataIn1 = 32'd9597
; 
32'd184893: dataIn1 = 32'd9598
; 
32'd184894: dataIn1 = 32'd10103
; 
32'd184895: dataIn1 = 32'd9599
; 
32'd184896: dataIn1 = 32'd10104
; 
32'd184897: dataIn1 = 32'd10106
; 
32'd184898: dataIn1 = 32'd10107
; 
32'd184899: dataIn1 = 32'd10108
; 
32'd184900: dataIn1 = 32'd10215
; 
32'd184901: dataIn1 = 32'd10216
; 
32'd184902: dataIn1 = 32'd9600
; 
32'd184903: dataIn1 = 32'd10110
; 
32'd184904: dataIn1 = 32'd10111
; 
32'd184905: dataIn1 = 32'd10112
; 
32'd184906: dataIn1 = 32'd10113
; 
32'd184907: dataIn1 = 32'd10217
; 
32'd184908: dataIn1 = 32'd10218
; 
32'd184909: dataIn1 = 32'd3770
; 
32'd184910: dataIn1 = 32'd9601
; 
32'd184911: dataIn1 = 32'd10114
; 
32'd184912: dataIn1 = 32'd10116
; 
32'd184913: dataIn1 = 32'd10117
; 
32'd184914: dataIn1 = 32'd10174
; 
32'd184915: dataIn1 = 32'd10219
; 
32'd184916: dataIn1 = 32'd4684
; 
32'd184917: dataIn1 = 32'd4687
; 
32'd184918: dataIn1 = 32'd4688
; 
32'd184919: dataIn1 = 32'd9602
; 
32'd184920: dataIn1 = 32'd9603
; 
32'd184921: dataIn1 = 32'd9604
; 
32'd184922: dataIn1 = 32'd133
; 
32'd184923: dataIn1 = 32'd4688
; 
32'd184924: dataIn1 = 32'd7576
; 
32'd184925: dataIn1 = 32'd9602
; 
32'd184926: dataIn1 = 32'd9603
; 
32'd184927: dataIn1 = 32'd9604
; 
32'd184928: dataIn1 = 32'd9629
; 
32'd184929: dataIn1 = 32'd133
; 
32'd184930: dataIn1 = 32'd4687
; 
32'd184931: dataIn1 = 32'd7489
; 
32'd184932: dataIn1 = 32'd9602
; 
32'd184933: dataIn1 = 32'd9603
; 
32'd184934: dataIn1 = 32'd9604
; 
32'd184935: dataIn1 = 32'd9617
; 
32'd184936: dataIn1 = 32'd7
; 
32'd184937: dataIn1 = 32'd4699
; 
32'd184938: dataIn1 = 32'd7712
; 
32'd184939: dataIn1 = 32'd9605
; 
32'd184940: dataIn1 = 32'd9606
; 
32'd184941: dataIn1 = 32'd9607
; 
32'd184942: dataIn1 = 32'd9660
; 
32'd184943: dataIn1 = 32'd4694
; 
32'd184944: dataIn1 = 32'd4698
; 
32'd184945: dataIn1 = 32'd4699
; 
32'd184946: dataIn1 = 32'd9605
; 
32'd184947: dataIn1 = 32'd9606
; 
32'd184948: dataIn1 = 32'd9607
; 
32'd184949: dataIn1 = 32'd7
; 
32'd184950: dataIn1 = 32'd4698
; 
32'd184951: dataIn1 = 32'd7606
; 
32'd184952: dataIn1 = 32'd9605
; 
32'd184953: dataIn1 = 32'd9606
; 
32'd184954: dataIn1 = 32'd9607
; 
32'd184955: dataIn1 = 32'd9643
; 
32'd184956: dataIn1 = 32'd4702
; 
32'd184957: dataIn1 = 32'd4705
; 
32'd184958: dataIn1 = 32'd4706
; 
32'd184959: dataIn1 = 32'd9608
; 
32'd184960: dataIn1 = 32'd9609
; 
32'd184961: dataIn1 = 32'd9610
; 
32'd184962: dataIn1 = 32'd136
; 
32'd184963: dataIn1 = 32'd4706
; 
32'd184964: dataIn1 = 32'd7829
; 
32'd184965: dataIn1 = 32'd9608
; 
32'd184966: dataIn1 = 32'd9609
; 
32'd184967: dataIn1 = 32'd9610
; 
32'd184968: dataIn1 = 32'd9665
; 
32'd184969: dataIn1 = 32'd136
; 
32'd184970: dataIn1 = 32'd4705
; 
32'd184971: dataIn1 = 32'd7742
; 
32'd184972: dataIn1 = 32'd9608
; 
32'd184973: dataIn1 = 32'd9609
; 
32'd184974: dataIn1 = 32'd9610
; 
32'd184975: dataIn1 = 32'd9650
; 
32'd184976: dataIn1 = 32'd1107
; 
32'd184977: dataIn1 = 32'd4892
; 
32'd184978: dataIn1 = 32'd7494
; 
32'd184979: dataIn1 = 32'd9611
; 
32'd184980: dataIn1 = 32'd9612
; 
32'd184981: dataIn1 = 32'd9613
; 
32'd184982: dataIn1 = 32'd9622
; 
32'd184983: dataIn1 = 32'd1107
; 
32'd184984: dataIn1 = 32'd4891
; 
32'd184985: dataIn1 = 32'd7472
; 
32'd184986: dataIn1 = 32'd9611
; 
32'd184987: dataIn1 = 32'd9612
; 
32'd184988: dataIn1 = 32'd9613
; 
32'd184989: dataIn1 = 32'd9763
; 
32'd184990: dataIn1 = 32'd4886
; 
32'd184991: dataIn1 = 32'd4891
; 
32'd184992: dataIn1 = 32'd4892
; 
32'd184993: dataIn1 = 32'd9611
; 
32'd184994: dataIn1 = 32'd9612
; 
32'd184995: dataIn1 = 32'd9613
; 
32'd184996: dataIn1 = 32'd2635
; 
32'd184997: dataIn1 = 32'd4895
; 
32'd184998: dataIn1 = 32'd7493
; 
32'd184999: dataIn1 = 32'd9614
; 
32'd185000: dataIn1 = 32'd9615
; 
32'd185001: dataIn1 = 32'd9616
; 
32'd185002: dataIn1 = 32'd9621
; 
32'd185003: dataIn1 = 32'd4893
; 
32'd185004: dataIn1 = 32'd4894
; 
32'd185005: dataIn1 = 32'd4895
; 
32'd185006: dataIn1 = 32'd9614
; 
32'd185007: dataIn1 = 32'd9615
; 
32'd185008: dataIn1 = 32'd9616
; 
32'd185009: dataIn1 = 32'd2635
; 
32'd185010: dataIn1 = 32'd4893
; 
32'd185011: dataIn1 = 32'd7488
; 
32'd185012: dataIn1 = 32'd9614
; 
32'd185013: dataIn1 = 32'd9615
; 
32'd185014: dataIn1 = 32'd9616
; 
32'd185015: dataIn1 = 32'd9618
; 
32'd185016: dataIn1 = 32'd4687
; 
32'd185017: dataIn1 = 32'd4896
; 
32'd185018: dataIn1 = 32'd7489
; 
32'd185019: dataIn1 = 32'd9604
; 
32'd185020: dataIn1 = 32'd9617
; 
32'd185021: dataIn1 = 32'd9618
; 
32'd185022: dataIn1 = 32'd9619
; 
32'd185023: dataIn1 = 32'd4893
; 
32'd185024: dataIn1 = 32'd4896
; 
32'd185025: dataIn1 = 32'd7488
; 
32'd185026: dataIn1 = 32'd9616
; 
32'd185027: dataIn1 = 32'd9617
; 
32'd185028: dataIn1 = 32'd9618
; 
32'd185029: dataIn1 = 32'd9619
; 
32'd185030: dataIn1 = 32'd2573
; 
32'd185031: dataIn1 = 32'd4687
; 
32'd185032: dataIn1 = 32'd4893
; 
32'd185033: dataIn1 = 32'd9617
; 
32'd185034: dataIn1 = 32'd9618
; 
32'd185035: dataIn1 = 32'd9619
; 
32'd185036: dataIn1 = 32'd2632
; 
32'd185037: dataIn1 = 32'd4892
; 
32'd185038: dataIn1 = 32'd4895
; 
32'd185039: dataIn1 = 32'd9620
; 
32'd185040: dataIn1 = 32'd9621
; 
32'd185041: dataIn1 = 32'd9622
; 
32'd185042: dataIn1 = 32'd4895
; 
32'd185043: dataIn1 = 32'd4897
; 
32'd185044: dataIn1 = 32'd7493
; 
32'd185045: dataIn1 = 32'd9614
; 
32'd185046: dataIn1 = 32'd9620
; 
32'd185047: dataIn1 = 32'd9621
; 
32'd185048: dataIn1 = 32'd9622
; 
32'd185049: dataIn1 = 32'd4892
; 
32'd185050: dataIn1 = 32'd4897
; 
32'd185051: dataIn1 = 32'd7494
; 
32'd185052: dataIn1 = 32'd9611
; 
32'd185053: dataIn1 = 32'd9620
; 
32'd185054: dataIn1 = 32'd9621
; 
32'd185055: dataIn1 = 32'd9622
; 
32'd185056: dataIn1 = 32'd1108
; 
32'd185057: dataIn1 = 32'd4909
; 
32'd185058: dataIn1 = 32'd7571
; 
32'd185059: dataIn1 = 32'd9623
; 
32'd185060: dataIn1 = 32'd9624
; 
32'd185061: dataIn1 = 32'd9625
; 
32'd185062: dataIn1 = 32'd9633
; 
32'd185063: dataIn1 = 32'd4904
; 
32'd185064: dataIn1 = 32'd4908
; 
32'd185065: dataIn1 = 32'd4909
; 
32'd185066: dataIn1 = 32'd9623
; 
32'd185067: dataIn1 = 32'd9624
; 
32'd185068: dataIn1 = 32'd9625
; 
32'd185069: dataIn1 = 32'd1108
; 
32'd185070: dataIn1 = 32'd4908
; 
32'd185071: dataIn1 = 32'd7593
; 
32'd185072: dataIn1 = 32'd9623
; 
32'd185073: dataIn1 = 32'd9624
; 
32'd185074: dataIn1 = 32'd9625
; 
32'd185075: dataIn1 = 32'd9639
; 
32'd185076: dataIn1 = 32'd2640
; 
32'd185077: dataIn1 = 32'd4913
; 
32'd185078: dataIn1 = 32'd7572
; 
32'd185079: dataIn1 = 32'd9626
; 
32'd185080: dataIn1 = 32'd9627
; 
32'd185081: dataIn1 = 32'd9628
; 
32'd185082: dataIn1 = 32'd9634
; 
32'd185083: dataIn1 = 32'd2640
; 
32'd185084: dataIn1 = 32'd4912
; 
32'd185085: dataIn1 = 32'd7577
; 
32'd185086: dataIn1 = 32'd9626
; 
32'd185087: dataIn1 = 32'd9627
; 
32'd185088: dataIn1 = 32'd9628
; 
32'd185089: dataIn1 = 32'd9631
; 
32'd185090: dataIn1 = 32'd4912
; 
32'd185091: dataIn1 = 32'd4913
; 
32'd185092: dataIn1 = 32'd4914
; 
32'd185093: dataIn1 = 32'd9626
; 
32'd185094: dataIn1 = 32'd9627
; 
32'd185095: dataIn1 = 32'd9628
; 
32'd185096: dataIn1 = 32'd4688
; 
32'd185097: dataIn1 = 32'd4915
; 
32'd185098: dataIn1 = 32'd7576
; 
32'd185099: dataIn1 = 32'd9603
; 
32'd185100: dataIn1 = 32'd9629
; 
32'd185101: dataIn1 = 32'd9630
; 
32'd185102: dataIn1 = 32'd9631
; 
32'd185103: dataIn1 = 32'd2572
; 
32'd185104: dataIn1 = 32'd4688
; 
32'd185105: dataIn1 = 32'd4912
; 
32'd185106: dataIn1 = 32'd9629
; 
32'd185107: dataIn1 = 32'd9630
; 
32'd185108: dataIn1 = 32'd9631
; 
32'd185109: dataIn1 = 32'd4912
; 
32'd185110: dataIn1 = 32'd4915
; 
32'd185111: dataIn1 = 32'd7577
; 
32'd185112: dataIn1 = 32'd9627
; 
32'd185113: dataIn1 = 32'd9629
; 
32'd185114: dataIn1 = 32'd9630
; 
32'd185115: dataIn1 = 32'd9631
; 
32'd185116: dataIn1 = 32'd2637
; 
32'd185117: dataIn1 = 32'd4909
; 
32'd185118: dataIn1 = 32'd4913
; 
32'd185119: dataIn1 = 32'd9632
; 
32'd185120: dataIn1 = 32'd9633
; 
32'd185121: dataIn1 = 32'd9634
; 
32'd185122: dataIn1 = 32'd4909
; 
32'd185123: dataIn1 = 32'd4916
; 
32'd185124: dataIn1 = 32'd7571
; 
32'd185125: dataIn1 = 32'd9623
; 
32'd185126: dataIn1 = 32'd9632
; 
32'd185127: dataIn1 = 32'd9633
; 
32'd185128: dataIn1 = 32'd9634
; 
32'd185129: dataIn1 = 32'd4913
; 
32'd185130: dataIn1 = 32'd4916
; 
32'd185131: dataIn1 = 32'd7572
; 
32'd185132: dataIn1 = 32'd9626
; 
32'd185133: dataIn1 = 32'd9632
; 
32'd185134: dataIn1 = 32'd9633
; 
32'd185135: dataIn1 = 32'd9634
; 
32'd185136: dataIn1 = 32'd4917
; 
32'd185137: dataIn1 = 32'd4918
; 
32'd185138: dataIn1 = 32'd4919
; 
32'd185139: dataIn1 = 32'd9635
; 
32'd185140: dataIn1 = 32'd9636
; 
32'd185141: dataIn1 = 32'd9637
; 
32'd185142: dataIn1 = 32'd2641
; 
32'd185143: dataIn1 = 32'd4919
; 
32'd185144: dataIn1 = 32'd7604
; 
32'd185145: dataIn1 = 32'd9635
; 
32'd185146: dataIn1 = 32'd9636
; 
32'd185147: dataIn1 = 32'd9637
; 
32'd185148: dataIn1 = 32'd9641
; 
32'd185149: dataIn1 = 32'd2641
; 
32'd185150: dataIn1 = 32'd4918
; 
32'd185151: dataIn1 = 32'd7594
; 
32'd185152: dataIn1 = 32'd9635
; 
32'd185153: dataIn1 = 32'd9636
; 
32'd185154: dataIn1 = 32'd9637
; 
32'd185155: dataIn1 = 32'd9638
; 
32'd185156: dataIn1 = 32'd4918
; 
32'd185157: dataIn1 = 32'd4920
; 
32'd185158: dataIn1 = 32'd7594
; 
32'd185159: dataIn1 = 32'd9637
; 
32'd185160: dataIn1 = 32'd9638
; 
32'd185161: dataIn1 = 32'd9639
; 
32'd185162: dataIn1 = 32'd9640
; 
32'd185163: dataIn1 = 32'd4908
; 
32'd185164: dataIn1 = 32'd4920
; 
32'd185165: dataIn1 = 32'd7593
; 
32'd185166: dataIn1 = 32'd9625
; 
32'd185167: dataIn1 = 32'd9638
; 
32'd185168: dataIn1 = 32'd9639
; 
32'd185169: dataIn1 = 32'd9640
; 
32'd185170: dataIn1 = 32'd2639
; 
32'd185171: dataIn1 = 32'd4908
; 
32'd185172: dataIn1 = 32'd4918
; 
32'd185173: dataIn1 = 32'd9638
; 
32'd185174: dataIn1 = 32'd9639
; 
32'd185175: dataIn1 = 32'd9640
; 
32'd185176: dataIn1 = 32'd4919
; 
32'd185177: dataIn1 = 32'd4921
; 
32'd185178: dataIn1 = 32'd7604
; 
32'd185179: dataIn1 = 32'd9636
; 
32'd185180: dataIn1 = 32'd9641
; 
32'd185181: dataIn1 = 32'd9642
; 
32'd185182: dataIn1 = 32'd9643
; 
32'd185183: dataIn1 = 32'd2576
; 
32'd185184: dataIn1 = 32'd4698
; 
32'd185185: dataIn1 = 32'd4919
; 
32'd185186: dataIn1 = 32'd9641
; 
32'd185187: dataIn1 = 32'd9642
; 
32'd185188: dataIn1 = 32'd9643
; 
32'd185189: dataIn1 = 32'd4698
; 
32'd185190: dataIn1 = 32'd4921
; 
32'd185191: dataIn1 = 32'd7606
; 
32'd185192: dataIn1 = 32'd9607
; 
32'd185193: dataIn1 = 32'd9641
; 
32'd185194: dataIn1 = 32'd9642
; 
32'd185195: dataIn1 = 32'd9643
; 
32'd185196: dataIn1 = 32'd1109
; 
32'd185197: dataIn1 = 32'd4930
; 
32'd185198: dataIn1 = 32'd7747
; 
32'd185199: dataIn1 = 32'd9644
; 
32'd185200: dataIn1 = 32'd9645
; 
32'd185201: dataIn1 = 32'd9646
; 
32'd185202: dataIn1 = 32'd9655
; 
32'd185203: dataIn1 = 32'd1109
; 
32'd185204: dataIn1 = 32'd4929
; 
32'd185205: dataIn1 = 32'd7725
; 
32'd185206: dataIn1 = 32'd9644
; 
32'd185207: dataIn1 = 32'd9645
; 
32'd185208: dataIn1 = 32'd9646
; 
32'd185209: dataIn1 = 32'd9664
; 
32'd185210: dataIn1 = 32'd4924
; 
32'd185211: dataIn1 = 32'd4929
; 
32'd185212: dataIn1 = 32'd4930
; 
32'd185213: dataIn1 = 32'd9644
; 
32'd185214: dataIn1 = 32'd9645
; 
32'd185215: dataIn1 = 32'd9646
; 
32'd185216: dataIn1 = 32'd2645
; 
32'd185217: dataIn1 = 32'd4933
; 
32'd185218: dataIn1 = 32'd7746
; 
32'd185219: dataIn1 = 32'd9647
; 
32'd185220: dataIn1 = 32'd9648
; 
32'd185221: dataIn1 = 32'd9649
; 
32'd185222: dataIn1 = 32'd9654
; 
32'd185223: dataIn1 = 32'd4931
; 
32'd185224: dataIn1 = 32'd4932
; 
32'd185225: dataIn1 = 32'd4933
; 
32'd185226: dataIn1 = 32'd9647
; 
32'd185227: dataIn1 = 32'd9648
; 
32'd185228: dataIn1 = 32'd9649
; 
32'd185229: dataIn1 = 32'd2645
; 
32'd185230: dataIn1 = 32'd4931
; 
32'd185231: dataIn1 = 32'd7741
; 
32'd185232: dataIn1 = 32'd9647
; 
32'd185233: dataIn1 = 32'd9648
; 
32'd185234: dataIn1 = 32'd9649
; 
32'd185235: dataIn1 = 32'd9651
; 
32'd185236: dataIn1 = 32'd4705
; 
32'd185237: dataIn1 = 32'd4934
; 
32'd185238: dataIn1 = 32'd7742
; 
32'd185239: dataIn1 = 32'd9610
; 
32'd185240: dataIn1 = 32'd9650
; 
32'd185241: dataIn1 = 32'd9651
; 
32'd185242: dataIn1 = 32'd9652
; 
32'd185243: dataIn1 = 32'd4931
; 
32'd185244: dataIn1 = 32'd4934
; 
32'd185245: dataIn1 = 32'd7741
; 
32'd185246: dataIn1 = 32'd9649
; 
32'd185247: dataIn1 = 32'd9650
; 
32'd185248: dataIn1 = 32'd9651
; 
32'd185249: dataIn1 = 32'd9652
; 
32'd185250: dataIn1 = 32'd2579
; 
32'd185251: dataIn1 = 32'd4705
; 
32'd185252: dataIn1 = 32'd4931
; 
32'd185253: dataIn1 = 32'd9650
; 
32'd185254: dataIn1 = 32'd9651
; 
32'd185255: dataIn1 = 32'd9652
; 
32'd185256: dataIn1 = 32'd2642
; 
32'd185257: dataIn1 = 32'd4930
; 
32'd185258: dataIn1 = 32'd4933
; 
32'd185259: dataIn1 = 32'd9653
; 
32'd185260: dataIn1 = 32'd9654
; 
32'd185261: dataIn1 = 32'd9655
; 
32'd185262: dataIn1 = 32'd4933
; 
32'd185263: dataIn1 = 32'd4935
; 
32'd185264: dataIn1 = 32'd7746
; 
32'd185265: dataIn1 = 32'd9647
; 
32'd185266: dataIn1 = 32'd9653
; 
32'd185267: dataIn1 = 32'd9654
; 
32'd185268: dataIn1 = 32'd9655
; 
32'd185269: dataIn1 = 32'd4930
; 
32'd185270: dataIn1 = 32'd4935
; 
32'd185271: dataIn1 = 32'd7747
; 
32'd185272: dataIn1 = 32'd9644
; 
32'd185273: dataIn1 = 32'd9653
; 
32'd185274: dataIn1 = 32'd9654
; 
32'd185275: dataIn1 = 32'd9655
; 
32'd185276: dataIn1 = 32'd4936
; 
32'd185277: dataIn1 = 32'd4937
; 
32'd185278: dataIn1 = 32'd4938
; 
32'd185279: dataIn1 = 32'd9656
; 
32'd185280: dataIn1 = 32'd9657
; 
32'd185281: dataIn1 = 32'd9658
; 
32'd185282: dataIn1 = 32'd2646
; 
32'd185283: dataIn1 = 32'd4938
; 
32'd185284: dataIn1 = 32'd7724
; 
32'd185285: dataIn1 = 32'd9656
; 
32'd185286: dataIn1 = 32'd9657
; 
32'd185287: dataIn1 = 32'd9658
; 
32'd185288: dataIn1 = 32'd9662
; 
32'd185289: dataIn1 = 32'd2646
; 
32'd185290: dataIn1 = 32'd4937
; 
32'd185291: dataIn1 = 32'd7714
; 
32'd185292: dataIn1 = 32'd9656
; 
32'd185293: dataIn1 = 32'd9657
; 
32'd185294: dataIn1 = 32'd9658
; 
32'd185295: dataIn1 = 32'd9659
; 
32'd185296: dataIn1 = 32'd4937
; 
32'd185297: dataIn1 = 32'd4939
; 
32'd185298: dataIn1 = 32'd7714
; 
32'd185299: dataIn1 = 32'd9658
; 
32'd185300: dataIn1 = 32'd9659
; 
32'd185301: dataIn1 = 32'd9660
; 
32'd185302: dataIn1 = 32'd9661
; 
32'd185303: dataIn1 = 32'd4699
; 
32'd185304: dataIn1 = 32'd4939
; 
32'd185305: dataIn1 = 32'd7712
; 
32'd185306: dataIn1 = 32'd9605
; 
32'd185307: dataIn1 = 32'd9659
; 
32'd185308: dataIn1 = 32'd9660
; 
32'd185309: dataIn1 = 32'd9661
; 
32'd185310: dataIn1 = 32'd2574
; 
32'd185311: dataIn1 = 32'd4699
; 
32'd185312: dataIn1 = 32'd4937
; 
32'd185313: dataIn1 = 32'd9659
; 
32'd185314: dataIn1 = 32'd9660
; 
32'd185315: dataIn1 = 32'd9661
; 
32'd185316: dataIn1 = 32'd4938
; 
32'd185317: dataIn1 = 32'd4940
; 
32'd185318: dataIn1 = 32'd7724
; 
32'd185319: dataIn1 = 32'd9657
; 
32'd185320: dataIn1 = 32'd9662
; 
32'd185321: dataIn1 = 32'd9663
; 
32'd185322: dataIn1 = 32'd9664
; 
32'd185323: dataIn1 = 32'd2643
; 
32'd185324: dataIn1 = 32'd4929
; 
32'd185325: dataIn1 = 32'd4938
; 
32'd185326: dataIn1 = 32'd9662
; 
32'd185327: dataIn1 = 32'd9663
; 
32'd185328: dataIn1 = 32'd9664
; 
32'd185329: dataIn1 = 32'd4929
; 
32'd185330: dataIn1 = 32'd4940
; 
32'd185331: dataIn1 = 32'd7725
; 
32'd185332: dataIn1 = 32'd9645
; 
32'd185333: dataIn1 = 32'd9662
; 
32'd185334: dataIn1 = 32'd9663
; 
32'd185335: dataIn1 = 32'd9664
; 
32'd185336: dataIn1 = 32'd4706
; 
32'd185337: dataIn1 = 32'd4953
; 
32'd185338: dataIn1 = 32'd7829
; 
32'd185339: dataIn1 = 32'd9609
; 
32'd185340: dataIn1 = 32'd9665
; 
32'd185341: dataIn1 = 32'd9666
; 
32'd185342: dataIn1 = 32'd9667
; 
32'd185343: dataIn1 = 32'd2578
; 
32'd185344: dataIn1 = 32'd4706
; 
32'd185345: dataIn1 = 32'd4950
; 
32'd185346: dataIn1 = 32'd9665
; 
32'd185347: dataIn1 = 32'd9666
; 
32'd185348: dataIn1 = 32'd9667
; 
32'd185349: dataIn1 = 32'd4950
; 
32'd185350: dataIn1 = 32'd4953
; 
32'd185351: dataIn1 = 32'd7830
; 
32'd185352: dataIn1 = 32'd9665
; 
32'd185353: dataIn1 = 32'd9666
; 
32'd185354: dataIn1 = 32'd9667
; 
32'd185355: dataIn1 = 32'd9764
; 
32'd185356: dataIn1 = 32'd2700
; 
32'd185357: dataIn1 = 32'd5142
; 
32'd185358: dataIn1 = 32'd5144
; 
32'd185359: dataIn1 = 32'd6155
; 
32'd185360: dataIn1 = 32'd9668
; 
32'd185361: dataIn1 = 32'd9669
; 
32'd185362: dataIn1 = 32'd10150
; 
32'd185363: dataIn1 = 32'd2700
; 
32'd185364: dataIn1 = 32'd9668
; 
32'd185365: dataIn1 = 32'd9669
; 
32'd185366: dataIn1 = 32'd10119
; 
32'd185367: dataIn1 = 32'd10120
; 
32'd185368: dataIn1 = 32'd10122
; 
32'd185369: dataIn1 = 32'd10150
; 
32'd185370: dataIn1 = 32'd2700
; 
32'd185371: dataIn1 = 32'd9670
; 
32'd185372: dataIn1 = 32'd9671
; 
32'd185373: dataIn1 = 32'd10120
; 
32'd185374: dataIn1 = 32'd10121
; 
32'd185375: dataIn1 = 32'd10125
; 
32'd185376: dataIn1 = 32'd10134
; 
32'd185377: dataIn1 = 32'd2700
; 
32'd185378: dataIn1 = 32'd5269
; 
32'd185379: dataIn1 = 32'd5270
; 
32'd185380: dataIn1 = 32'd6597
; 
32'd185381: dataIn1 = 32'd9670
; 
32'd185382: dataIn1 = 32'd9671
; 
32'd185383: dataIn1 = 32'd10134
; 
32'd185384: dataIn1 = 32'd5451
; 
32'd185385: dataIn1 = 32'd5520
; 
32'd185386: dataIn1 = 32'd6738
; 
32'd185387: dataIn1 = 32'd9672
; 
32'd185388: dataIn1 = 32'd9673
; 
32'd185389: dataIn1 = 32'd10126
; 
32'd185390: dataIn1 = 32'd10132
; 
32'd185391: dataIn1 = 32'd10276
; 
32'd185392: dataIn1 = 32'd10277
; 
32'd185393: dataIn1 = 32'd9672
; 
32'd185394: dataIn1 = 32'd9673
; 
32'd185395: dataIn1 = 32'd10126
; 
32'd185396: dataIn1 = 32'd10127
; 
32'd185397: dataIn1 = 32'd10128
; 
32'd185398: dataIn1 = 32'd10130
; 
32'd185399: dataIn1 = 32'd10132
; 
32'd185400: dataIn1 = 32'd20
; 
32'd185401: dataIn1 = 32'd9674
; 
32'd185402: dataIn1 = 32'd9822
; 
32'd185403: dataIn1 = 32'd9825
; 
32'd185404: dataIn1 = 32'd10129
; 
32'd185405: dataIn1 = 32'd10130
; 
32'd185406: dataIn1 = 32'd10133
; 
32'd185407: dataIn1 = 32'd20
; 
32'd185408: dataIn1 = 32'd6739
; 
32'd185409: dataIn1 = 32'd9675
; 
32'd185410: dataIn1 = 32'd9755
; 
32'd185411: dataIn1 = 32'd10128
; 
32'd185412: dataIn1 = 32'd10129
; 
32'd185413: dataIn1 = 32'd10131
; 
32'd185414: dataIn1 = 32'd1140
; 
32'd185415: dataIn1 = 32'd2111
; 
32'd185416: dataIn1 = 32'd2112
; 
32'd185417: dataIn1 = 32'd5521
; 
32'd185418: dataIn1 = 32'd9452
; 
32'd185419: dataIn1 = 32'd9676
; 
32'd185420: dataIn1 = 32'd124
; 
32'd185421: dataIn1 = 32'd6088
; 
32'd185422: dataIn1 = 32'd9677
; 
32'd185423: dataIn1 = 32'd9678
; 
32'd185424: dataIn1 = 32'd9679
; 
32'd185425: dataIn1 = 32'd9722
; 
32'd185426: dataIn1 = 32'd9724
; 
32'd185427: dataIn1 = 32'd6087
; 
32'd185428: dataIn1 = 32'd6088
; 
32'd185429: dataIn1 = 32'd9677
; 
32'd185430: dataIn1 = 32'd9678
; 
32'd185431: dataIn1 = 32'd9679
; 
32'd185432: dataIn1 = 32'd9792
; 
32'd185433: dataIn1 = 32'd9793
; 
32'd185434: dataIn1 = 32'd124
; 
32'd185435: dataIn1 = 32'd6087
; 
32'd185436: dataIn1 = 32'd9677
; 
32'd185437: dataIn1 = 32'd9678
; 
32'd185438: dataIn1 = 32'd9679
; 
32'd185439: dataIn1 = 32'd9701
; 
32'd185440: dataIn1 = 32'd9704
; 
32'd185441: dataIn1 = 32'd1102
; 
32'd185442: dataIn1 = 32'd6105
; 
32'd185443: dataIn1 = 32'd9680
; 
32'd185444: dataIn1 = 32'd9681
; 
32'd185445: dataIn1 = 32'd9682
; 
32'd185446: dataIn1 = 32'd9694
; 
32'd185447: dataIn1 = 32'd9696
; 
32'd185448: dataIn1 = 32'd1102
; 
32'd185449: dataIn1 = 32'd6104
; 
32'd185450: dataIn1 = 32'd9680
; 
32'd185451: dataIn1 = 32'd9681
; 
32'd185452: dataIn1 = 32'd9682
; 
32'd185453: dataIn1 = 32'd9707
; 
32'd185454: dataIn1 = 32'd9709
; 
32'd185455: dataIn1 = 32'd6104
; 
32'd185456: dataIn1 = 32'd6105
; 
32'd185457: dataIn1 = 32'd9680
; 
32'd185458: dataIn1 = 32'd9681
; 
32'd185459: dataIn1 = 32'd9682
; 
32'd185460: dataIn1 = 32'd9800
; 
32'd185461: dataIn1 = 32'd9801
; 
32'd185462: dataIn1 = 32'd2611
; 
32'd185463: dataIn1 = 32'd6108
; 
32'd185464: dataIn1 = 32'd9683
; 
32'd185465: dataIn1 = 32'd9684
; 
32'd185466: dataIn1 = 32'd9685
; 
32'd185467: dataIn1 = 32'd9693
; 
32'd185468: dataIn1 = 32'd9695
; 
32'd185469: dataIn1 = 32'd6106
; 
32'd185470: dataIn1 = 32'd6108
; 
32'd185471: dataIn1 = 32'd9683
; 
32'd185472: dataIn1 = 32'd9684
; 
32'd185473: dataIn1 = 32'd9685
; 
32'd185474: dataIn1 = 32'd9804
; 
32'd185475: dataIn1 = 32'd9805
; 
32'd185476: dataIn1 = 32'd2611
; 
32'd185477: dataIn1 = 32'd6106
; 
32'd185478: dataIn1 = 32'd9683
; 
32'd185479: dataIn1 = 32'd9684
; 
32'd185480: dataIn1 = 32'd9685
; 
32'd185481: dataIn1 = 32'd9687
; 
32'd185482: dataIn1 = 32'd9691
; 
32'd185483: dataIn1 = 32'd4803
; 
32'd185484: dataIn1 = 32'd6109
; 
32'd185485: dataIn1 = 32'd9686
; 
32'd185486: dataIn1 = 32'd9687
; 
32'd185487: dataIn1 = 32'd9688
; 
32'd185488: dataIn1 = 32'd9689
; 
32'd185489: dataIn1 = 32'd9690
; 
32'd185490: dataIn1 = 32'd4803
; 
32'd185491: dataIn1 = 32'd6106
; 
32'd185492: dataIn1 = 32'd9685
; 
32'd185493: dataIn1 = 32'd9686
; 
32'd185494: dataIn1 = 32'd9687
; 
32'd185495: dataIn1 = 32'd9688
; 
32'd185496: dataIn1 = 32'd9691
; 
32'd185497: dataIn1 = 32'd6106
; 
32'd185498: dataIn1 = 32'd6109
; 
32'd185499: dataIn1 = 32'd9686
; 
32'd185500: dataIn1 = 32'd9687
; 
32'd185501: dataIn1 = 32'd9688
; 
32'd185502: dataIn1 = 32'd9806
; 
32'd185503: dataIn1 = 32'd9807
; 
32'd185504: dataIn1 = 32'd3
; 
32'd185505: dataIn1 = 32'd4638
; 
32'd185506: dataIn1 = 32'd4803
; 
32'd185507: dataIn1 = 32'd9686
; 
32'd185508: dataIn1 = 32'd9689
; 
32'd185509: dataIn1 = 32'd9690
; 
32'd185510: dataIn1 = 32'd3
; 
32'd185511: dataIn1 = 32'd6109
; 
32'd185512: dataIn1 = 32'd9686
; 
32'd185513: dataIn1 = 32'd9689
; 
32'd185514: dataIn1 = 32'd9690
; 
32'd185515: dataIn1 = 32'd9756
; 
32'd185516: dataIn1 = 32'd9757
; 
32'd185517: dataIn1 = 32'd2611
; 
32'd185518: dataIn1 = 32'd4801
; 
32'd185519: dataIn1 = 32'd4803
; 
32'd185520: dataIn1 = 32'd9685
; 
32'd185521: dataIn1 = 32'd9687
; 
32'd185522: dataIn1 = 32'd9691
; 
32'd185523: dataIn1 = 32'd6105
; 
32'd185524: dataIn1 = 32'd6108
; 
32'd185525: dataIn1 = 32'd9692
; 
32'd185526: dataIn1 = 32'd9693
; 
32'd185527: dataIn1 = 32'd9694
; 
32'd185528: dataIn1 = 32'd9802
; 
32'd185529: dataIn1 = 32'd9803
; 
32'd185530: dataIn1 = 32'd4804
; 
32'd185531: dataIn1 = 32'd6108
; 
32'd185532: dataIn1 = 32'd9683
; 
32'd185533: dataIn1 = 32'd9692
; 
32'd185534: dataIn1 = 32'd9693
; 
32'd185535: dataIn1 = 32'd9694
; 
32'd185536: dataIn1 = 32'd9695
; 
32'd185537: dataIn1 = 32'd4804
; 
32'd185538: dataIn1 = 32'd6105
; 
32'd185539: dataIn1 = 32'd9680
; 
32'd185540: dataIn1 = 32'd9692
; 
32'd185541: dataIn1 = 32'd9693
; 
32'd185542: dataIn1 = 32'd9694
; 
32'd185543: dataIn1 = 32'd9696
; 
32'd185544: dataIn1 = 32'd2611
; 
32'd185545: dataIn1 = 32'd4802
; 
32'd185546: dataIn1 = 32'd4804
; 
32'd185547: dataIn1 = 32'd9683
; 
32'd185548: dataIn1 = 32'd9693
; 
32'd185549: dataIn1 = 32'd9695
; 
32'd185550: dataIn1 = 32'd1102
; 
32'd185551: dataIn1 = 32'd4792
; 
32'd185552: dataIn1 = 32'd4804
; 
32'd185553: dataIn1 = 32'd9680
; 
32'd185554: dataIn1 = 32'd9694
; 
32'd185555: dataIn1 = 32'd9696
; 
32'd185556: dataIn1 = 32'd6112
; 
32'd185557: dataIn1 = 32'd6113
; 
32'd185558: dataIn1 = 32'd9697
; 
32'd185559: dataIn1 = 32'd9698
; 
32'd185560: dataIn1 = 32'd9699
; 
32'd185561: dataIn1 = 32'd9796
; 
32'd185562: dataIn1 = 32'd9797
; 
32'd185563: dataIn1 = 32'd2610
; 
32'd185564: dataIn1 = 32'd6113
; 
32'd185565: dataIn1 = 32'd9697
; 
32'd185566: dataIn1 = 32'd9698
; 
32'd185567: dataIn1 = 32'd9699
; 
32'd185568: dataIn1 = 32'd9705
; 
32'd185569: dataIn1 = 32'd9708
; 
32'd185570: dataIn1 = 32'd2610
; 
32'd185571: dataIn1 = 32'd6112
; 
32'd185572: dataIn1 = 32'd9697
; 
32'd185573: dataIn1 = 32'd9698
; 
32'd185574: dataIn1 = 32'd9699
; 
32'd185575: dataIn1 = 32'd9700
; 
32'd185576: dataIn1 = 32'd9703
; 
32'd185577: dataIn1 = 32'd4798
; 
32'd185578: dataIn1 = 32'd6112
; 
32'd185579: dataIn1 = 32'd9699
; 
32'd185580: dataIn1 = 32'd9700
; 
32'd185581: dataIn1 = 32'd9701
; 
32'd185582: dataIn1 = 32'd9702
; 
32'd185583: dataIn1 = 32'd9703
; 
32'd185584: dataIn1 = 32'd4798
; 
32'd185585: dataIn1 = 32'd6087
; 
32'd185586: dataIn1 = 32'd9679
; 
32'd185587: dataIn1 = 32'd9700
; 
32'd185588: dataIn1 = 32'd9701
; 
32'd185589: dataIn1 = 32'd9702
; 
32'd185590: dataIn1 = 32'd9704
; 
32'd185591: dataIn1 = 32'd6087
; 
32'd185592: dataIn1 = 32'd6112
; 
32'd185593: dataIn1 = 32'd9700
; 
32'd185594: dataIn1 = 32'd9701
; 
32'd185595: dataIn1 = 32'd9702
; 
32'd185596: dataIn1 = 32'd9794
; 
32'd185597: dataIn1 = 32'd9795
; 
32'd185598: dataIn1 = 32'd2610
; 
32'd185599: dataIn1 = 32'd4795
; 
32'd185600: dataIn1 = 32'd4798
; 
32'd185601: dataIn1 = 32'd9699
; 
32'd185602: dataIn1 = 32'd9700
; 
32'd185603: dataIn1 = 32'd9703
; 
32'd185604: dataIn1 = 32'd124
; 
32'd185605: dataIn1 = 32'd4640
; 
32'd185606: dataIn1 = 32'd4798
; 
32'd185607: dataIn1 = 32'd9679
; 
32'd185608: dataIn1 = 32'd9701
; 
32'd185609: dataIn1 = 32'd9704
; 
32'd185610: dataIn1 = 32'd4799
; 
32'd185611: dataIn1 = 32'd6113
; 
32'd185612: dataIn1 = 32'd9698
; 
32'd185613: dataIn1 = 32'd9705
; 
32'd185614: dataIn1 = 32'd9706
; 
32'd185615: dataIn1 = 32'd9707
; 
32'd185616: dataIn1 = 32'd9708
; 
32'd185617: dataIn1 = 32'd6104
; 
32'd185618: dataIn1 = 32'd6113
; 
32'd185619: dataIn1 = 32'd9705
; 
32'd185620: dataIn1 = 32'd9706
; 
32'd185621: dataIn1 = 32'd9707
; 
32'd185622: dataIn1 = 32'd9798
; 
32'd185623: dataIn1 = 32'd9799
; 
32'd185624: dataIn1 = 32'd4799
; 
32'd185625: dataIn1 = 32'd6104
; 
32'd185626: dataIn1 = 32'd9681
; 
32'd185627: dataIn1 = 32'd9705
; 
32'd185628: dataIn1 = 32'd9706
; 
32'd185629: dataIn1 = 32'd9707
; 
32'd185630: dataIn1 = 32'd9709
; 
32'd185631: dataIn1 = 32'd2610
; 
32'd185632: dataIn1 = 32'd4797
; 
32'd185633: dataIn1 = 32'd4799
; 
32'd185634: dataIn1 = 32'd9698
; 
32'd185635: dataIn1 = 32'd9705
; 
32'd185636: dataIn1 = 32'd9708
; 
32'd185637: dataIn1 = 32'd1102
; 
32'd185638: dataIn1 = 32'd4793
; 
32'd185639: dataIn1 = 32'd4799
; 
32'd185640: dataIn1 = 32'd9681
; 
32'd185641: dataIn1 = 32'd9707
; 
32'd185642: dataIn1 = 32'd9709
; 
32'd185643: dataIn1 = 32'd6122
; 
32'd185644: dataIn1 = 32'd6123
; 
32'd185645: dataIn1 = 32'd9710
; 
32'd185646: dataIn1 = 32'd9711
; 
32'd185647: dataIn1 = 32'd9712
; 
32'd185648: dataIn1 = 32'd9777
; 
32'd185649: dataIn1 = 32'd9785
; 
32'd185650: dataIn1 = 32'd1103
; 
32'd185651: dataIn1 = 32'd6123
; 
32'd185652: dataIn1 = 32'd9710
; 
32'd185653: dataIn1 = 32'd9711
; 
32'd185654: dataIn1 = 32'd9712
; 
32'd185655: dataIn1 = 32'd9716
; 
32'd185656: dataIn1 = 32'd9719
; 
32'd185657: dataIn1 = 32'd1103
; 
32'd185658: dataIn1 = 32'd6122
; 
32'd185659: dataIn1 = 32'd9710
; 
32'd185660: dataIn1 = 32'd9711
; 
32'd185661: dataIn1 = 32'd9712
; 
32'd185662: dataIn1 = 32'd9726
; 
32'd185663: dataIn1 = 32'd9729
; 
32'd185664: dataIn1 = 32'd2615
; 
32'd185665: dataIn1 = 32'd6134
; 
32'd185666: dataIn1 = 32'd9713
; 
32'd185667: dataIn1 = 32'd9714
; 
32'd185668: dataIn1 = 32'd9715
; 
32'd185669: dataIn1 = 32'd9723
; 
32'd185670: dataIn1 = 32'd9725
; 
32'd185671: dataIn1 = 32'd2615
; 
32'd185672: dataIn1 = 32'd6133
; 
32'd185673: dataIn1 = 32'd9713
; 
32'd185674: dataIn1 = 32'd9714
; 
32'd185675: dataIn1 = 32'd9715
; 
32'd185676: dataIn1 = 32'd9718
; 
32'd185677: dataIn1 = 32'd9720
; 
32'd185678: dataIn1 = 32'd6133
; 
32'd185679: dataIn1 = 32'd6134
; 
32'd185680: dataIn1 = 32'd9713
; 
32'd185681: dataIn1 = 32'd9714
; 
32'd185682: dataIn1 = 32'd9715
; 
32'd185683: dataIn1 = 32'd9788
; 
32'd185684: dataIn1 = 32'd9789
; 
32'd185685: dataIn1 = 32'd4812
; 
32'd185686: dataIn1 = 32'd6123
; 
32'd185687: dataIn1 = 32'd9711
; 
32'd185688: dataIn1 = 32'd9716
; 
32'd185689: dataIn1 = 32'd9717
; 
32'd185690: dataIn1 = 32'd9718
; 
32'd185691: dataIn1 = 32'd9719
; 
32'd185692: dataIn1 = 32'd6123
; 
32'd185693: dataIn1 = 32'd6133
; 
32'd185694: dataIn1 = 32'd9716
; 
32'd185695: dataIn1 = 32'd9717
; 
32'd185696: dataIn1 = 32'd9718
; 
32'd185697: dataIn1 = 32'd9786
; 
32'd185698: dataIn1 = 32'd9787
; 
32'd185699: dataIn1 = 32'd4812
; 
32'd185700: dataIn1 = 32'd6133
; 
32'd185701: dataIn1 = 32'd9714
; 
32'd185702: dataIn1 = 32'd9716
; 
32'd185703: dataIn1 = 32'd9717
; 
32'd185704: dataIn1 = 32'd9718
; 
32'd185705: dataIn1 = 32'd9720
; 
32'd185706: dataIn1 = 32'd1103
; 
32'd185707: dataIn1 = 32'd4807
; 
32'd185708: dataIn1 = 32'd4812
; 
32'd185709: dataIn1 = 32'd9711
; 
32'd185710: dataIn1 = 32'd9716
; 
32'd185711: dataIn1 = 32'd9719
; 
32'd185712: dataIn1 = 32'd2615
; 
32'd185713: dataIn1 = 32'd4809
; 
32'd185714: dataIn1 = 32'd4812
; 
32'd185715: dataIn1 = 32'd9714
; 
32'd185716: dataIn1 = 32'd9718
; 
32'd185717: dataIn1 = 32'd9720
; 
32'd185718: dataIn1 = 32'd6088
; 
32'd185719: dataIn1 = 32'd6134
; 
32'd185720: dataIn1 = 32'd9721
; 
32'd185721: dataIn1 = 32'd9722
; 
32'd185722: dataIn1 = 32'd9723
; 
32'd185723: dataIn1 = 32'd9790
; 
32'd185724: dataIn1 = 32'd9791
; 
32'd185725: dataIn1 = 32'd4811
; 
32'd185726: dataIn1 = 32'd6088
; 
32'd185727: dataIn1 = 32'd9677
; 
32'd185728: dataIn1 = 32'd9721
; 
32'd185729: dataIn1 = 32'd9722
; 
32'd185730: dataIn1 = 32'd9723
; 
32'd185731: dataIn1 = 32'd9724
; 
32'd185732: dataIn1 = 32'd4811
; 
32'd185733: dataIn1 = 32'd6134
; 
32'd185734: dataIn1 = 32'd9713
; 
32'd185735: dataIn1 = 32'd9721
; 
32'd185736: dataIn1 = 32'd9722
; 
32'd185737: dataIn1 = 32'd9723
; 
32'd185738: dataIn1 = 32'd9725
; 
32'd185739: dataIn1 = 32'd124
; 
32'd185740: dataIn1 = 32'd4641
; 
32'd185741: dataIn1 = 32'd4811
; 
32'd185742: dataIn1 = 32'd9677
; 
32'd185743: dataIn1 = 32'd9722
; 
32'd185744: dataIn1 = 32'd9724
; 
32'd185745: dataIn1 = 32'd2615
; 
32'd185746: dataIn1 = 32'd4808
; 
32'd185747: dataIn1 = 32'd4811
; 
32'd185748: dataIn1 = 32'd9713
; 
32'd185749: dataIn1 = 32'd9723
; 
32'd185750: dataIn1 = 32'd9725
; 
32'd185751: dataIn1 = 32'd4816
; 
32'd185752: dataIn1 = 32'd6122
; 
32'd185753: dataIn1 = 32'd9712
; 
32'd185754: dataIn1 = 32'd9726
; 
32'd185755: dataIn1 = 32'd9727
; 
32'd185756: dataIn1 = 32'd9728
; 
32'd185757: dataIn1 = 32'd9729
; 
32'd185758: dataIn1 = 32'd4816
; 
32'd185759: dataIn1 = 32'd6136
; 
32'd185760: dataIn1 = 32'd9726
; 
32'd185761: dataIn1 = 32'd9727
; 
32'd185762: dataIn1 = 32'd9728
; 
32'd185763: dataIn1 = 32'd9730
; 
32'd185764: dataIn1 = 32'd9731
; 
32'd185765: dataIn1 = 32'd6122
; 
32'd185766: dataIn1 = 32'd6136
; 
32'd185767: dataIn1 = 32'd7214
; 
32'd185768: dataIn1 = 32'd9726
; 
32'd185769: dataIn1 = 32'd9727
; 
32'd185770: dataIn1 = 32'd9728
; 
32'd185771: dataIn1 = 32'd9759
; 
32'd185772: dataIn1 = 32'd1103
; 
32'd185773: dataIn1 = 32'd4805
; 
32'd185774: dataIn1 = 32'd4816
; 
32'd185775: dataIn1 = 32'd9712
; 
32'd185776: dataIn1 = 32'd9726
; 
32'd185777: dataIn1 = 32'd9729
; 
32'd185778: dataIn1 = 32'd2616
; 
32'd185779: dataIn1 = 32'd4814
; 
32'd185780: dataIn1 = 32'd4816
; 
32'd185781: dataIn1 = 32'd9727
; 
32'd185782: dataIn1 = 32'd9730
; 
32'd185783: dataIn1 = 32'd9731
; 
32'd185784: dataIn1 = 32'd2616
; 
32'd185785: dataIn1 = 32'd6136
; 
32'd185786: dataIn1 = 32'd7209
; 
32'd185787: dataIn1 = 32'd9727
; 
32'd185788: dataIn1 = 32'd9730
; 
32'd185789: dataIn1 = 32'd9731
; 
32'd185790: dataIn1 = 32'd9758
; 
32'd185791: dataIn1 = 32'd6155
; 
32'd185792: dataIn1 = 32'd6156
; 
32'd185793: dataIn1 = 32'd7250
; 
32'd185794: dataIn1 = 32'd9732
; 
32'd185795: dataIn1 = 32'd9733
; 
32'd185796: dataIn1 = 32'd9734
; 
32'd185797: dataIn1 = 32'd9760
; 
32'd185798: dataIn1 = 32'd6154
; 
32'd185799: dataIn1 = 32'd6156
; 
32'd185800: dataIn1 = 32'd7252
; 
32'd185801: dataIn1 = 32'd9732
; 
32'd185802: dataIn1 = 32'd9733
; 
32'd185803: dataIn1 = 32'd9734
; 
32'd185804: dataIn1 = 32'd9761
; 
32'd185805: dataIn1 = 32'd5142
; 
32'd185806: dataIn1 = 32'd6154
; 
32'd185807: dataIn1 = 32'd6155
; 
32'd185808: dataIn1 = 32'd9732
; 
32'd185809: dataIn1 = 32'd9733
; 
32'd185810: dataIn1 = 32'd9734
; 
32'd185811: dataIn1 = 32'd6393
; 
32'd185812: dataIn1 = 32'd6394
; 
32'd185813: dataIn1 = 32'd8139
; 
32'd185814: dataIn1 = 32'd9735
; 
32'd185815: dataIn1 = 32'd9736
; 
32'd185816: dataIn1 = 32'd9737
; 
32'd185817: dataIn1 = 32'd9765
; 
32'd185818: dataIn1 = 32'd6392
; 
32'd185819: dataIn1 = 32'd6394
; 
32'd185820: dataIn1 = 32'd8140
; 
32'd185821: dataIn1 = 32'd9735
; 
32'd185822: dataIn1 = 32'd9736
; 
32'd185823: dataIn1 = 32'd9737
; 
32'd185824: dataIn1 = 32'd9766
; 
32'd185825: dataIn1 = 32'd6392
; 
32'd185826: dataIn1 = 32'd6393
; 
32'd185827: dataIn1 = 32'd9735
; 
32'd185828: dataIn1 = 32'd9736
; 
32'd185829: dataIn1 = 32'd9737
; 
32'd185830: dataIn1 = 32'd9738
; 
32'd185831: dataIn1 = 32'd9739
; 
32'd185832: dataIn1 = 32'd5211
; 
32'd185833: dataIn1 = 32'd6393
; 
32'd185834: dataIn1 = 32'd6397
; 
32'd185835: dataIn1 = 32'd9737
; 
32'd185836: dataIn1 = 32'd9738
; 
32'd185837: dataIn1 = 32'd9739
; 
32'd185838: dataIn1 = 32'd5211
; 
32'd185839: dataIn1 = 32'd6392
; 
32'd185840: dataIn1 = 32'd9737
; 
32'd185841: dataIn1 = 32'd9738
; 
32'd185842: dataIn1 = 32'd9739
; 
32'd185843: dataIn1 = 32'd9740
; 
32'd185844: dataIn1 = 32'd9741
; 
32'd185845: dataIn1 = 32'd5211
; 
32'd185846: dataIn1 = 32'd6395
; 
32'd185847: dataIn1 = 32'd9739
; 
32'd185848: dataIn1 = 32'd9740
; 
32'd185849: dataIn1 = 32'd9741
; 
32'd185850: dataIn1 = 32'd10140
; 
32'd185851: dataIn1 = 32'd10221
; 
32'd185852: dataIn1 = 32'd6392
; 
32'd185853: dataIn1 = 32'd6395
; 
32'd185854: dataIn1 = 32'd9739
; 
32'd185855: dataIn1 = 32'd9740
; 
32'd185856: dataIn1 = 32'd9741
; 
32'd185857: dataIn1 = 32'd10279
; 
32'd185858: dataIn1 = 32'd10282
; 
32'd185859: dataIn1 = 32'd5269
; 
32'd185860: dataIn1 = 32'd6596
; 
32'd185861: dataIn1 = 32'd6597
; 
32'd185862: dataIn1 = 32'd9742
; 
32'd185863: dataIn1 = 32'd9743
; 
32'd185864: dataIn1 = 32'd9744
; 
32'd185865: dataIn1 = 32'd6595
; 
32'd185866: dataIn1 = 32'd6597
; 
32'd185867: dataIn1 = 32'd9742
; 
32'd185868: dataIn1 = 32'd9743
; 
32'd185869: dataIn1 = 32'd9744
; 
32'd185870: dataIn1 = 32'd9745
; 
32'd185871: dataIn1 = 32'd9746
; 
32'd185872: dataIn1 = 32'd6595
; 
32'd185873: dataIn1 = 32'd6596
; 
32'd185874: dataIn1 = 32'd8926
; 
32'd185875: dataIn1 = 32'd9742
; 
32'd185876: dataIn1 = 32'd9743
; 
32'd185877: dataIn1 = 32'd9744
; 
32'd185878: dataIn1 = 32'd9768
; 
32'd185879: dataIn1 = 32'd5143
; 
32'd185880: dataIn1 = 32'd6597
; 
32'd185881: dataIn1 = 32'd9743
; 
32'd185882: dataIn1 = 32'd9745
; 
32'd185883: dataIn1 = 32'd9746
; 
32'd185884: dataIn1 = 32'd10125
; 
32'd185885: dataIn1 = 32'd10134
; 
32'd185886: dataIn1 = 32'd5143
; 
32'd185887: dataIn1 = 32'd6595
; 
32'd185888: dataIn1 = 32'd8922
; 
32'd185889: dataIn1 = 32'd9743
; 
32'd185890: dataIn1 = 32'd9745
; 
32'd185891: dataIn1 = 32'd9746
; 
32'd185892: dataIn1 = 32'd9767
; 
32'd185893: dataIn1 = 32'd9747
; 
32'd185894: dataIn1 = 32'd9748
; 
32'd185895: dataIn1 = 32'd10136
; 
32'd185896: dataIn1 = 32'd10137
; 
32'd185897: dataIn1 = 32'd10139
; 
32'd185898: dataIn1 = 32'd10140
; 
32'd185899: dataIn1 = 32'd10221
; 
32'd185900: dataIn1 = 32'd5211
; 
32'd185901: dataIn1 = 32'd6397
; 
32'd185902: dataIn1 = 32'd6712
; 
32'd185903: dataIn1 = 32'd9747
; 
32'd185904: dataIn1 = 32'd9748
; 
32'd185905: dataIn1 = 32'd9749
; 
32'd185906: dataIn1 = 32'd9776
; 
32'd185907: dataIn1 = 32'd10136
; 
32'd185908: dataIn1 = 32'd10221
; 
32'd185909: dataIn1 = 32'd6712
; 
32'd185910: dataIn1 = 32'd9748
; 
32'd185911: dataIn1 = 32'd9749
; 
32'd185912: dataIn1 = 32'd9752
; 
32'd185913: dataIn1 = 32'd10135
; 
32'd185914: dataIn1 = 32'd10136
; 
32'd185915: dataIn1 = 32'd10142
; 
32'd185916: dataIn1 = 32'd1129
; 
32'd185917: dataIn1 = 32'd9750
; 
32'd185918: dataIn1 = 32'd10138
; 
32'd185919: dataIn1 = 32'd10139
; 
32'd185920: dataIn1 = 32'd10141
; 
32'd185921: dataIn1 = 32'd10222
; 
32'd185922: dataIn1 = 32'd10223
; 
32'd185923: dataIn1 = 32'd9751
; 
32'd185924: dataIn1 = 32'd9752
; 
32'd185925: dataIn1 = 32'd10142
; 
32'd185926: dataIn1 = 32'd10143
; 
32'd185927: dataIn1 = 32'd10144
; 
32'd185928: dataIn1 = 32'd10145
; 
32'd185929: dataIn1 = 32'd10147
; 
32'd185930: dataIn1 = 32'd5440
; 
32'd185931: dataIn1 = 32'd6712
; 
32'd185932: dataIn1 = 32'd6739
; 
32'd185933: dataIn1 = 32'd9749
; 
32'd185934: dataIn1 = 32'd9751
; 
32'd185935: dataIn1 = 32'd9752
; 
32'd185936: dataIn1 = 32'd10142
; 
32'd185937: dataIn1 = 32'd10147
; 
32'd185938: dataIn1 = 32'd6738
; 
32'd185939: dataIn1 = 32'd9753
; 
32'd185940: dataIn1 = 32'd10145
; 
32'd185941: dataIn1 = 32'd10146
; 
32'd185942: dataIn1 = 32'd10149
; 
32'd185943: dataIn1 = 32'd10223
; 
32'd185944: dataIn1 = 32'd10224
; 
32'd185945: dataIn1 = 32'd6738
; 
32'd185946: dataIn1 = 32'd9754
; 
32'd185947: dataIn1 = 32'd10126
; 
32'd185948: dataIn1 = 32'd10127
; 
32'd185949: dataIn1 = 32'd10144
; 
32'd185950: dataIn1 = 32'd10146
; 
32'd185951: dataIn1 = 32'd10148
; 
32'd185952: dataIn1 = 32'd20
; 
32'd185953: dataIn1 = 32'd5439
; 
32'd185954: dataIn1 = 32'd5521
; 
32'd185955: dataIn1 = 32'd6739
; 
32'd185956: dataIn1 = 32'd9675
; 
32'd185957: dataIn1 = 32'd9755
; 
32'd185958: dataIn1 = 32'd6109
; 
32'd185959: dataIn1 = 32'd6814
; 
32'd185960: dataIn1 = 32'd9690
; 
32'd185961: dataIn1 = 32'd9756
; 
32'd185962: dataIn1 = 32'd9757
; 
32'd185963: dataIn1 = 32'd9808
; 
32'd185964: dataIn1 = 32'd9809
; 
32'd185965: dataIn1 = 32'd3
; 
32'd185966: dataIn1 = 32'd6814
; 
32'd185967: dataIn1 = 32'd9690
; 
32'd185968: dataIn1 = 32'd9756
; 
32'd185969: dataIn1 = 32'd9757
; 
32'd185970: dataIn1 = 32'd2616
; 
32'd185971: dataIn1 = 32'd4817
; 
32'd185972: dataIn1 = 32'd6138
; 
32'd185973: dataIn1 = 32'd7209
; 
32'd185974: dataIn1 = 32'd9731
; 
32'd185975: dataIn1 = 32'd9758
; 
32'd185976: dataIn1 = 32'd5128
; 
32'd185977: dataIn1 = 32'd6122
; 
32'd185978: dataIn1 = 32'd7171
; 
32'd185979: dataIn1 = 32'd7214
; 
32'd185980: dataIn1 = 32'd9728
; 
32'd185981: dataIn1 = 32'd9759
; 
32'd185982: dataIn1 = 32'd9777
; 
32'd185983: dataIn1 = 32'd5140
; 
32'd185984: dataIn1 = 32'd6155
; 
32'd185985: dataIn1 = 32'd7250
; 
32'd185986: dataIn1 = 32'd9732
; 
32'd185987: dataIn1 = 32'd9760
; 
32'd185988: dataIn1 = 32'd10122
; 
32'd185989: dataIn1 = 32'd10150
; 
32'd185990: dataIn1 = 32'd5141
; 
32'd185991: dataIn1 = 32'd6154
; 
32'd185992: dataIn1 = 32'd7252
; 
32'd185993: dataIn1 = 32'd7275
; 
32'd185994: dataIn1 = 32'd9733
; 
32'd185995: dataIn1 = 32'd9761
; 
32'd185996: dataIn1 = 32'd9762
; 
32'd185997: dataIn1 = 32'd6154
; 
32'd185998: dataIn1 = 32'd6157
; 
32'd185999: dataIn1 = 32'd6158
; 
32'd186000: dataIn1 = 32'd7275
; 
32'd186001: dataIn1 = 32'd9761
; 
32'd186002: dataIn1 = 32'd9762
; 
32'd186003: dataIn1 = 32'd4891
; 
32'd186004: dataIn1 = 32'd4900
; 
32'd186005: dataIn1 = 32'd4902
; 
32'd186006: dataIn1 = 32'd7472
; 
32'd186007: dataIn1 = 32'd9612
; 
32'd186008: dataIn1 = 32'd9763
; 
32'd186009: dataIn1 = 32'd2650
; 
32'd186010: dataIn1 = 32'd4950
; 
32'd186011: dataIn1 = 32'd4951
; 
32'd186012: dataIn1 = 32'd7830
; 
32'd186013: dataIn1 = 32'd9667
; 
32'd186014: dataIn1 = 32'd9764
; 
32'd186015: dataIn1 = 32'd5207
; 
32'd186016: dataIn1 = 32'd6389
; 
32'd186017: dataIn1 = 32'd6393
; 
32'd186018: dataIn1 = 32'd8139
; 
32'd186019: dataIn1 = 32'd9735
; 
32'd186020: dataIn1 = 32'd9765
; 
32'd186021: dataIn1 = 32'd5210
; 
32'd186022: dataIn1 = 32'd6392
; 
32'd186023: dataIn1 = 32'd8140
; 
32'd186024: dataIn1 = 32'd9736
; 
32'd186025: dataIn1 = 32'd9766
; 
32'd186026: dataIn1 = 32'd10278
; 
32'd186027: dataIn1 = 32'd10279
; 
32'd186028: dataIn1 = 32'd5143
; 
32'd186029: dataIn1 = 32'd6164
; 
32'd186030: dataIn1 = 32'd7258
; 
32'd186031: dataIn1 = 32'd8922
; 
32'd186032: dataIn1 = 32'd9746
; 
32'd186033: dataIn1 = 32'd9767
; 
32'd186034: dataIn1 = 32'd9778
; 
32'd186035: dataIn1 = 32'd3985
; 
32'd186036: dataIn1 = 32'd6596
; 
32'd186037: dataIn1 = 32'd7050
; 
32'd186038: dataIn1 = 32'd8926
; 
32'd186039: dataIn1 = 32'd9744
; 
32'd186040: dataIn1 = 32'd9768
; 
32'd186041: dataIn1 = 32'd9779
; 
32'd186042: dataIn1 = 32'd42
; 
32'd186043: dataIn1 = 32'd2149
; 
32'd186044: dataIn1 = 32'd2150
; 
32'd186045: dataIn1 = 32'd9461
; 
32'd186046: dataIn1 = 32'd9477
; 
32'd186047: dataIn1 = 32'd9769
; 
32'd186048: dataIn1 = 32'd2175
; 
32'd186049: dataIn1 = 32'd9770
; 
32'd186050: dataIn1 = 32'd9771
; 
32'd186051: dataIn1 = 32'd9781
; 
32'd186052: dataIn1 = 32'd10160
; 
32'd186053: dataIn1 = 32'd10161
; 
32'd186054: dataIn1 = 32'd10227
; 
32'd186055: dataIn1 = 32'd2175
; 
32'd186056: dataIn1 = 32'd2176
; 
32'd186057: dataIn1 = 32'd3589
; 
32'd186058: dataIn1 = 32'd3631
; 
32'd186059: dataIn1 = 32'd9471
; 
32'd186060: dataIn1 = 32'd9770
; 
32'd186061: dataIn1 = 32'd9771
; 
32'd186062: dataIn1 = 32'd9780
; 
32'd186063: dataIn1 = 32'd10160
; 
32'd186064: dataIn1 = 32'd2218
; 
32'd186065: dataIn1 = 32'd9772
; 
32'd186066: dataIn1 = 32'd9783
; 
32'd186067: dataIn1 = 32'd10205
; 
32'd186068: dataIn1 = 32'd10206
; 
32'd186069: dataIn1 = 32'd10238
; 
32'd186070: dataIn1 = 32'd10239
; 
32'd186071: dataIn1 = 32'd2218
; 
32'd186072: dataIn1 = 32'd5310
; 
32'd186073: dataIn1 = 32'd9773
; 
32'd186074: dataIn1 = 32'd9782
; 
32'd186075: dataIn1 = 32'd10203
; 
32'd186076: dataIn1 = 32'd10204
; 
32'd186077: dataIn1 = 32'd10238
; 
32'd186078: dataIn1 = 32'd2219
; 
32'd186079: dataIn1 = 32'd9774
; 
32'd186080: dataIn1 = 32'd9783
; 
32'd186081: dataIn1 = 32'd10207
; 
32'd186082: dataIn1 = 32'd10208
; 
32'd186083: dataIn1 = 32'd10239
; 
32'd186084: dataIn1 = 32'd10240
; 
32'd186085: dataIn1 = 32'd2219
; 
32'd186086: dataIn1 = 32'd9775
; 
32'd186087: dataIn1 = 32'd9784
; 
32'd186088: dataIn1 = 32'd10209
; 
32'd186089: dataIn1 = 32'd10210
; 
32'd186090: dataIn1 = 32'd10240
; 
32'd186091: dataIn1 = 32'd10241
; 
32'd186092: dataIn1 = 32'd2720
; 
32'd186093: dataIn1 = 32'd6397
; 
32'd186094: dataIn1 = 32'd6712
; 
32'd186095: dataIn1 = 32'd6716
; 
32'd186096: dataIn1 = 32'd9748
; 
32'd186097: dataIn1 = 32'd9776
; 
32'd186098: dataIn1 = 32'd6119
; 
32'd186099: dataIn1 = 32'd6122
; 
32'd186100: dataIn1 = 32'd7171
; 
32'd186101: dataIn1 = 32'd9710
; 
32'd186102: dataIn1 = 32'd9759
; 
32'd186103: dataIn1 = 32'd9777
; 
32'd186104: dataIn1 = 32'd9785
; 
32'd186105: dataIn1 = 32'd5143
; 
32'd186106: dataIn1 = 32'd6161
; 
32'd186107: dataIn1 = 32'd7258
; 
32'd186108: dataIn1 = 32'd9767
; 
32'd186109: dataIn1 = 32'd9778
; 
32'd186110: dataIn1 = 32'd10124
; 
32'd186111: dataIn1 = 32'd10151
; 
32'd186112: dataIn1 = 32'd5887
; 
32'd186113: dataIn1 = 32'd6596
; 
32'd186114: dataIn1 = 32'd6598
; 
32'd186115: dataIn1 = 32'd7050
; 
32'd186116: dataIn1 = 32'd9768
; 
32'd186117: dataIn1 = 32'd9779
; 
32'd186118: dataIn1 = 32'd51
; 
32'd186119: dataIn1 = 32'd2174
; 
32'd186120: dataIn1 = 32'd2175
; 
32'd186121: dataIn1 = 32'd3631
; 
32'd186122: dataIn1 = 32'd9771
; 
32'd186123: dataIn1 = 32'd9780
; 
32'd186124: dataIn1 = 32'd41
; 
32'd186125: dataIn1 = 32'd2145
; 
32'd186126: dataIn1 = 32'd2175
; 
32'd186127: dataIn1 = 32'd9467
; 
32'd186128: dataIn1 = 32'd9770
; 
32'd186129: dataIn1 = 32'd9781
; 
32'd186130: dataIn1 = 32'd10227
; 
32'd186131: dataIn1 = 32'd56
; 
32'd186132: dataIn1 = 32'd2215
; 
32'd186133: dataIn1 = 32'd2218
; 
32'd186134: dataIn1 = 32'd5310
; 
32'd186135: dataIn1 = 32'd9773
; 
32'd186136: dataIn1 = 32'd9782
; 
32'd186137: dataIn1 = 32'd2189
; 
32'd186138: dataIn1 = 32'd2218
; 
32'd186139: dataIn1 = 32'd2219
; 
32'd186140: dataIn1 = 32'd9772
; 
32'd186141: dataIn1 = 32'd9774
; 
32'd186142: dataIn1 = 32'd9783
; 
32'd186143: dataIn1 = 32'd10239
; 
32'd186144: dataIn1 = 32'd57
; 
32'd186145: dataIn1 = 32'd2219
; 
32'd186146: dataIn1 = 32'd2221
; 
32'd186147: dataIn1 = 32'd3661
; 
32'd186148: dataIn1 = 32'd9775
; 
32'd186149: dataIn1 = 32'd9784
; 
32'd186150: dataIn1 = 32'd10241
; 
32'd186151: dataIn1 = 32'd6119
; 
32'd186152: dataIn1 = 32'd6123
; 
32'd186153: dataIn1 = 32'd7169
; 
32'd186154: dataIn1 = 32'd9710
; 
32'd186155: dataIn1 = 32'd9777
; 
32'd186156: dataIn1 = 32'd9785
; 
32'd186157: dataIn1 = 32'd9786
; 
32'd186158: dataIn1 = 32'd5127
; 
32'd186159: dataIn1 = 32'd6123
; 
32'd186160: dataIn1 = 32'd7169
; 
32'd186161: dataIn1 = 32'd9717
; 
32'd186162: dataIn1 = 32'd9785
; 
32'd186163: dataIn1 = 32'd9786
; 
32'd186164: dataIn1 = 32'd9787
; 
32'd186165: dataIn1 = 32'd5127
; 
32'd186166: dataIn1 = 32'd6133
; 
32'd186167: dataIn1 = 32'd7207
; 
32'd186168: dataIn1 = 32'd9717
; 
32'd186169: dataIn1 = 32'd9786
; 
32'd186170: dataIn1 = 32'd9787
; 
32'd186171: dataIn1 = 32'd9788
; 
32'd186172: dataIn1 = 32'd6133
; 
32'd186173: dataIn1 = 32'd6135
; 
32'd186174: dataIn1 = 32'd7207
; 
32'd186175: dataIn1 = 32'd9715
; 
32'd186176: dataIn1 = 32'd9787
; 
32'd186177: dataIn1 = 32'd9788
; 
32'd186178: dataIn1 = 32'd9789
; 
32'd186179: dataIn1 = 32'd6134
; 
32'd186180: dataIn1 = 32'd6135
; 
32'd186181: dataIn1 = 32'd7206
; 
32'd186182: dataIn1 = 32'd9715
; 
32'd186183: dataIn1 = 32'd9788
; 
32'd186184: dataIn1 = 32'd9789
; 
32'd186185: dataIn1 = 32'd9790
; 
32'd186186: dataIn1 = 32'd5117
; 
32'd186187: dataIn1 = 32'd6134
; 
32'd186188: dataIn1 = 32'd7206
; 
32'd186189: dataIn1 = 32'd9721
; 
32'd186190: dataIn1 = 32'd9789
; 
32'd186191: dataIn1 = 32'd9790
; 
32'd186192: dataIn1 = 32'd9791
; 
32'd186193: dataIn1 = 32'd5117
; 
32'd186194: dataIn1 = 32'd6088
; 
32'd186195: dataIn1 = 32'd7089
; 
32'd186196: dataIn1 = 32'd9721
; 
32'd186197: dataIn1 = 32'd9790
; 
32'd186198: dataIn1 = 32'd9791
; 
32'd186199: dataIn1 = 32'd9792
; 
32'd186200: dataIn1 = 32'd6084
; 
32'd186201: dataIn1 = 32'd6088
; 
32'd186202: dataIn1 = 32'd7089
; 
32'd186203: dataIn1 = 32'd9678
; 
32'd186204: dataIn1 = 32'd9791
; 
32'd186205: dataIn1 = 32'd9792
; 
32'd186206: dataIn1 = 32'd9793
; 
32'd186207: dataIn1 = 32'd6084
; 
32'd186208: dataIn1 = 32'd6087
; 
32'd186209: dataIn1 = 32'd7092
; 
32'd186210: dataIn1 = 32'd9678
; 
32'd186211: dataIn1 = 32'd9792
; 
32'd186212: dataIn1 = 32'd9793
; 
32'd186213: dataIn1 = 32'd9794
; 
32'd186214: dataIn1 = 32'd5118
; 
32'd186215: dataIn1 = 32'd6087
; 
32'd186216: dataIn1 = 32'd7092
; 
32'd186217: dataIn1 = 32'd9702
; 
32'd186218: dataIn1 = 32'd9793
; 
32'd186219: dataIn1 = 32'd9794
; 
32'd186220: dataIn1 = 32'd9795
; 
32'd186221: dataIn1 = 32'd5118
; 
32'd186222: dataIn1 = 32'd6112
; 
32'd186223: dataIn1 = 32'd7145
; 
32'd186224: dataIn1 = 32'd9702
; 
32'd186225: dataIn1 = 32'd9794
; 
32'd186226: dataIn1 = 32'd9795
; 
32'd186227: dataIn1 = 32'd9796
; 
32'd186228: dataIn1 = 32'd6111
; 
32'd186229: dataIn1 = 32'd6112
; 
32'd186230: dataIn1 = 32'd7145
; 
32'd186231: dataIn1 = 32'd9697
; 
32'd186232: dataIn1 = 32'd9795
; 
32'd186233: dataIn1 = 32'd9796
; 
32'd186234: dataIn1 = 32'd9797
; 
32'd186235: dataIn1 = 32'd6111
; 
32'd186236: dataIn1 = 32'd6113
; 
32'd186237: dataIn1 = 32'd7144
; 
32'd186238: dataIn1 = 32'd9697
; 
32'd186239: dataIn1 = 32'd9796
; 
32'd186240: dataIn1 = 32'd9797
; 
32'd186241: dataIn1 = 32'd9798
; 
32'd186242: dataIn1 = 32'd5122
; 
32'd186243: dataIn1 = 32'd6113
; 
32'd186244: dataIn1 = 32'd7144
; 
32'd186245: dataIn1 = 32'd9706
; 
32'd186246: dataIn1 = 32'd9797
; 
32'd186247: dataIn1 = 32'd9798
; 
32'd186248: dataIn1 = 32'd9799
; 
32'd186249: dataIn1 = 32'd5122
; 
32'd186250: dataIn1 = 32'd6104
; 
32'd186251: dataIn1 = 32'd7116
; 
32'd186252: dataIn1 = 32'd9706
; 
32'd186253: dataIn1 = 32'd9798
; 
32'd186254: dataIn1 = 32'd9799
; 
32'd186255: dataIn1 = 32'd9800
; 
32'd186256: dataIn1 = 32'd6099
; 
32'd186257: dataIn1 = 32'd6104
; 
32'd186258: dataIn1 = 32'd7116
; 
32'd186259: dataIn1 = 32'd9682
; 
32'd186260: dataIn1 = 32'd9799
; 
32'd186261: dataIn1 = 32'd9800
; 
32'd186262: dataIn1 = 32'd9801
; 
32'd186263: dataIn1 = 32'd6099
; 
32'd186264: dataIn1 = 32'd6105
; 
32'd186265: dataIn1 = 32'd7114
; 
32'd186266: dataIn1 = 32'd9682
; 
32'd186267: dataIn1 = 32'd9800
; 
32'd186268: dataIn1 = 32'd9801
; 
32'd186269: dataIn1 = 32'd9802
; 
32'd186270: dataIn1 = 32'd5121
; 
32'd186271: dataIn1 = 32'd6105
; 
32'd186272: dataIn1 = 32'd7114
; 
32'd186273: dataIn1 = 32'd9692
; 
32'd186274: dataIn1 = 32'd9801
; 
32'd186275: dataIn1 = 32'd9802
; 
32'd186276: dataIn1 = 32'd9803
; 
32'd186277: dataIn1 = 32'd5121
; 
32'd186278: dataIn1 = 32'd6108
; 
32'd186279: dataIn1 = 32'd7137
; 
32'd186280: dataIn1 = 32'd9692
; 
32'd186281: dataIn1 = 32'd9802
; 
32'd186282: dataIn1 = 32'd9803
; 
32'd186283: dataIn1 = 32'd9804
; 
32'd186284: dataIn1 = 32'd6107
; 
32'd186285: dataIn1 = 32'd6108
; 
32'd186286: dataIn1 = 32'd7137
; 
32'd186287: dataIn1 = 32'd9684
; 
32'd186288: dataIn1 = 32'd9803
; 
32'd186289: dataIn1 = 32'd9804
; 
32'd186290: dataIn1 = 32'd9805
; 
32'd186291: dataIn1 = 32'd6106
; 
32'd186292: dataIn1 = 32'd6107
; 
32'd186293: dataIn1 = 32'd7139
; 
32'd186294: dataIn1 = 32'd9684
; 
32'd186295: dataIn1 = 32'd9804
; 
32'd186296: dataIn1 = 32'd9805
; 
32'd186297: dataIn1 = 32'd9806
; 
32'd186298: dataIn1 = 32'd5124
; 
32'd186299: dataIn1 = 32'd6106
; 
32'd186300: dataIn1 = 32'd7139
; 
32'd186301: dataIn1 = 32'd9688
; 
32'd186302: dataIn1 = 32'd9805
; 
32'd186303: dataIn1 = 32'd9806
; 
32'd186304: dataIn1 = 32'd9807
; 
32'd186305: dataIn1 = 32'd5124
; 
32'd186306: dataIn1 = 32'd6109
; 
32'd186307: dataIn1 = 32'd9369
; 
32'd186308: dataIn1 = 32'd9688
; 
32'd186309: dataIn1 = 32'd9806
; 
32'd186310: dataIn1 = 32'd9807
; 
32'd186311: dataIn1 = 32'd9808
; 
32'd186312: dataIn1 = 32'd6109
; 
32'd186313: dataIn1 = 32'd6811
; 
32'd186314: dataIn1 = 32'd9369
; 
32'd186315: dataIn1 = 32'd9756
; 
32'd186316: dataIn1 = 32'd9807
; 
32'd186317: dataIn1 = 32'd9808
; 
32'd186318: dataIn1 = 32'd9809
; 
32'd186319: dataIn1 = 32'd6811
; 
32'd186320: dataIn1 = 32'd6814
; 
32'd186321: dataIn1 = 32'd9371
; 
32'd186322: dataIn1 = 32'd9756
; 
32'd186323: dataIn1 = 32'd9808
; 
32'd186324: dataIn1 = 32'd9809
; 
32'd186325: dataIn1 = 32'd9810
; 
32'd186326: dataIn1 = 32'd5638
; 
32'd186327: dataIn1 = 32'd6814
; 
32'd186328: dataIn1 = 32'd9371
; 
32'd186329: dataIn1 = 32'd9809
; 
32'd186330: dataIn1 = 32'd9810
; 
32'd186331: dataIn1 = 32'd2114
; 
32'd186332: dataIn1 = 32'd9451
; 
32'd186333: dataIn1 = 32'd9811
; 
32'd186334: dataIn1 = 32'd9812
; 
32'd186335: dataIn1 = 32'd9813
; 
32'd186336: dataIn1 = 32'd9817
; 
32'd186337: dataIn1 = 32'd9821
; 
32'd186338: dataIn1 = 32'd9449
; 
32'd186339: dataIn1 = 32'd9450
; 
32'd186340: dataIn1 = 32'd9451
; 
32'd186341: dataIn1 = 32'd9811
; 
32'd186342: dataIn1 = 32'd9812
; 
32'd186343: dataIn1 = 32'd9813
; 
32'd186344: dataIn1 = 32'd2114
; 
32'd186345: dataIn1 = 32'd9449
; 
32'd186346: dataIn1 = 32'd9811
; 
32'd186347: dataIn1 = 32'd9812
; 
32'd186348: dataIn1 = 32'd9813
; 
32'd186349: dataIn1 = 32'd9814
; 
32'd186350: dataIn1 = 32'd9815
; 
32'd186351: dataIn1 = 32'd2114
; 
32'd186352: dataIn1 = 32'd9453
; 
32'd186353: dataIn1 = 32'd9813
; 
32'd186354: dataIn1 = 32'd9814
; 
32'd186355: dataIn1 = 32'd9815
; 
32'd186356: dataIn1 = 32'd9824
; 
32'd186357: dataIn1 = 32'd9826
; 
32'd186358: dataIn1 = 32'd9449
; 
32'd186359: dataIn1 = 32'd9452
; 
32'd186360: dataIn1 = 32'd9453
; 
32'd186361: dataIn1 = 32'd9813
; 
32'd186362: dataIn1 = 32'd9814
; 
32'd186363: dataIn1 = 32'd9815
; 
32'd186364: dataIn1 = 32'd9451
; 
32'd186365: dataIn1 = 32'd9455
; 
32'd186366: dataIn1 = 32'd9816
; 
32'd186367: dataIn1 = 32'd9817
; 
32'd186368: dataIn1 = 32'd9818
; 
32'd186369: dataIn1 = 32'd9819
; 
32'd186370: dataIn1 = 32'd9820
; 
32'd186371: dataIn1 = 32'd9451
; 
32'd186372: dataIn1 = 32'd9454
; 
32'd186373: dataIn1 = 32'd9811
; 
32'd186374: dataIn1 = 32'd9816
; 
32'd186375: dataIn1 = 32'd9817
; 
32'd186376: dataIn1 = 32'd9818
; 
32'd186377: dataIn1 = 32'd9821
; 
32'd186378: dataIn1 = 32'd31
; 
32'd186379: dataIn1 = 32'd9454
; 
32'd186380: dataIn1 = 32'd9455
; 
32'd186381: dataIn1 = 32'd9816
; 
32'd186382: dataIn1 = 32'd9817
; 
32'd186383: dataIn1 = 32'd9818
; 
32'd186384: dataIn1 = 32'd2113
; 
32'd186385: dataIn1 = 32'd9450
; 
32'd186386: dataIn1 = 32'd9451
; 
32'd186387: dataIn1 = 32'd9816
; 
32'd186388: dataIn1 = 32'd9819
; 
32'd186389: dataIn1 = 32'd9820
; 
32'd186390: dataIn1 = 32'd2113
; 
32'd186391: dataIn1 = 32'd9455
; 
32'd186392: dataIn1 = 32'd9816
; 
32'd186393: dataIn1 = 32'd9819
; 
32'd186394: dataIn1 = 32'd9820
; 
32'd186395: dataIn1 = 32'd9828
; 
32'd186396: dataIn1 = 32'd9832
; 
32'd186397: dataIn1 = 32'd2114
; 
32'd186398: dataIn1 = 32'd9454
; 
32'd186399: dataIn1 = 32'd9811
; 
32'd186400: dataIn1 = 32'd9817
; 
32'd186401: dataIn1 = 32'd9821
; 
32'd186402: dataIn1 = 32'd10152
; 
32'd186403: dataIn1 = 32'd5520
; 
32'd186404: dataIn1 = 32'd9453
; 
32'd186405: dataIn1 = 32'd9674
; 
32'd186406: dataIn1 = 32'd9822
; 
32'd186407: dataIn1 = 32'd9823
; 
32'd186408: dataIn1 = 32'd9824
; 
32'd186409: dataIn1 = 32'd9825
; 
32'd186410: dataIn1 = 32'd10133
; 
32'd186411: dataIn1 = 32'd5520
; 
32'd186412: dataIn1 = 32'd9456
; 
32'd186413: dataIn1 = 32'd9822
; 
32'd186414: dataIn1 = 32'd9823
; 
32'd186415: dataIn1 = 32'd9824
; 
32'd186416: dataIn1 = 32'd10276
; 
32'd186417: dataIn1 = 32'd10283
; 
32'd186418: dataIn1 = 32'd9453
; 
32'd186419: dataIn1 = 32'd9456
; 
32'd186420: dataIn1 = 32'd9814
; 
32'd186421: dataIn1 = 32'd9822
; 
32'd186422: dataIn1 = 32'd9823
; 
32'd186423: dataIn1 = 32'd9824
; 
32'd186424: dataIn1 = 32'd9826
; 
32'd186425: dataIn1 = 32'd20
; 
32'd186426: dataIn1 = 32'd9452
; 
32'd186427: dataIn1 = 32'd9453
; 
32'd186428: dataIn1 = 32'd9674
; 
32'd186429: dataIn1 = 32'd9822
; 
32'd186430: dataIn1 = 32'd9825
; 
32'd186431: dataIn1 = 32'd2114
; 
32'd186432: dataIn1 = 32'd9456
; 
32'd186433: dataIn1 = 32'd9814
; 
32'd186434: dataIn1 = 32'd9824
; 
32'd186435: dataIn1 = 32'd9826
; 
32'd186436: dataIn1 = 32'd10152
; 
32'd186437: dataIn1 = 32'd9457
; 
32'd186438: dataIn1 = 32'd9458
; 
32'd186439: dataIn1 = 32'd9827
; 
32'd186440: dataIn1 = 32'd9828
; 
32'd186441: dataIn1 = 32'd9829
; 
32'd186442: dataIn1 = 32'd9830
; 
32'd186443: dataIn1 = 32'd9831
; 
32'd186444: dataIn1 = 32'd9455
; 
32'd186445: dataIn1 = 32'd9458
; 
32'd186446: dataIn1 = 32'd9820
; 
32'd186447: dataIn1 = 32'd9827
; 
32'd186448: dataIn1 = 32'd9828
; 
32'd186449: dataIn1 = 32'd9829
; 
32'd186450: dataIn1 = 32'd9832
; 
32'd186451: dataIn1 = 32'd31
; 
32'd186452: dataIn1 = 32'd9455
; 
32'd186453: dataIn1 = 32'd9457
; 
32'd186454: dataIn1 = 32'd9827
; 
32'd186455: dataIn1 = 32'd9828
; 
32'd186456: dataIn1 = 32'd9829
; 
32'd186457: dataIn1 = 32'd2147
; 
32'd186458: dataIn1 = 32'd9458
; 
32'd186459: dataIn1 = 32'd9827
; 
32'd186460: dataIn1 = 32'd9830
; 
32'd186461: dataIn1 = 32'd9831
; 
32'd186462: dataIn1 = 32'd10156
; 
32'd186463: dataIn1 = 32'd2147
; 
32'd186464: dataIn1 = 32'd9457
; 
32'd186465: dataIn1 = 32'd9827
; 
32'd186466: dataIn1 = 32'd9830
; 
32'd186467: dataIn1 = 32'd9831
; 
32'd186468: dataIn1 = 32'd9834
; 
32'd186469: dataIn1 = 32'd9836
; 
32'd186470: dataIn1 = 32'd2113
; 
32'd186471: dataIn1 = 32'd9458
; 
32'd186472: dataIn1 = 32'd9820
; 
32'd186473: dataIn1 = 32'd9828
; 
32'd186474: dataIn1 = 32'd9832
; 
32'd186475: dataIn1 = 32'd10155
; 
32'd186476: dataIn1 = 32'd2147
; 
32'd186477: dataIn1 = 32'd9460
; 
32'd186478: dataIn1 = 32'd9833
; 
32'd186479: dataIn1 = 32'd9834
; 
32'd186480: dataIn1 = 32'd9835
; 
32'd186481: dataIn1 = 32'd9839
; 
32'd186482: dataIn1 = 32'd9842
; 
32'd186483: dataIn1 = 32'd2147
; 
32'd186484: dataIn1 = 32'd9459
; 
32'd186485: dataIn1 = 32'd9831
; 
32'd186486: dataIn1 = 32'd9833
; 
32'd186487: dataIn1 = 32'd9834
; 
32'd186488: dataIn1 = 32'd9835
; 
32'd186489: dataIn1 = 32'd9836
; 
32'd186490: dataIn1 = 32'd9459
; 
32'd186491: dataIn1 = 32'd9460
; 
32'd186492: dataIn1 = 32'd9461
; 
32'd186493: dataIn1 = 32'd9833
; 
32'd186494: dataIn1 = 32'd9834
; 
32'd186495: dataIn1 = 32'd9835
; 
32'd186496: dataIn1 = 32'd9457
; 
32'd186497: dataIn1 = 32'd9459
; 
32'd186498: dataIn1 = 32'd9462
; 
32'd186499: dataIn1 = 32'd9831
; 
32'd186500: dataIn1 = 32'd9834
; 
32'd186501: dataIn1 = 32'd9836
; 
32'd186502: dataIn1 = 32'd9460
; 
32'd186503: dataIn1 = 32'd9464
; 
32'd186504: dataIn1 = 32'd9837
; 
32'd186505: dataIn1 = 32'd9838
; 
32'd186506: dataIn1 = 32'd9839
; 
32'd186507: dataIn1 = 32'd9840
; 
32'd186508: dataIn1 = 32'd9841
; 
32'd186509: dataIn1 = 32'd41
; 
32'd186510: dataIn1 = 32'd9463
; 
32'd186511: dataIn1 = 32'd9464
; 
32'd186512: dataIn1 = 32'd9837
; 
32'd186513: dataIn1 = 32'd9838
; 
32'd186514: dataIn1 = 32'd9839
; 
32'd186515: dataIn1 = 32'd9460
; 
32'd186516: dataIn1 = 32'd9463
; 
32'd186517: dataIn1 = 32'd9833
; 
32'd186518: dataIn1 = 32'd9837
; 
32'd186519: dataIn1 = 32'd9838
; 
32'd186520: dataIn1 = 32'd9839
; 
32'd186521: dataIn1 = 32'd9842
; 
32'd186522: dataIn1 = 32'd2148
; 
32'd186523: dataIn1 = 32'd9464
; 
32'd186524: dataIn1 = 32'd9837
; 
32'd186525: dataIn1 = 32'd9840
; 
32'd186526: dataIn1 = 32'd9841
; 
32'd186527: dataIn1 = 32'd9846
; 
32'd186528: dataIn1 = 32'd9848
; 
32'd186529: dataIn1 = 32'd2148
; 
32'd186530: dataIn1 = 32'd9460
; 
32'd186531: dataIn1 = 32'd9461
; 
32'd186532: dataIn1 = 32'd9837
; 
32'd186533: dataIn1 = 32'd9840
; 
32'd186534: dataIn1 = 32'd9841
; 
32'd186535: dataIn1 = 32'd2147
; 
32'd186536: dataIn1 = 32'd9463
; 
32'd186537: dataIn1 = 32'd9833
; 
32'd186538: dataIn1 = 32'd9839
; 
32'd186539: dataIn1 = 32'd9842
; 
32'd186540: dataIn1 = 32'd10156
; 
32'd186541: dataIn1 = 32'd2177
; 
32'd186542: dataIn1 = 32'd9465
; 
32'd186543: dataIn1 = 32'd9475
; 
32'd186544: dataIn1 = 32'd9843
; 
32'd186545: dataIn1 = 32'd9844
; 
32'd186546: dataIn1 = 32'd9847
; 
32'd186547: dataIn1 = 32'd9849
; 
32'd186548: dataIn1 = 32'd9865
; 
32'd186549: dataIn1 = 32'd3590
; 
32'd186550: dataIn1 = 32'd9465
; 
32'd186551: dataIn1 = 32'd9466
; 
32'd186552: dataIn1 = 32'd9475
; 
32'd186553: dataIn1 = 32'd9843
; 
32'd186554: dataIn1 = 32'd9844
; 
32'd186555: dataIn1 = 32'd41
; 
32'd186556: dataIn1 = 32'd9464
; 
32'd186557: dataIn1 = 32'd9467
; 
32'd186558: dataIn1 = 32'd9845
; 
32'd186559: dataIn1 = 32'd9846
; 
32'd186560: dataIn1 = 32'd9847
; 
32'd186561: dataIn1 = 32'd9464
; 
32'd186562: dataIn1 = 32'd9465
; 
32'd186563: dataIn1 = 32'd9840
; 
32'd186564: dataIn1 = 32'd9845
; 
32'd186565: dataIn1 = 32'd9846
; 
32'd186566: dataIn1 = 32'd9847
; 
32'd186567: dataIn1 = 32'd9848
; 
32'd186568: dataIn1 = 32'd9465
; 
32'd186569: dataIn1 = 32'd9467
; 
32'd186570: dataIn1 = 32'd9843
; 
32'd186571: dataIn1 = 32'd9845
; 
32'd186572: dataIn1 = 32'd9846
; 
32'd186573: dataIn1 = 32'd9847
; 
32'd186574: dataIn1 = 32'd9849
; 
32'd186575: dataIn1 = 32'd2148
; 
32'd186576: dataIn1 = 32'd9465
; 
32'd186577: dataIn1 = 32'd9466
; 
32'd186578: dataIn1 = 32'd9840
; 
32'd186579: dataIn1 = 32'd9846
; 
32'd186580: dataIn1 = 32'd9848
; 
32'd186581: dataIn1 = 32'd2177
; 
32'd186582: dataIn1 = 32'd9467
; 
32'd186583: dataIn1 = 32'd9843
; 
32'd186584: dataIn1 = 32'd9847
; 
32'd186585: dataIn1 = 32'd9849
; 
32'd186586: dataIn1 = 32'd10161
; 
32'd186587: dataIn1 = 32'd10227
; 
32'd186588: dataIn1 = 32'd3587
; 
32'd186589: dataIn1 = 32'd9469
; 
32'd186590: dataIn1 = 32'd9470
; 
32'd186591: dataIn1 = 32'd9850
; 
32'd186592: dataIn1 = 32'd9851
; 
32'd186593: dataIn1 = 32'd9852
; 
32'd186594: dataIn1 = 32'd9468
; 
32'd186595: dataIn1 = 32'd9470
; 
32'd186596: dataIn1 = 32'd9850
; 
32'd186597: dataIn1 = 32'd9851
; 
32'd186598: dataIn1 = 32'd9852
; 
32'd186599: dataIn1 = 32'd9853
; 
32'd186600: dataIn1 = 32'd9854
; 
32'd186601: dataIn1 = 32'd9468
; 
32'd186602: dataIn1 = 32'd9469
; 
32'd186603: dataIn1 = 32'd9850
; 
32'd186604: dataIn1 = 32'd9851
; 
32'd186605: dataIn1 = 32'd9852
; 
32'd186606: dataIn1 = 32'd9855
; 
32'd186607: dataIn1 = 32'd9856
; 
32'd186608: dataIn1 = 32'd3588
; 
32'd186609: dataIn1 = 32'd9470
; 
32'd186610: dataIn1 = 32'd9851
; 
32'd186611: dataIn1 = 32'd9853
; 
32'd186612: dataIn1 = 32'd9854
; 
32'd186613: dataIn1 = 32'd10158
; 
32'd186614: dataIn1 = 32'd3588
; 
32'd186615: dataIn1 = 32'd9468
; 
32'd186616: dataIn1 = 32'd9851
; 
32'd186617: dataIn1 = 32'd9853
; 
32'd186618: dataIn1 = 32'd9854
; 
32'd186619: dataIn1 = 32'd9857
; 
32'd186620: dataIn1 = 32'd9858
; 
32'd186621: dataIn1 = 32'd3589
; 
32'd186622: dataIn1 = 32'd9469
; 
32'd186623: dataIn1 = 32'd9852
; 
32'd186624: dataIn1 = 32'd9855
; 
32'd186625: dataIn1 = 32'd9856
; 
32'd186626: dataIn1 = 32'd9861
; 
32'd186627: dataIn1 = 32'd9864
; 
32'd186628: dataIn1 = 32'd3589
; 
32'd186629: dataIn1 = 32'd9468
; 
32'd186630: dataIn1 = 32'd9471
; 
32'd186631: dataIn1 = 32'd9852
; 
32'd186632: dataIn1 = 32'd9855
; 
32'd186633: dataIn1 = 32'd9856
; 
32'd186634: dataIn1 = 32'd3588
; 
32'd186635: dataIn1 = 32'd9472
; 
32'd186636: dataIn1 = 32'd9854
; 
32'd186637: dataIn1 = 32'd9857
; 
32'd186638: dataIn1 = 32'd9858
; 
32'd186639: dataIn1 = 32'd9906
; 
32'd186640: dataIn1 = 32'd9909
; 
32'd186641: dataIn1 = 32'd9468
; 
32'd186642: dataIn1 = 32'd9471
; 
32'd186643: dataIn1 = 32'd9472
; 
32'd186644: dataIn1 = 32'd9854
; 
32'd186645: dataIn1 = 32'd9857
; 
32'd186646: dataIn1 = 32'd9858
; 
32'd186647: dataIn1 = 32'd3587
; 
32'd186648: dataIn1 = 32'd9469
; 
32'd186649: dataIn1 = 32'd9474
; 
32'd186650: dataIn1 = 32'd9859
; 
32'd186651: dataIn1 = 32'd9860
; 
32'd186652: dataIn1 = 32'd9861
; 
32'd186653: dataIn1 = 32'd9473
; 
32'd186654: dataIn1 = 32'd9474
; 
32'd186655: dataIn1 = 32'd9859
; 
32'd186656: dataIn1 = 32'd9860
; 
32'd186657: dataIn1 = 32'd9861
; 
32'd186658: dataIn1 = 32'd9862
; 
32'd186659: dataIn1 = 32'd9863
; 
32'd186660: dataIn1 = 32'd9469
; 
32'd186661: dataIn1 = 32'd9473
; 
32'd186662: dataIn1 = 32'd9855
; 
32'd186663: dataIn1 = 32'd9859
; 
32'd186664: dataIn1 = 32'd9860
; 
32'd186665: dataIn1 = 32'd9861
; 
32'd186666: dataIn1 = 32'd9864
; 
32'd186667: dataIn1 = 32'd2177
; 
32'd186668: dataIn1 = 32'd9474
; 
32'd186669: dataIn1 = 32'd9860
; 
32'd186670: dataIn1 = 32'd9862
; 
32'd186671: dataIn1 = 32'd9863
; 
32'd186672: dataIn1 = 32'd9865
; 
32'd186673: dataIn1 = 32'd9866
; 
32'd186674: dataIn1 = 32'd2177
; 
32'd186675: dataIn1 = 32'd9473
; 
32'd186676: dataIn1 = 32'd9860
; 
32'd186677: dataIn1 = 32'd9862
; 
32'd186678: dataIn1 = 32'd9863
; 
32'd186679: dataIn1 = 32'd10161
; 
32'd186680: dataIn1 = 32'd3589
; 
32'd186681: dataIn1 = 32'd9473
; 
32'd186682: dataIn1 = 32'd9855
; 
32'd186683: dataIn1 = 32'd9861
; 
32'd186684: dataIn1 = 32'd9864
; 
32'd186685: dataIn1 = 32'd10160
; 
32'd186686: dataIn1 = 32'd2177
; 
32'd186687: dataIn1 = 32'd9475
; 
32'd186688: dataIn1 = 32'd9843
; 
32'd186689: dataIn1 = 32'd9862
; 
32'd186690: dataIn1 = 32'd9865
; 
32'd186691: dataIn1 = 32'd9866
; 
32'd186692: dataIn1 = 32'd9474
; 
32'd186693: dataIn1 = 32'd9475
; 
32'd186694: dataIn1 = 32'd9476
; 
32'd186695: dataIn1 = 32'd9862
; 
32'd186696: dataIn1 = 32'd9865
; 
32'd186697: dataIn1 = 32'd9866
; 
32'd186698: dataIn1 = 32'd3622
; 
32'd186699: dataIn1 = 32'd9479
; 
32'd186700: dataIn1 = 32'd9867
; 
32'd186701: dataIn1 = 32'd9868
; 
32'd186702: dataIn1 = 32'd9869
; 
32'd186703: dataIn1 = 32'd9876
; 
32'd186704: dataIn1 = 32'd9877
; 
32'd186705: dataIn1 = 32'd3622
; 
32'd186706: dataIn1 = 32'd9478
; 
32'd186707: dataIn1 = 32'd9867
; 
32'd186708: dataIn1 = 32'd9868
; 
32'd186709: dataIn1 = 32'd9869
; 
32'd186710: dataIn1 = 32'd9872
; 
32'd186711: dataIn1 = 32'd9875
; 
32'd186712: dataIn1 = 32'd9478
; 
32'd186713: dataIn1 = 32'd9479
; 
32'd186714: dataIn1 = 32'd9480
; 
32'd186715: dataIn1 = 32'd9867
; 
32'd186716: dataIn1 = 32'd9868
; 
32'd186717: dataIn1 = 32'd9869
; 
32'd186718: dataIn1 = 32'd2204
; 
32'd186719: dataIn1 = 32'd9481
; 
32'd186720: dataIn1 = 32'd9482
; 
32'd186721: dataIn1 = 32'd9870
; 
32'd186722: dataIn1 = 32'd9871
; 
32'd186723: dataIn1 = 32'd9872
; 
32'd186724: dataIn1 = 32'd9478
; 
32'd186725: dataIn1 = 32'd9482
; 
32'd186726: dataIn1 = 32'd9870
; 
32'd186727: dataIn1 = 32'd9871
; 
32'd186728: dataIn1 = 32'd9872
; 
32'd186729: dataIn1 = 32'd9873
; 
32'd186730: dataIn1 = 32'd9874
; 
32'd186731: dataIn1 = 32'd9478
; 
32'd186732: dataIn1 = 32'd9481
; 
32'd186733: dataIn1 = 32'd9868
; 
32'd186734: dataIn1 = 32'd9870
; 
32'd186735: dataIn1 = 32'd9871
; 
32'd186736: dataIn1 = 32'd9872
; 
32'd186737: dataIn1 = 32'd9875
; 
32'd186738: dataIn1 = 32'd3621
; 
32'd186739: dataIn1 = 32'd9482
; 
32'd186740: dataIn1 = 32'd9871
; 
32'd186741: dataIn1 = 32'd9873
; 
32'd186742: dataIn1 = 32'd9874
; 
32'd186743: dataIn1 = 32'd9879
; 
32'd186744: dataIn1 = 32'd9881
; 
32'd186745: dataIn1 = 32'd3621
; 
32'd186746: dataIn1 = 32'd9478
; 
32'd186747: dataIn1 = 32'd9480
; 
32'd186748: dataIn1 = 32'd9871
; 
32'd186749: dataIn1 = 32'd9873
; 
32'd186750: dataIn1 = 32'd9874
; 
32'd186751: dataIn1 = 32'd3622
; 
32'd186752: dataIn1 = 32'd9481
; 
32'd186753: dataIn1 = 32'd9868
; 
32'd186754: dataIn1 = 32'd9872
; 
32'd186755: dataIn1 = 32'd9875
; 
32'd186756: dataIn1 = 32'd10162
; 
32'd186757: dataIn1 = 32'd3622
; 
32'd186758: dataIn1 = 32'd9483
; 
32'd186759: dataIn1 = 32'd9867
; 
32'd186760: dataIn1 = 32'd9876
; 
32'd186761: dataIn1 = 32'd9877
; 
32'd186762: dataIn1 = 32'd9886
; 
32'd186763: dataIn1 = 32'd9889
; 
32'd186764: dataIn1 = 32'd9479
; 
32'd186765: dataIn1 = 32'd9483
; 
32'd186766: dataIn1 = 32'd9484
; 
32'd186767: dataIn1 = 32'd9867
; 
32'd186768: dataIn1 = 32'd9876
; 
32'd186769: dataIn1 = 32'd9877
; 
32'd186770: dataIn1 = 32'd2204
; 
32'd186771: dataIn1 = 32'd9482
; 
32'd186772: dataIn1 = 32'd9486
; 
32'd186773: dataIn1 = 32'd9878
; 
32'd186774: dataIn1 = 32'd9879
; 
32'd186775: dataIn1 = 32'd9880
; 
32'd186776: dataIn1 = 32'd9482
; 
32'd186777: dataIn1 = 32'd9485
; 
32'd186778: dataIn1 = 32'd9873
; 
32'd186779: dataIn1 = 32'd9878
; 
32'd186780: dataIn1 = 32'd9879
; 
32'd186781: dataIn1 = 32'd9880
; 
32'd186782: dataIn1 = 32'd9881
; 
32'd186783: dataIn1 = 32'd9485
; 
32'd186784: dataIn1 = 32'd9486
; 
32'd186785: dataIn1 = 32'd9878
; 
32'd186786: dataIn1 = 32'd9879
; 
32'd186787: dataIn1 = 32'd9880
; 
32'd186788: dataIn1 = 32'd9882
; 
32'd186789: dataIn1 = 32'd9883
; 
32'd186790: dataIn1 = 32'd3621
; 
32'd186791: dataIn1 = 32'd9485
; 
32'd186792: dataIn1 = 32'd9873
; 
32'd186793: dataIn1 = 32'd9879
; 
32'd186794: dataIn1 = 32'd9881
; 
32'd186795: dataIn1 = 32'd10165
; 
32'd186796: dataIn1 = 32'd3625
; 
32'd186797: dataIn1 = 32'd9486
; 
32'd186798: dataIn1 = 32'd9880
; 
32'd186799: dataIn1 = 32'd9882
; 
32'd186800: dataIn1 = 32'd9883
; 
32'd186801: dataIn1 = 32'd10018
; 
32'd186802: dataIn1 = 32'd10026
; 
32'd186803: dataIn1 = 32'd3625
; 
32'd186804: dataIn1 = 32'd9485
; 
32'd186805: dataIn1 = 32'd9880
; 
32'd186806: dataIn1 = 32'd9882
; 
32'd186807: dataIn1 = 32'd9883
; 
32'd186808: dataIn1 = 32'd10164
; 
32'd186809: dataIn1 = 32'd3626
; 
32'd186810: dataIn1 = 32'd9487
; 
32'd186811: dataIn1 = 32'd9488
; 
32'd186812: dataIn1 = 32'd9884
; 
32'd186813: dataIn1 = 32'd9885
; 
32'd186814: dataIn1 = 32'd9886
; 
32'd186815: dataIn1 = 32'd9483
; 
32'd186816: dataIn1 = 32'd9488
; 
32'd186817: dataIn1 = 32'd9884
; 
32'd186818: dataIn1 = 32'd9885
; 
32'd186819: dataIn1 = 32'd9886
; 
32'd186820: dataIn1 = 32'd9887
; 
32'd186821: dataIn1 = 32'd9888
; 
32'd186822: dataIn1 = 32'd9483
; 
32'd186823: dataIn1 = 32'd9487
; 
32'd186824: dataIn1 = 32'd9876
; 
32'd186825: dataIn1 = 32'd9884
; 
32'd186826: dataIn1 = 32'd9885
; 
32'd186827: dataIn1 = 32'd9886
; 
32'd186828: dataIn1 = 32'd9889
; 
32'd186829: dataIn1 = 32'd2205
; 
32'd186830: dataIn1 = 32'd9488
; 
32'd186831: dataIn1 = 32'd9885
; 
32'd186832: dataIn1 = 32'd9887
; 
32'd186833: dataIn1 = 32'd9888
; 
32'd186834: dataIn1 = 32'd9904
; 
32'd186835: dataIn1 = 32'd9905
; 
32'd186836: dataIn1 = 32'd2205
; 
32'd186837: dataIn1 = 32'd9483
; 
32'd186838: dataIn1 = 32'd9484
; 
32'd186839: dataIn1 = 32'd9885
; 
32'd186840: dataIn1 = 32'd9887
; 
32'd186841: dataIn1 = 32'd9888
; 
32'd186842: dataIn1 = 32'd3622
; 
32'd186843: dataIn1 = 32'd9487
; 
32'd186844: dataIn1 = 32'd9876
; 
32'd186845: dataIn1 = 32'd9886
; 
32'd186846: dataIn1 = 32'd9889
; 
32'd186847: dataIn1 = 32'd10162
; 
32'd186848: dataIn1 = 32'd9490
; 
32'd186849: dataIn1 = 32'd9491
; 
32'd186850: dataIn1 = 32'd9890
; 
32'd186851: dataIn1 = 32'd9891
; 
32'd186852: dataIn1 = 32'd9892
; 
32'd186853: dataIn1 = 32'd9893
; 
32'd186854: dataIn1 = 32'd9894
; 
32'd186855: dataIn1 = 32'd3629
; 
32'd186856: dataIn1 = 32'd9489
; 
32'd186857: dataIn1 = 32'd9491
; 
32'd186858: dataIn1 = 32'd9890
; 
32'd186859: dataIn1 = 32'd9891
; 
32'd186860: dataIn1 = 32'd9892
; 
32'd186861: dataIn1 = 32'd9489
; 
32'd186862: dataIn1 = 32'd9490
; 
32'd186863: dataIn1 = 32'd9890
; 
32'd186864: dataIn1 = 32'd9891
; 
32'd186865: dataIn1 = 32'd9892
; 
32'd186866: dataIn1 = 32'd9895
; 
32'd186867: dataIn1 = 32'd9896
; 
32'd186868: dataIn1 = 32'd3628
; 
32'd186869: dataIn1 = 32'd9491
; 
32'd186870: dataIn1 = 32'd9890
; 
32'd186871: dataIn1 = 32'd9893
; 
32'd186872: dataIn1 = 32'd9894
; 
32'd186873: dataIn1 = 32'd9899
; 
32'd186874: dataIn1 = 32'd9902
; 
32'd186875: dataIn1 = 32'd3628
; 
32'd186876: dataIn1 = 32'd9490
; 
32'd186877: dataIn1 = 32'd9493
; 
32'd186878: dataIn1 = 32'd9890
; 
32'd186879: dataIn1 = 32'd9893
; 
32'd186880: dataIn1 = 32'd9894
; 
32'd186881: dataIn1 = 32'd3630
; 
32'd186882: dataIn1 = 32'd9490
; 
32'd186883: dataIn1 = 32'd9892
; 
32'd186884: dataIn1 = 32'd9895
; 
32'd186885: dataIn1 = 32'd9896
; 
32'd186886: dataIn1 = 32'd9897
; 
32'd186887: dataIn1 = 32'd9898
; 
32'd186888: dataIn1 = 32'd3630
; 
32'd186889: dataIn1 = 32'd9489
; 
32'd186890: dataIn1 = 32'd9892
; 
32'd186891: dataIn1 = 32'd9895
; 
32'd186892: dataIn1 = 32'd9896
; 
32'd186893: dataIn1 = 32'd10167
; 
32'd186894: dataIn1 = 32'd3630
; 
32'd186895: dataIn1 = 32'd9492
; 
32'd186896: dataIn1 = 32'd9895
; 
32'd186897: dataIn1 = 32'd9897
; 
32'd186898: dataIn1 = 32'd9898
; 
32'd186899: dataIn1 = 32'd9908
; 
32'd186900: dataIn1 = 32'd9910
; 
32'd186901: dataIn1 = 32'd9490
; 
32'd186902: dataIn1 = 32'd9492
; 
32'd186903: dataIn1 = 32'd9493
; 
32'd186904: dataIn1 = 32'd9895
; 
32'd186905: dataIn1 = 32'd9897
; 
32'd186906: dataIn1 = 32'd9898
; 
32'd186907: dataIn1 = 32'd9491
; 
32'd186908: dataIn1 = 32'd9495
; 
32'd186909: dataIn1 = 32'd9893
; 
32'd186910: dataIn1 = 32'd9899
; 
32'd186911: dataIn1 = 32'd9900
; 
32'd186912: dataIn1 = 32'd9901
; 
32'd186913: dataIn1 = 32'd9902
; 
32'd186914: dataIn1 = 32'd3629
; 
32'd186915: dataIn1 = 32'd9491
; 
32'd186916: dataIn1 = 32'd9494
; 
32'd186917: dataIn1 = 32'd9899
; 
32'd186918: dataIn1 = 32'd9900
; 
32'd186919: dataIn1 = 32'd9901
; 
32'd186920: dataIn1 = 32'd9494
; 
32'd186921: dataIn1 = 32'd9495
; 
32'd186922: dataIn1 = 32'd9899
; 
32'd186923: dataIn1 = 32'd9900
; 
32'd186924: dataIn1 = 32'd9901
; 
32'd186925: dataIn1 = 32'd9903
; 
32'd186926: dataIn1 = 32'd9904
; 
32'd186927: dataIn1 = 32'd3628
; 
32'd186928: dataIn1 = 32'd9495
; 
32'd186929: dataIn1 = 32'd9893
; 
32'd186930: dataIn1 = 32'd9899
; 
32'd186931: dataIn1 = 32'd9902
; 
32'd186932: dataIn1 = 32'd10170
; 
32'd186933: dataIn1 = 32'd2205
; 
32'd186934: dataIn1 = 32'd9495
; 
32'd186935: dataIn1 = 32'd9901
; 
32'd186936: dataIn1 = 32'd9903
; 
32'd186937: dataIn1 = 32'd9904
; 
32'd186938: dataIn1 = 32'd10169
; 
32'd186939: dataIn1 = 32'd2205
; 
32'd186940: dataIn1 = 32'd9494
; 
32'd186941: dataIn1 = 32'd9887
; 
32'd186942: dataIn1 = 32'd9901
; 
32'd186943: dataIn1 = 32'd9903
; 
32'd186944: dataIn1 = 32'd9904
; 
32'd186945: dataIn1 = 32'd9905
; 
32'd186946: dataIn1 = 32'd9488
; 
32'd186947: dataIn1 = 32'd9494
; 
32'd186948: dataIn1 = 32'd9496
; 
32'd186949: dataIn1 = 32'd9887
; 
32'd186950: dataIn1 = 32'd9904
; 
32'd186951: dataIn1 = 32'd9905
; 
32'd186952: dataIn1 = 32'd9472
; 
32'd186953: dataIn1 = 32'd9497
; 
32'd186954: dataIn1 = 32'd9857
; 
32'd186955: dataIn1 = 32'd9906
; 
32'd186956: dataIn1 = 32'd9907
; 
32'd186957: dataIn1 = 32'd9908
; 
32'd186958: dataIn1 = 32'd9909
; 
32'd186959: dataIn1 = 32'd2176
; 
32'd186960: dataIn1 = 32'd9472
; 
32'd186961: dataIn1 = 32'd9492
; 
32'd186962: dataIn1 = 32'd9906
; 
32'd186963: dataIn1 = 32'd9907
; 
32'd186964: dataIn1 = 32'd9908
; 
32'd186965: dataIn1 = 32'd9492
; 
32'd186966: dataIn1 = 32'd9497
; 
32'd186967: dataIn1 = 32'd9897
; 
32'd186968: dataIn1 = 32'd9906
; 
32'd186969: dataIn1 = 32'd9907
; 
32'd186970: dataIn1 = 32'd9908
; 
32'd186971: dataIn1 = 32'd9910
; 
32'd186972: dataIn1 = 32'd3588
; 
32'd186973: dataIn1 = 32'd9497
; 
32'd186974: dataIn1 = 32'd9857
; 
32'd186975: dataIn1 = 32'd9906
; 
32'd186976: dataIn1 = 32'd9909
; 
32'd186977: dataIn1 = 32'd10172
; 
32'd186978: dataIn1 = 32'd3630
; 
32'd186979: dataIn1 = 32'd9497
; 
32'd186980: dataIn1 = 32'd9897
; 
32'd186981: dataIn1 = 32'd9908
; 
32'd186982: dataIn1 = 32'd9910
; 
32'd186983: dataIn1 = 32'd10171
; 
32'd186984: dataIn1 = 32'd3669
; 
32'd186985: dataIn1 = 32'd9500
; 
32'd186986: dataIn1 = 32'd9911
; 
32'd186987: dataIn1 = 32'd9912
; 
32'd186988: dataIn1 = 32'd9913
; 
32'd186989: dataIn1 = 32'd9917
; 
32'd186990: dataIn1 = 32'd9919
; 
32'd186991: dataIn1 = 32'd9498
; 
32'd186992: dataIn1 = 32'd9499
; 
32'd186993: dataIn1 = 32'd9500
; 
32'd186994: dataIn1 = 32'd9911
; 
32'd186995: dataIn1 = 32'd9912
; 
32'd186996: dataIn1 = 32'd9913
; 
32'd186997: dataIn1 = 32'd3669
; 
32'd186998: dataIn1 = 32'd9498
; 
32'd186999: dataIn1 = 32'd9911
; 
32'd187000: dataIn1 = 32'd9912
; 
32'd187001: dataIn1 = 32'd9913
; 
32'd187002: dataIn1 = 32'd9914
; 
32'd187003: dataIn1 = 32'd9915
; 
32'd187004: dataIn1 = 32'd3669
; 
32'd187005: dataIn1 = 32'd9502
; 
32'd187006: dataIn1 = 32'd9913
; 
32'd187007: dataIn1 = 32'd9914
; 
32'd187008: dataIn1 = 32'd9915
; 
32'd187009: dataIn1 = 32'd10114
; 
32'd187010: dataIn1 = 32'd10117
; 
32'd187011: dataIn1 = 32'd9498
; 
32'd187012: dataIn1 = 32'd9501
; 
32'd187013: dataIn1 = 32'd9502
; 
32'd187014: dataIn1 = 32'd9913
; 
32'd187015: dataIn1 = 32'd9914
; 
32'd187016: dataIn1 = 32'd9915
; 
32'd187017: dataIn1 = 32'd3668
; 
32'd187018: dataIn1 = 32'd9500
; 
32'd187019: dataIn1 = 32'd9504
; 
32'd187020: dataIn1 = 32'd9916
; 
32'd187021: dataIn1 = 32'd9917
; 
32'd187022: dataIn1 = 32'd9918
; 
32'd187023: dataIn1 = 32'd9500
; 
32'd187024: dataIn1 = 32'd9503
; 
32'd187025: dataIn1 = 32'd9911
; 
32'd187026: dataIn1 = 32'd9916
; 
32'd187027: dataIn1 = 32'd9917
; 
32'd187028: dataIn1 = 32'd9918
; 
32'd187029: dataIn1 = 32'd9919
; 
32'd187030: dataIn1 = 32'd9503
; 
32'd187031: dataIn1 = 32'd9504
; 
32'd187032: dataIn1 = 32'd9916
; 
32'd187033: dataIn1 = 32'd9917
; 
32'd187034: dataIn1 = 32'd9918
; 
32'd187035: dataIn1 = 32'd9920
; 
32'd187036: dataIn1 = 32'd9921
; 
32'd187037: dataIn1 = 32'd3669
; 
32'd187038: dataIn1 = 32'd9503
; 
32'd187039: dataIn1 = 32'd9911
; 
32'd187040: dataIn1 = 32'd9917
; 
32'd187041: dataIn1 = 32'd9919
; 
32'd187042: dataIn1 = 32'd10174
; 
32'd187043: dataIn1 = 32'd69
; 
32'd187044: dataIn1 = 32'd9504
; 
32'd187045: dataIn1 = 32'd9918
; 
32'd187046: dataIn1 = 32'd9920
; 
32'd187047: dataIn1 = 32'd9921
; 
32'd187048: dataIn1 = 32'd9922
; 
32'd187049: dataIn1 = 32'd9923
; 
32'd187050: dataIn1 = 32'd69
; 
32'd187051: dataIn1 = 32'd9503
; 
32'd187052: dataIn1 = 32'd9918
; 
32'd187053: dataIn1 = 32'd9920
; 
32'd187054: dataIn1 = 32'd9921
; 
32'd187055: dataIn1 = 32'd10173
; 
32'd187056: dataIn1 = 32'd9504
; 
32'd187057: dataIn1 = 32'd9505
; 
32'd187058: dataIn1 = 32'd9506
; 
32'd187059: dataIn1 = 32'd9920
; 
32'd187060: dataIn1 = 32'd9922
; 
32'd187061: dataIn1 = 32'd9923
; 
32'd187062: dataIn1 = 32'd69
; 
32'd187063: dataIn1 = 32'd9505
; 
32'd187064: dataIn1 = 32'd9920
; 
32'd187065: dataIn1 = 32'd9922
; 
32'd187066: dataIn1 = 32'd9923
; 
32'd187067: dataIn1 = 32'd9940
; 
32'd187068: dataIn1 = 32'd9942
; 
32'd187069: dataIn1 = 32'd9508
; 
32'd187070: dataIn1 = 32'd9509
; 
32'd187071: dataIn1 = 32'd9924
; 
32'd187072: dataIn1 = 32'd9925
; 
32'd187073: dataIn1 = 32'd9926
; 
32'd187074: dataIn1 = 32'd9927
; 
32'd187075: dataIn1 = 32'd9928
; 
32'd187076: dataIn1 = 32'd3673
; 
32'd187077: dataIn1 = 32'd9507
; 
32'd187078: dataIn1 = 32'd9509
; 
32'd187079: dataIn1 = 32'd9924
; 
32'd187080: dataIn1 = 32'd9925
; 
32'd187081: dataIn1 = 32'd9926
; 
32'd187082: dataIn1 = 32'd9507
; 
32'd187083: dataIn1 = 32'd9508
; 
32'd187084: dataIn1 = 32'd9924
; 
32'd187085: dataIn1 = 32'd9925
; 
32'd187086: dataIn1 = 32'd9926
; 
32'd187087: dataIn1 = 32'd9929
; 
32'd187088: dataIn1 = 32'd9930
; 
32'd187089: dataIn1 = 32'd2226
; 
32'd187090: dataIn1 = 32'd9509
; 
32'd187091: dataIn1 = 32'd9924
; 
32'd187092: dataIn1 = 32'd9927
; 
32'd187093: dataIn1 = 32'd9928
; 
32'd187094: dataIn1 = 32'd9934
; 
32'd187095: dataIn1 = 32'd9937
; 
32'd187096: dataIn1 = 32'd2226
; 
32'd187097: dataIn1 = 32'd9508
; 
32'd187098: dataIn1 = 32'd9518
; 
32'd187099: dataIn1 = 32'd9924
; 
32'd187100: dataIn1 = 32'd9927
; 
32'd187101: dataIn1 = 32'd9928
; 
32'd187102: dataIn1 = 32'd3674
; 
32'd187103: dataIn1 = 32'd9508
; 
32'd187104: dataIn1 = 32'd9926
; 
32'd187105: dataIn1 = 32'd9929
; 
32'd187106: dataIn1 = 32'd9930
; 
32'd187107: dataIn1 = 32'd9950
; 
32'd187108: dataIn1 = 32'd9951
; 
32'd187109: dataIn1 = 32'd3674
; 
32'd187110: dataIn1 = 32'd9507
; 
32'd187111: dataIn1 = 32'd9926
; 
32'd187112: dataIn1 = 32'd9929
; 
32'd187113: dataIn1 = 32'd9930
; 
32'd187114: dataIn1 = 32'd10175
; 
32'd187115: dataIn1 = 32'd3677
; 
32'd187116: dataIn1 = 32'd9511
; 
32'd187117: dataIn1 = 32'd9931
; 
32'd187118: dataIn1 = 32'd9932
; 
32'd187119: dataIn1 = 32'd9933
; 
32'd187120: dataIn1 = 32'd9941
; 
32'd187121: dataIn1 = 32'd9943
; 
32'd187122: dataIn1 = 32'd3677
; 
32'd187123: dataIn1 = 32'd9510
; 
32'd187124: dataIn1 = 32'd9931
; 
32'd187125: dataIn1 = 32'd9932
; 
32'd187126: dataIn1 = 32'd9933
; 
32'd187127: dataIn1 = 32'd9936
; 
32'd187128: dataIn1 = 32'd9938
; 
32'd187129: dataIn1 = 32'd9510
; 
32'd187130: dataIn1 = 32'd9511
; 
32'd187131: dataIn1 = 32'd9512
; 
32'd187132: dataIn1 = 32'd9931
; 
32'd187133: dataIn1 = 32'd9932
; 
32'd187134: dataIn1 = 32'd9933
; 
32'd187135: dataIn1 = 32'd9509
; 
32'd187136: dataIn1 = 32'd9513
; 
32'd187137: dataIn1 = 32'd9927
; 
32'd187138: dataIn1 = 32'd9934
; 
32'd187139: dataIn1 = 32'd9935
; 
32'd187140: dataIn1 = 32'd9936
; 
32'd187141: dataIn1 = 32'd9937
; 
32'd187142: dataIn1 = 32'd3673
; 
32'd187143: dataIn1 = 32'd9509
; 
32'd187144: dataIn1 = 32'd9510
; 
32'd187145: dataIn1 = 32'd9934
; 
32'd187146: dataIn1 = 32'd9935
; 
32'd187147: dataIn1 = 32'd9936
; 
32'd187148: dataIn1 = 32'd9510
; 
32'd187149: dataIn1 = 32'd9513
; 
32'd187150: dataIn1 = 32'd9932
; 
32'd187151: dataIn1 = 32'd9934
; 
32'd187152: dataIn1 = 32'd9935
; 
32'd187153: dataIn1 = 32'd9936
; 
32'd187154: dataIn1 = 32'd9938
; 
32'd187155: dataIn1 = 32'd2226
; 
32'd187156: dataIn1 = 32'd9513
; 
32'd187157: dataIn1 = 32'd9927
; 
32'd187158: dataIn1 = 32'd9934
; 
32'd187159: dataIn1 = 32'd9937
; 
32'd187160: dataIn1 = 32'd10178
; 
32'd187161: dataIn1 = 32'd3677
; 
32'd187162: dataIn1 = 32'd9513
; 
32'd187163: dataIn1 = 32'd9932
; 
32'd187164: dataIn1 = 32'd9936
; 
32'd187165: dataIn1 = 32'd9938
; 
32'd187166: dataIn1 = 32'd10177
; 
32'd187167: dataIn1 = 32'd3671
; 
32'd187168: dataIn1 = 32'd9505
; 
32'd187169: dataIn1 = 32'd9511
; 
32'd187170: dataIn1 = 32'd9939
; 
32'd187171: dataIn1 = 32'd9940
; 
32'd187172: dataIn1 = 32'd9941
; 
32'd187173: dataIn1 = 32'd9505
; 
32'd187174: dataIn1 = 32'd9514
; 
32'd187175: dataIn1 = 32'd9923
; 
32'd187176: dataIn1 = 32'd9939
; 
32'd187177: dataIn1 = 32'd9940
; 
32'd187178: dataIn1 = 32'd9941
; 
32'd187179: dataIn1 = 32'd9942
; 
32'd187180: dataIn1 = 32'd9511
; 
32'd187181: dataIn1 = 32'd9514
; 
32'd187182: dataIn1 = 32'd9931
; 
32'd187183: dataIn1 = 32'd9939
; 
32'd187184: dataIn1 = 32'd9940
; 
32'd187185: dataIn1 = 32'd9941
; 
32'd187186: dataIn1 = 32'd9943
; 
32'd187187: dataIn1 = 32'd69
; 
32'd187188: dataIn1 = 32'd9514
; 
32'd187189: dataIn1 = 32'd9923
; 
32'd187190: dataIn1 = 32'd9940
; 
32'd187191: dataIn1 = 32'd9942
; 
32'd187192: dataIn1 = 32'd10180
; 
32'd187193: dataIn1 = 32'd3677
; 
32'd187194: dataIn1 = 32'd9514
; 
32'd187195: dataIn1 = 32'd9931
; 
32'd187196: dataIn1 = 32'd9941
; 
32'd187197: dataIn1 = 32'd9943
; 
32'd187198: dataIn1 = 32'd10179
; 
32'd187199: dataIn1 = 32'd9516
; 
32'd187200: dataIn1 = 32'd9517
; 
32'd187201: dataIn1 = 32'd9944
; 
32'd187202: dataIn1 = 32'd9945
; 
32'd187203: dataIn1 = 32'd9946
; 
32'd187204: dataIn1 = 32'd9947
; 
32'd187205: dataIn1 = 32'd9948
; 
32'd187206: dataIn1 = 32'd3679
; 
32'd187207: dataIn1 = 32'd9515
; 
32'd187208: dataIn1 = 32'd9517
; 
32'd187209: dataIn1 = 32'd9944
; 
32'd187210: dataIn1 = 32'd9945
; 
32'd187211: dataIn1 = 32'd9946
; 
32'd187212: dataIn1 = 32'd9515
; 
32'd187213: dataIn1 = 32'd9516
; 
32'd187214: dataIn1 = 32'd9944
; 
32'd187215: dataIn1 = 32'd9945
; 
32'd187216: dataIn1 = 32'd9946
; 
32'd187217: dataIn1 = 32'd9949
; 
32'd187218: dataIn1 = 32'd9950
; 
32'd187219: dataIn1 = 32'd3678
; 
32'd187220: dataIn1 = 32'd9517
; 
32'd187221: dataIn1 = 32'd9944
; 
32'd187222: dataIn1 = 32'd9947
; 
32'd187223: dataIn1 = 32'd9948
; 
32'd187224: dataIn1 = 32'd9952
; 
32'd187225: dataIn1 = 32'd9953
; 
32'd187226: dataIn1 = 32'd3678
; 
32'd187227: dataIn1 = 32'd9516
; 
32'd187228: dataIn1 = 32'd9944
; 
32'd187229: dataIn1 = 32'd9947
; 
32'd187230: dataIn1 = 32'd9948
; 
32'd187231: dataIn1 = 32'd10182
; 
32'd187232: dataIn1 = 32'd3674
; 
32'd187233: dataIn1 = 32'd9516
; 
32'd187234: dataIn1 = 32'd9946
; 
32'd187235: dataIn1 = 32'd9949
; 
32'd187236: dataIn1 = 32'd9950
; 
32'd187237: dataIn1 = 32'd10181
; 
32'd187238: dataIn1 = 32'd3674
; 
32'd187239: dataIn1 = 32'd9515
; 
32'd187240: dataIn1 = 32'd9929
; 
32'd187241: dataIn1 = 32'd9946
; 
32'd187242: dataIn1 = 32'd9949
; 
32'd187243: dataIn1 = 32'd9950
; 
32'd187244: dataIn1 = 32'd9951
; 
32'd187245: dataIn1 = 32'd9508
; 
32'd187246: dataIn1 = 32'd9515
; 
32'd187247: dataIn1 = 32'd9518
; 
32'd187248: dataIn1 = 32'd9929
; 
32'd187249: dataIn1 = 32'd9950
; 
32'd187250: dataIn1 = 32'd9951
; 
32'd187251: dataIn1 = 32'd9517
; 
32'd187252: dataIn1 = 32'd9519
; 
32'd187253: dataIn1 = 32'd9520
; 
32'd187254: dataIn1 = 32'd9947
; 
32'd187255: dataIn1 = 32'd9952
; 
32'd187256: dataIn1 = 32'd9953
; 
32'd187257: dataIn1 = 32'd3678
; 
32'd187258: dataIn1 = 32'd9520
; 
32'd187259: dataIn1 = 32'd9947
; 
32'd187260: dataIn1 = 32'd9952
; 
32'd187261: dataIn1 = 32'd9953
; 
32'd187262: dataIn1 = 32'd9959
; 
32'd187263: dataIn1 = 32'd9962
; 
32'd187264: dataIn1 = 32'd3684
; 
32'd187265: dataIn1 = 32'd9522
; 
32'd187266: dataIn1 = 32'd9954
; 
32'd187267: dataIn1 = 32'd9955
; 
32'd187268: dataIn1 = 32'd9956
; 
32'd187269: dataIn1 = 32'd9961
; 
32'd187270: dataIn1 = 32'd9963
; 
32'd187271: dataIn1 = 32'd3684
; 
32'd187272: dataIn1 = 32'd9521
; 
32'd187273: dataIn1 = 32'd9954
; 
32'd187274: dataIn1 = 32'd9955
; 
32'd187275: dataIn1 = 32'd9956
; 
32'd187276: dataIn1 = 32'd9957
; 
32'd187277: dataIn1 = 32'd9958
; 
32'd187278: dataIn1 = 32'd9521
; 
32'd187279: dataIn1 = 32'd9522
; 
32'd187280: dataIn1 = 32'd9523
; 
32'd187281: dataIn1 = 32'd9954
; 
32'd187282: dataIn1 = 32'd9955
; 
32'd187283: dataIn1 = 32'd9956
; 
32'd187284: dataIn1 = 32'd3684
; 
32'd187285: dataIn1 = 32'd9524
; 
32'd187286: dataIn1 = 32'd9955
; 
32'd187287: dataIn1 = 32'd9957
; 
32'd187288: dataIn1 = 32'd9958
; 
32'd187289: dataIn1 = 32'd9979
; 
32'd187290: dataIn1 = 32'd9982
; 
32'd187291: dataIn1 = 32'd9521
; 
32'd187292: dataIn1 = 32'd9524
; 
32'd187293: dataIn1 = 32'd9525
; 
32'd187294: dataIn1 = 32'd9955
; 
32'd187295: dataIn1 = 32'd9957
; 
32'd187296: dataIn1 = 32'd9958
; 
32'd187297: dataIn1 = 32'd9520
; 
32'd187298: dataIn1 = 32'd9522
; 
32'd187299: dataIn1 = 32'd9953
; 
32'd187300: dataIn1 = 32'd9959
; 
32'd187301: dataIn1 = 32'd9960
; 
32'd187302: dataIn1 = 32'd9961
; 
32'd187303: dataIn1 = 32'd9962
; 
32'd187304: dataIn1 = 32'd70
; 
32'd187305: dataIn1 = 32'd9520
; 
32'd187306: dataIn1 = 32'd9526
; 
32'd187307: dataIn1 = 32'd9959
; 
32'd187308: dataIn1 = 32'd9960
; 
32'd187309: dataIn1 = 32'd9961
; 
32'd187310: dataIn1 = 32'd9522
; 
32'd187311: dataIn1 = 32'd9526
; 
32'd187312: dataIn1 = 32'd9954
; 
32'd187313: dataIn1 = 32'd9959
; 
32'd187314: dataIn1 = 32'd9960
; 
32'd187315: dataIn1 = 32'd9961
; 
32'd187316: dataIn1 = 32'd9963
; 
32'd187317: dataIn1 = 32'd3678
; 
32'd187318: dataIn1 = 32'd9522
; 
32'd187319: dataIn1 = 32'd9523
; 
32'd187320: dataIn1 = 32'd9953
; 
32'd187321: dataIn1 = 32'd9959
; 
32'd187322: dataIn1 = 32'd9962
; 
32'd187323: dataIn1 = 32'd3684
; 
32'd187324: dataIn1 = 32'd9526
; 
32'd187325: dataIn1 = 32'd9954
; 
32'd187326: dataIn1 = 32'd9961
; 
32'd187327: dataIn1 = 32'd9963
; 
32'd187328: dataIn1 = 32'd10184
; 
32'd187329: dataIn1 = 32'd9528
; 
32'd187330: dataIn1 = 32'd9529
; 
32'd187331: dataIn1 = 32'd9964
; 
32'd187332: dataIn1 = 32'd9965
; 
32'd187333: dataIn1 = 32'd9966
; 
32'd187334: dataIn1 = 32'd9967
; 
32'd187335: dataIn1 = 32'd9968
; 
32'd187336: dataIn1 = 32'd9527
; 
32'd187337: dataIn1 = 32'd9529
; 
32'd187338: dataIn1 = 32'd9964
; 
32'd187339: dataIn1 = 32'd9965
; 
32'd187340: dataIn1 = 32'd9966
; 
32'd187341: dataIn1 = 32'd9969
; 
32'd187342: dataIn1 = 32'd9970
; 
32'd187343: dataIn1 = 32'd3689
; 
32'd187344: dataIn1 = 32'd9527
; 
32'd187345: dataIn1 = 32'd9528
; 
32'd187346: dataIn1 = 32'd9964
; 
32'd187347: dataIn1 = 32'd9965
; 
32'd187348: dataIn1 = 32'd9966
; 
32'd187349: dataIn1 = 32'd3687
; 
32'd187350: dataIn1 = 32'd9529
; 
32'd187351: dataIn1 = 32'd9533
; 
32'd187352: dataIn1 = 32'd9964
; 
32'd187353: dataIn1 = 32'd9967
; 
32'd187354: dataIn1 = 32'd9968
; 
32'd187355: dataIn1 = 32'd3687
; 
32'd187356: dataIn1 = 32'd9528
; 
32'd187357: dataIn1 = 32'd9964
; 
32'd187358: dataIn1 = 32'd9967
; 
32'd187359: dataIn1 = 32'd9968
; 
32'd187360: dataIn1 = 32'd9971
; 
32'd187361: dataIn1 = 32'd9974
; 
32'd187362: dataIn1 = 32'd3688
; 
32'd187363: dataIn1 = 32'd9529
; 
32'd187364: dataIn1 = 32'd9965
; 
32'd187365: dataIn1 = 32'd9969
; 
32'd187366: dataIn1 = 32'd9970
; 
32'd187367: dataIn1 = 32'd9977
; 
32'd187368: dataIn1 = 32'd9978
; 
32'd187369: dataIn1 = 32'd3688
; 
32'd187370: dataIn1 = 32'd9527
; 
32'd187371: dataIn1 = 32'd9965
; 
32'd187372: dataIn1 = 32'd9969
; 
32'd187373: dataIn1 = 32'd9970
; 
32'd187374: dataIn1 = 32'd10186
; 
32'd187375: dataIn1 = 32'd9528
; 
32'd187376: dataIn1 = 32'd9531
; 
32'd187377: dataIn1 = 32'd9968
; 
32'd187378: dataIn1 = 32'd9971
; 
32'd187379: dataIn1 = 32'd9972
; 
32'd187380: dataIn1 = 32'd9973
; 
32'd187381: dataIn1 = 32'd9974
; 
32'd187382: dataIn1 = 32'd9530
; 
32'd187383: dataIn1 = 32'd9531
; 
32'd187384: dataIn1 = 32'd9971
; 
32'd187385: dataIn1 = 32'd9972
; 
32'd187386: dataIn1 = 32'd9973
; 
32'd187387: dataIn1 = 32'd9975
; 
32'd187388: dataIn1 = 32'd9976
; 
32'd187389: dataIn1 = 32'd3689
; 
32'd187390: dataIn1 = 32'd9528
; 
32'd187391: dataIn1 = 32'd9530
; 
32'd187392: dataIn1 = 32'd9971
; 
32'd187393: dataIn1 = 32'd9972
; 
32'd187394: dataIn1 = 32'd9973
; 
32'd187395: dataIn1 = 32'd3687
; 
32'd187396: dataIn1 = 32'd9531
; 
32'd187397: dataIn1 = 32'd9968
; 
32'd187398: dataIn1 = 32'd9971
; 
32'd187399: dataIn1 = 32'd9974
; 
32'd187400: dataIn1 = 32'd10188
; 
32'd187401: dataIn1 = 32'd2230
; 
32'd187402: dataIn1 = 32'd9531
; 
32'd187403: dataIn1 = 32'd9972
; 
32'd187404: dataIn1 = 32'd9975
; 
32'd187405: dataIn1 = 32'd9976
; 
32'd187406: dataIn1 = 32'd10187
; 
32'd187407: dataIn1 = 32'd2230
; 
32'd187408: dataIn1 = 32'd9530
; 
32'd187409: dataIn1 = 32'd9972
; 
32'd187410: dataIn1 = 32'd9975
; 
32'd187411: dataIn1 = 32'd9976
; 
32'd187412: dataIn1 = 32'd9984
; 
32'd187413: dataIn1 = 32'd9985
; 
32'd187414: dataIn1 = 32'd9529
; 
32'd187415: dataIn1 = 32'd9532
; 
32'd187416: dataIn1 = 32'd9533
; 
32'd187417: dataIn1 = 32'd9969
; 
32'd187418: dataIn1 = 32'd9977
; 
32'd187419: dataIn1 = 32'd9978
; 
32'd187420: dataIn1 = 32'd3688
; 
32'd187421: dataIn1 = 32'd9532
; 
32'd187422: dataIn1 = 32'd9969
; 
32'd187423: dataIn1 = 32'd9977
; 
32'd187424: dataIn1 = 32'd9978
; 
32'd187425: dataIn1 = 32'd9980
; 
32'd187426: dataIn1 = 32'd9983
; 
32'd187427: dataIn1 = 32'd9524
; 
32'd187428: dataIn1 = 32'd9534
; 
32'd187429: dataIn1 = 32'd9957
; 
32'd187430: dataIn1 = 32'd9979
; 
32'd187431: dataIn1 = 32'd9980
; 
32'd187432: dataIn1 = 32'd9981
; 
32'd187433: dataIn1 = 32'd9982
; 
32'd187434: dataIn1 = 32'd9532
; 
32'd187435: dataIn1 = 32'd9534
; 
32'd187436: dataIn1 = 32'd9978
; 
32'd187437: dataIn1 = 32'd9979
; 
32'd187438: dataIn1 = 32'd9980
; 
32'd187439: dataIn1 = 32'd9981
; 
32'd187440: dataIn1 = 32'd9983
; 
32'd187441: dataIn1 = 32'd2228
; 
32'd187442: dataIn1 = 32'd9524
; 
32'd187443: dataIn1 = 32'd9532
; 
32'd187444: dataIn1 = 32'd9979
; 
32'd187445: dataIn1 = 32'd9980
; 
32'd187446: dataIn1 = 32'd9981
; 
32'd187447: dataIn1 = 32'd3684
; 
32'd187448: dataIn1 = 32'd9534
; 
32'd187449: dataIn1 = 32'd9957
; 
32'd187450: dataIn1 = 32'd9979
; 
32'd187451: dataIn1 = 32'd9982
; 
32'd187452: dataIn1 = 32'd10184
; 
32'd187453: dataIn1 = 32'd3688
; 
32'd187454: dataIn1 = 32'd9534
; 
32'd187455: dataIn1 = 32'd9978
; 
32'd187456: dataIn1 = 32'd9980
; 
32'd187457: dataIn1 = 32'd9983
; 
32'd187458: dataIn1 = 32'd10189
; 
32'd187459: dataIn1 = 32'd2230
; 
32'd187460: dataIn1 = 32'd9536
; 
32'd187461: dataIn1 = 32'd9976
; 
32'd187462: dataIn1 = 32'd9984
; 
32'd187463: dataIn1 = 32'd9985
; 
32'd187464: dataIn1 = 32'd10000
; 
32'd187465: dataIn1 = 32'd10001
; 
32'd187466: dataIn1 = 32'd9530
; 
32'd187467: dataIn1 = 32'd9535
; 
32'd187468: dataIn1 = 32'd9536
; 
32'd187469: dataIn1 = 32'd9976
; 
32'd187470: dataIn1 = 32'd9984
; 
32'd187471: dataIn1 = 32'd9985
; 
32'd187472: dataIn1 = 32'd3695
; 
32'd187473: dataIn1 = 32'd9539
; 
32'd187474: dataIn1 = 32'd9986
; 
32'd187475: dataIn1 = 32'd9987
; 
32'd187476: dataIn1 = 32'd9988
; 
32'd187477: dataIn1 = 32'd9996
; 
32'd187478: dataIn1 = 32'd9998
; 
32'd187479: dataIn1 = 32'd9537
; 
32'd187480: dataIn1 = 32'd9538
; 
32'd187481: dataIn1 = 32'd9539
; 
32'd187482: dataIn1 = 32'd9986
; 
32'd187483: dataIn1 = 32'd9987
; 
32'd187484: dataIn1 = 32'd9988
; 
32'd187485: dataIn1 = 32'd3695
; 
32'd187486: dataIn1 = 32'd9537
; 
32'd187487: dataIn1 = 32'd9986
; 
32'd187488: dataIn1 = 32'd9987
; 
32'd187489: dataIn1 = 32'd9988
; 
32'd187490: dataIn1 = 32'd9990
; 
32'd187491: dataIn1 = 32'd9992
; 
32'd187492: dataIn1 = 32'd2231
; 
32'd187493: dataIn1 = 32'd9540
; 
32'd187494: dataIn1 = 32'd9541
; 
32'd187495: dataIn1 = 32'd9989
; 
32'd187496: dataIn1 = 32'd9990
; 
32'd187497: dataIn1 = 32'd9991
; 
32'd187498: dataIn1 = 32'd9537
; 
32'd187499: dataIn1 = 32'd9541
; 
32'd187500: dataIn1 = 32'd9988
; 
32'd187501: dataIn1 = 32'd9989
; 
32'd187502: dataIn1 = 32'd9990
; 
32'd187503: dataIn1 = 32'd9991
; 
32'd187504: dataIn1 = 32'd9992
; 
32'd187505: dataIn1 = 32'd9537
; 
32'd187506: dataIn1 = 32'd9540
; 
32'd187507: dataIn1 = 32'd9989
; 
32'd187508: dataIn1 = 32'd9990
; 
32'd187509: dataIn1 = 32'd9991
; 
32'd187510: dataIn1 = 32'd9993
; 
32'd187511: dataIn1 = 32'd9994
; 
32'd187512: dataIn1 = 32'd3695
; 
32'd187513: dataIn1 = 32'd9541
; 
32'd187514: dataIn1 = 32'd9988
; 
32'd187515: dataIn1 = 32'd9990
; 
32'd187516: dataIn1 = 32'd9992
; 
32'd187517: dataIn1 = 32'd10190
; 
32'd187518: dataIn1 = 32'd3696
; 
32'd187519: dataIn1 = 32'd9540
; 
32'd187520: dataIn1 = 32'd9991
; 
32'd187521: dataIn1 = 32'd9993
; 
32'd187522: dataIn1 = 32'd9994
; 
32'd187523: dataIn1 = 32'd10007
; 
32'd187524: dataIn1 = 32'd10009
; 
32'd187525: dataIn1 = 32'd3696
; 
32'd187526: dataIn1 = 32'd9537
; 
32'd187527: dataIn1 = 32'd9538
; 
32'd187528: dataIn1 = 32'd9991
; 
32'd187529: dataIn1 = 32'd9993
; 
32'd187530: dataIn1 = 32'd9994
; 
32'd187531: dataIn1 = 32'd3694
; 
32'd187532: dataIn1 = 32'd9539
; 
32'd187533: dataIn1 = 32'd9543
; 
32'd187534: dataIn1 = 32'd9995
; 
32'd187535: dataIn1 = 32'd9996
; 
32'd187536: dataIn1 = 32'd9997
; 
32'd187537: dataIn1 = 32'd9539
; 
32'd187538: dataIn1 = 32'd9542
; 
32'd187539: dataIn1 = 32'd9986
; 
32'd187540: dataIn1 = 32'd9995
; 
32'd187541: dataIn1 = 32'd9996
; 
32'd187542: dataIn1 = 32'd9997
; 
32'd187543: dataIn1 = 32'd9998
; 
32'd187544: dataIn1 = 32'd9542
; 
32'd187545: dataIn1 = 32'd9543
; 
32'd187546: dataIn1 = 32'd9995
; 
32'd187547: dataIn1 = 32'd9996
; 
32'd187548: dataIn1 = 32'd9997
; 
32'd187549: dataIn1 = 32'd9999
; 
32'd187550: dataIn1 = 32'd10000
; 
32'd187551: dataIn1 = 32'd3695
; 
32'd187552: dataIn1 = 32'd9542
; 
32'd187553: dataIn1 = 32'd9544
; 
32'd187554: dataIn1 = 32'd9986
; 
32'd187555: dataIn1 = 32'd9996
; 
32'd187556: dataIn1 = 32'd9998
; 
32'd187557: dataIn1 = 32'd2230
; 
32'd187558: dataIn1 = 32'd9543
; 
32'd187559: dataIn1 = 32'd9997
; 
32'd187560: dataIn1 = 32'd9999
; 
32'd187561: dataIn1 = 32'd10000
; 
32'd187562: dataIn1 = 32'd10187
; 
32'd187563: dataIn1 = 32'd2230
; 
32'd187564: dataIn1 = 32'd9542
; 
32'd187565: dataIn1 = 32'd9984
; 
32'd187566: dataIn1 = 32'd9997
; 
32'd187567: dataIn1 = 32'd9999
; 
32'd187568: dataIn1 = 32'd10000
; 
32'd187569: dataIn1 = 32'd10001
; 
32'd187570: dataIn1 = 32'd9536
; 
32'd187571: dataIn1 = 32'd9542
; 
32'd187572: dataIn1 = 32'd9544
; 
32'd187573: dataIn1 = 32'd9984
; 
32'd187574: dataIn1 = 32'd10000
; 
32'd187575: dataIn1 = 32'd10001
; 
32'd187576: dataIn1 = 32'd3698
; 
32'd187577: dataIn1 = 32'd9547
; 
32'd187578: dataIn1 = 32'd10002
; 
32'd187579: dataIn1 = 32'd10003
; 
32'd187580: dataIn1 = 32'd10004
; 
32'd187581: dataIn1 = 32'd10010
; 
32'd187582: dataIn1 = 32'd10011
; 
32'd187583: dataIn1 = 32'd9545
; 
32'd187584: dataIn1 = 32'd9546
; 
32'd187585: dataIn1 = 32'd9547
; 
32'd187586: dataIn1 = 32'd10002
; 
32'd187587: dataIn1 = 32'd10003
; 
32'd187588: dataIn1 = 32'd10004
; 
32'd187589: dataIn1 = 32'd3698
; 
32'd187590: dataIn1 = 32'd9545
; 
32'd187591: dataIn1 = 32'd10002
; 
32'd187592: dataIn1 = 32'd10003
; 
32'd187593: dataIn1 = 32'd10004
; 
32'd187594: dataIn1 = 32'd10006
; 
32'd187595: dataIn1 = 32'd10008
; 
32'd187596: dataIn1 = 32'd2231
; 
32'd187597: dataIn1 = 32'd9540
; 
32'd187598: dataIn1 = 32'd9548
; 
32'd187599: dataIn1 = 32'd10005
; 
32'd187600: dataIn1 = 32'd10006
; 
32'd187601: dataIn1 = 32'd10007
; 
32'd187602: dataIn1 = 32'd9545
; 
32'd187603: dataIn1 = 32'd9548
; 
32'd187604: dataIn1 = 32'd10004
; 
32'd187605: dataIn1 = 32'd10005
; 
32'd187606: dataIn1 = 32'd10006
; 
32'd187607: dataIn1 = 32'd10007
; 
32'd187608: dataIn1 = 32'd10008
; 
32'd187609: dataIn1 = 32'd9540
; 
32'd187610: dataIn1 = 32'd9545
; 
32'd187611: dataIn1 = 32'd9993
; 
32'd187612: dataIn1 = 32'd10005
; 
32'd187613: dataIn1 = 32'd10006
; 
32'd187614: dataIn1 = 32'd10007
; 
32'd187615: dataIn1 = 32'd10009
; 
32'd187616: dataIn1 = 32'd3698
; 
32'd187617: dataIn1 = 32'd9548
; 
32'd187618: dataIn1 = 32'd10004
; 
32'd187619: dataIn1 = 32'd10006
; 
32'd187620: dataIn1 = 32'd10008
; 
32'd187621: dataIn1 = 32'd10194
; 
32'd187622: dataIn1 = 32'd3696
; 
32'd187623: dataIn1 = 32'd9545
; 
32'd187624: dataIn1 = 32'd9546
; 
32'd187625: dataIn1 = 32'd9993
; 
32'd187626: dataIn1 = 32'd10007
; 
32'd187627: dataIn1 = 32'd10009
; 
32'd187628: dataIn1 = 32'd9547
; 
32'd187629: dataIn1 = 32'd9549
; 
32'd187630: dataIn1 = 32'd9550
; 
32'd187631: dataIn1 = 32'd10002
; 
32'd187632: dataIn1 = 32'd10010
; 
32'd187633: dataIn1 = 32'd10011
; 
32'd187634: dataIn1 = 32'd3698
; 
32'd187635: dataIn1 = 32'd9549
; 
32'd187636: dataIn1 = 32'd10002
; 
32'd187637: dataIn1 = 32'd10010
; 
32'd187638: dataIn1 = 32'd10011
; 
32'd187639: dataIn1 = 32'd10013
; 
32'd187640: dataIn1 = 32'd10015
; 
32'd187641: dataIn1 = 32'd61
; 
32'd187642: dataIn1 = 32'd9549
; 
32'd187643: dataIn1 = 32'd9552
; 
32'd187644: dataIn1 = 32'd10012
; 
32'd187645: dataIn1 = 32'd10013
; 
32'd187646: dataIn1 = 32'd10014
; 
32'd187647: dataIn1 = 32'd9549
; 
32'd187648: dataIn1 = 32'd9551
; 
32'd187649: dataIn1 = 32'd10011
; 
32'd187650: dataIn1 = 32'd10012
; 
32'd187651: dataIn1 = 32'd10013
; 
32'd187652: dataIn1 = 32'd10014
; 
32'd187653: dataIn1 = 32'd10015
; 
32'd187654: dataIn1 = 32'd9551
; 
32'd187655: dataIn1 = 32'd9552
; 
32'd187656: dataIn1 = 32'd10012
; 
32'd187657: dataIn1 = 32'd10013
; 
32'd187658: dataIn1 = 32'd10014
; 
32'd187659: dataIn1 = 32'd10016
; 
32'd187660: dataIn1 = 32'd10017
; 
32'd187661: dataIn1 = 32'd3698
; 
32'd187662: dataIn1 = 32'd9551
; 
32'd187663: dataIn1 = 32'd10011
; 
32'd187664: dataIn1 = 32'd10013
; 
32'd187665: dataIn1 = 32'd10015
; 
32'd187666: dataIn1 = 32'd10194
; 
32'd187667: dataIn1 = 32'd3702
; 
32'd187668: dataIn1 = 32'd9552
; 
32'd187669: dataIn1 = 32'd10014
; 
32'd187670: dataIn1 = 32'd10016
; 
32'd187671: dataIn1 = 32'd10017
; 
32'd187672: dataIn1 = 32'd10022
; 
32'd187673: dataIn1 = 32'd10024
; 
32'd187674: dataIn1 = 32'd3702
; 
32'd187675: dataIn1 = 32'd9551
; 
32'd187676: dataIn1 = 32'd10014
; 
32'd187677: dataIn1 = 32'd10016
; 
32'd187678: dataIn1 = 32'd10017
; 
32'd187679: dataIn1 = 32'd10195
; 
32'd187680: dataIn1 = 32'd3625
; 
32'd187681: dataIn1 = 32'd9554
; 
32'd187682: dataIn1 = 32'd9882
; 
32'd187683: dataIn1 = 32'd10018
; 
32'd187684: dataIn1 = 32'd10019
; 
32'd187685: dataIn1 = 32'd10020
; 
32'd187686: dataIn1 = 32'd10026
; 
32'd187687: dataIn1 = 32'd3625
; 
32'd187688: dataIn1 = 32'd9553
; 
32'd187689: dataIn1 = 32'd10018
; 
32'd187690: dataIn1 = 32'd10019
; 
32'd187691: dataIn1 = 32'd10020
; 
32'd187692: dataIn1 = 32'd10023
; 
32'd187693: dataIn1 = 32'd10025
; 
32'd187694: dataIn1 = 32'd9553
; 
32'd187695: dataIn1 = 32'd9554
; 
32'd187696: dataIn1 = 32'd9555
; 
32'd187697: dataIn1 = 32'd10018
; 
32'd187698: dataIn1 = 32'd10019
; 
32'd187699: dataIn1 = 32'd10020
; 
32'd187700: dataIn1 = 32'd61
; 
32'd187701: dataIn1 = 32'd9552
; 
32'd187702: dataIn1 = 32'd9556
; 
32'd187703: dataIn1 = 32'd10021
; 
32'd187704: dataIn1 = 32'd10022
; 
32'd187705: dataIn1 = 32'd10023
; 
32'd187706: dataIn1 = 32'd9552
; 
32'd187707: dataIn1 = 32'd9553
; 
32'd187708: dataIn1 = 32'd10016
; 
32'd187709: dataIn1 = 32'd10021
; 
32'd187710: dataIn1 = 32'd10022
; 
32'd187711: dataIn1 = 32'd10023
; 
32'd187712: dataIn1 = 32'd10024
; 
32'd187713: dataIn1 = 32'd9553
; 
32'd187714: dataIn1 = 32'd9556
; 
32'd187715: dataIn1 = 32'd10019
; 
32'd187716: dataIn1 = 32'd10021
; 
32'd187717: dataIn1 = 32'd10022
; 
32'd187718: dataIn1 = 32'd10023
; 
32'd187719: dataIn1 = 32'd10025
; 
32'd187720: dataIn1 = 32'd3702
; 
32'd187721: dataIn1 = 32'd9553
; 
32'd187722: dataIn1 = 32'd9555
; 
32'd187723: dataIn1 = 32'd10016
; 
32'd187724: dataIn1 = 32'd10022
; 
32'd187725: dataIn1 = 32'd10024
; 
32'd187726: dataIn1 = 32'd3625
; 
32'd187727: dataIn1 = 32'd9556
; 
32'd187728: dataIn1 = 32'd10019
; 
32'd187729: dataIn1 = 32'd10023
; 
32'd187730: dataIn1 = 32'd10025
; 
32'd187731: dataIn1 = 32'd10164
; 
32'd187732: dataIn1 = 32'd9486
; 
32'd187733: dataIn1 = 32'd9554
; 
32'd187734: dataIn1 = 32'd9557
; 
32'd187735: dataIn1 = 32'd9882
; 
32'd187736: dataIn1 = 32'd10018
; 
32'd187737: dataIn1 = 32'd10026
; 
32'd187738: dataIn1 = 32'd66
; 
32'd187739: dataIn1 = 32'd9559
; 
32'd187740: dataIn1 = 32'd9560
; 
32'd187741: dataIn1 = 32'd10027
; 
32'd187742: dataIn1 = 32'd10028
; 
32'd187743: dataIn1 = 32'd10029
; 
32'd187744: dataIn1 = 32'd9558
; 
32'd187745: dataIn1 = 32'd9560
; 
32'd187746: dataIn1 = 32'd10027
; 
32'd187747: dataIn1 = 32'd10028
; 
32'd187748: dataIn1 = 32'd10029
; 
32'd187749: dataIn1 = 32'd10030
; 
32'd187750: dataIn1 = 32'd10031
; 
32'd187751: dataIn1 = 32'd9558
; 
32'd187752: dataIn1 = 32'd9559
; 
32'd187753: dataIn1 = 32'd10027
; 
32'd187754: dataIn1 = 32'd10028
; 
32'd187755: dataIn1 = 32'd10029
; 
32'd187756: dataIn1 = 32'd10032
; 
32'd187757: dataIn1 = 32'd10033
; 
32'd187758: dataIn1 = 32'd3735
; 
32'd187759: dataIn1 = 32'd9560
; 
32'd187760: dataIn1 = 32'd10028
; 
32'd187761: dataIn1 = 32'd10030
; 
32'd187762: dataIn1 = 32'd10031
; 
32'd187763: dataIn1 = 32'd3735
; 
32'd187764: dataIn1 = 32'd9558
; 
32'd187765: dataIn1 = 32'd10028
; 
32'd187766: dataIn1 = 32'd10030
; 
32'd187767: dataIn1 = 32'd10031
; 
32'd187768: dataIn1 = 32'd10198
; 
32'd187769: dataIn1 = 32'd10287
; 
32'd187770: dataIn1 = 32'd3736
; 
32'd187771: dataIn1 = 32'd9559
; 
32'd187772: dataIn1 = 32'd10029
; 
32'd187773: dataIn1 = 32'd10032
; 
32'd187774: dataIn1 = 32'd10033
; 
32'd187775: dataIn1 = 32'd10047
; 
32'd187776: dataIn1 = 32'd10048
; 
32'd187777: dataIn1 = 32'd3736
; 
32'd187778: dataIn1 = 32'd9558
; 
32'd187779: dataIn1 = 32'd10029
; 
32'd187780: dataIn1 = 32'd10032
; 
32'd187781: dataIn1 = 32'd10033
; 
32'd187782: dataIn1 = 32'd10197
; 
32'd187783: dataIn1 = 32'd10198
; 
32'd187784: dataIn1 = 32'd9562
; 
32'd187785: dataIn1 = 32'd9563
; 
32'd187786: dataIn1 = 32'd10034
; 
32'd187787: dataIn1 = 32'd10035
; 
32'd187788: dataIn1 = 32'd10036
; 
32'd187789: dataIn1 = 32'd10037
; 
32'd187790: dataIn1 = 32'd10038
; 
32'd187791: dataIn1 = 32'd9561
; 
32'd187792: dataIn1 = 32'd9563
; 
32'd187793: dataIn1 = 32'd10034
; 
32'd187794: dataIn1 = 32'd10035
; 
32'd187795: dataIn1 = 32'd10036
; 
32'd187796: dataIn1 = 32'd10039
; 
32'd187797: dataIn1 = 32'd10040
; 
32'd187798: dataIn1 = 32'd3743
; 
32'd187799: dataIn1 = 32'd9561
; 
32'd187800: dataIn1 = 32'd9562
; 
32'd187801: dataIn1 = 32'd10034
; 
32'd187802: dataIn1 = 32'd10035
; 
32'd187803: dataIn1 = 32'd10036
; 
32'd187804: dataIn1 = 32'd3741
; 
32'd187805: dataIn1 = 32'd9563
; 
32'd187806: dataIn1 = 32'd10034
; 
32'd187807: dataIn1 = 32'd10037
; 
32'd187808: dataIn1 = 32'd10038
; 
32'd187809: dataIn1 = 32'd10045
; 
32'd187810: dataIn1 = 32'd10049
; 
32'd187811: dataIn1 = 32'd3741
; 
32'd187812: dataIn1 = 32'd9562
; 
32'd187813: dataIn1 = 32'd10034
; 
32'd187814: dataIn1 = 32'd10037
; 
32'd187815: dataIn1 = 32'd10038
; 
32'd187816: dataIn1 = 32'd10200
; 
32'd187817: dataIn1 = 32'd2217
; 
32'd187818: dataIn1 = 32'd9563
; 
32'd187819: dataIn1 = 32'd9568
; 
32'd187820: dataIn1 = 32'd10035
; 
32'd187821: dataIn1 = 32'd10039
; 
32'd187822: dataIn1 = 32'd10040
; 
32'd187823: dataIn1 = 32'd2217
; 
32'd187824: dataIn1 = 32'd9561
; 
32'd187825: dataIn1 = 32'd10035
; 
32'd187826: dataIn1 = 32'd10039
; 
32'd187827: dataIn1 = 32'd10040
; 
32'd187828: dataIn1 = 32'd10054
; 
32'd187829: dataIn1 = 32'd10057
; 
32'd187830: dataIn1 = 32'd9565
; 
32'd187831: dataIn1 = 32'd9566
; 
32'd187832: dataIn1 = 32'd10041
; 
32'd187833: dataIn1 = 32'd10042
; 
32'd187834: dataIn1 = 32'd10043
; 
32'd187835: dataIn1 = 32'd10044
; 
32'd187836: dataIn1 = 32'd10045
; 
32'd187837: dataIn1 = 32'd9564
; 
32'd187838: dataIn1 = 32'd9566
; 
32'd187839: dataIn1 = 32'd10041
; 
32'd187840: dataIn1 = 32'd10042
; 
32'd187841: dataIn1 = 32'd10043
; 
32'd187842: dataIn1 = 32'd10046
; 
32'd187843: dataIn1 = 32'd10047
; 
32'd187844: dataIn1 = 32'd3744
; 
32'd187845: dataIn1 = 32'd9564
; 
32'd187846: dataIn1 = 32'd9565
; 
32'd187847: dataIn1 = 32'd10041
; 
32'd187848: dataIn1 = 32'd10042
; 
32'd187849: dataIn1 = 32'd10043
; 
32'd187850: dataIn1 = 32'd3741
; 
32'd187851: dataIn1 = 32'd9566
; 
32'd187852: dataIn1 = 32'd10041
; 
32'd187853: dataIn1 = 32'd10044
; 
32'd187854: dataIn1 = 32'd10045
; 
32'd187855: dataIn1 = 32'd10202
; 
32'd187856: dataIn1 = 32'd3741
; 
32'd187857: dataIn1 = 32'd9565
; 
32'd187858: dataIn1 = 32'd10037
; 
32'd187859: dataIn1 = 32'd10041
; 
32'd187860: dataIn1 = 32'd10044
; 
32'd187861: dataIn1 = 32'd10045
; 
32'd187862: dataIn1 = 32'd10049
; 
32'd187863: dataIn1 = 32'd3736
; 
32'd187864: dataIn1 = 32'd9566
; 
32'd187865: dataIn1 = 32'd10042
; 
32'd187866: dataIn1 = 32'd10046
; 
32'd187867: dataIn1 = 32'd10047
; 
32'd187868: dataIn1 = 32'd10201
; 
32'd187869: dataIn1 = 32'd3736
; 
32'd187870: dataIn1 = 32'd9564
; 
32'd187871: dataIn1 = 32'd10032
; 
32'd187872: dataIn1 = 32'd10042
; 
32'd187873: dataIn1 = 32'd10046
; 
32'd187874: dataIn1 = 32'd10047
; 
32'd187875: dataIn1 = 32'd10048
; 
32'd187876: dataIn1 = 32'd9559
; 
32'd187877: dataIn1 = 32'd9564
; 
32'd187878: dataIn1 = 32'd9567
; 
32'd187879: dataIn1 = 32'd10032
; 
32'd187880: dataIn1 = 32'd10047
; 
32'd187881: dataIn1 = 32'd10048
; 
32'd187882: dataIn1 = 32'd9563
; 
32'd187883: dataIn1 = 32'd9565
; 
32'd187884: dataIn1 = 32'd9568
; 
32'd187885: dataIn1 = 32'd10037
; 
32'd187886: dataIn1 = 32'd10045
; 
32'd187887: dataIn1 = 32'd10049
; 
32'd187888: dataIn1 = 32'd9569
; 
32'd187889: dataIn1 = 32'd9570
; 
32'd187890: dataIn1 = 32'd9571
; 
32'd187891: dataIn1 = 32'd10050
; 
32'd187892: dataIn1 = 32'd10051
; 
32'd187893: dataIn1 = 32'd10052
; 
32'd187894: dataIn1 = 32'd3746
; 
32'd187895: dataIn1 = 32'd9571
; 
32'd187896: dataIn1 = 32'd10050
; 
32'd187897: dataIn1 = 32'd10051
; 
32'd187898: dataIn1 = 32'd10052
; 
32'd187899: dataIn1 = 32'd10058
; 
32'd187900: dataIn1 = 32'd10061
; 
32'd187901: dataIn1 = 32'd3746
; 
32'd187902: dataIn1 = 32'd9570
; 
32'd187903: dataIn1 = 32'd10050
; 
32'd187904: dataIn1 = 32'd10051
; 
32'd187905: dataIn1 = 32'd10052
; 
32'd187906: dataIn1 = 32'd10053
; 
32'd187907: dataIn1 = 32'd10056
; 
32'd187908: dataIn1 = 32'd9570
; 
32'd187909: dataIn1 = 32'd9572
; 
32'd187910: dataIn1 = 32'd10052
; 
32'd187911: dataIn1 = 32'd10053
; 
32'd187912: dataIn1 = 32'd10054
; 
32'd187913: dataIn1 = 32'd10055
; 
32'd187914: dataIn1 = 32'd10056
; 
32'd187915: dataIn1 = 32'd9561
; 
32'd187916: dataIn1 = 32'd9572
; 
32'd187917: dataIn1 = 32'd10040
; 
32'd187918: dataIn1 = 32'd10053
; 
32'd187919: dataIn1 = 32'd10054
; 
32'd187920: dataIn1 = 32'd10055
; 
32'd187921: dataIn1 = 32'd10057
; 
32'd187922: dataIn1 = 32'd3743
; 
32'd187923: dataIn1 = 32'd9561
; 
32'd187924: dataIn1 = 32'd9570
; 
32'd187925: dataIn1 = 32'd10053
; 
32'd187926: dataIn1 = 32'd10054
; 
32'd187927: dataIn1 = 32'd10055
; 
32'd187928: dataIn1 = 32'd3746
; 
32'd187929: dataIn1 = 32'd9572
; 
32'd187930: dataIn1 = 32'd10052
; 
32'd187931: dataIn1 = 32'd10053
; 
32'd187932: dataIn1 = 32'd10056
; 
32'd187933: dataIn1 = 32'd10203
; 
32'd187934: dataIn1 = 32'd2217
; 
32'd187935: dataIn1 = 32'd9572
; 
32'd187936: dataIn1 = 32'd10040
; 
32'd187937: dataIn1 = 32'd10054
; 
32'd187938: dataIn1 = 32'd10057
; 
32'd187939: dataIn1 = 32'd10204
; 
32'd187940: dataIn1 = 32'd9571
; 
32'd187941: dataIn1 = 32'd9574
; 
32'd187942: dataIn1 = 32'd10051
; 
32'd187943: dataIn1 = 32'd10058
; 
32'd187944: dataIn1 = 32'd10059
; 
32'd187945: dataIn1 = 32'd10060
; 
32'd187946: dataIn1 = 32'd10061
; 
32'd187947: dataIn1 = 32'd3747
; 
32'd187948: dataIn1 = 32'd9571
; 
32'd187949: dataIn1 = 32'd9573
; 
32'd187950: dataIn1 = 32'd10058
; 
32'd187951: dataIn1 = 32'd10059
; 
32'd187952: dataIn1 = 32'd10060
; 
32'd187953: dataIn1 = 32'd9573
; 
32'd187954: dataIn1 = 32'd9574
; 
32'd187955: dataIn1 = 32'd10058
; 
32'd187956: dataIn1 = 32'd10059
; 
32'd187957: dataIn1 = 32'd10060
; 
32'd187958: dataIn1 = 32'd10062
; 
32'd187959: dataIn1 = 32'd10063
; 
32'd187960: dataIn1 = 32'd3746
; 
32'd187961: dataIn1 = 32'd9574
; 
32'd187962: dataIn1 = 32'd10051
; 
32'd187963: dataIn1 = 32'd10058
; 
32'd187964: dataIn1 = 32'd10061
; 
32'd187965: dataIn1 = 32'd10206
; 
32'd187966: dataIn1 = 32'd67
; 
32'd187967: dataIn1 = 32'd9574
; 
32'd187968: dataIn1 = 32'd10060
; 
32'd187969: dataIn1 = 32'd10062
; 
32'd187970: dataIn1 = 32'd10063
; 
32'd187971: dataIn1 = 32'd10205
; 
32'd187972: dataIn1 = 32'd67
; 
32'd187973: dataIn1 = 32'd9573
; 
32'd187974: dataIn1 = 32'd10060
; 
32'd187975: dataIn1 = 32'd10062
; 
32'd187976: dataIn1 = 32'd10063
; 
32'd187977: dataIn1 = 32'd10064
; 
32'd187978: dataIn1 = 32'd10065
; 
32'd187979: dataIn1 = 32'd9573
; 
32'd187980: dataIn1 = 32'd9575
; 
32'd187981: dataIn1 = 32'd9576
; 
32'd187982: dataIn1 = 32'd10063
; 
32'd187983: dataIn1 = 32'd10064
; 
32'd187984: dataIn1 = 32'd10065
; 
32'd187985: dataIn1 = 32'd67
; 
32'd187986: dataIn1 = 32'd9576
; 
32'd187987: dataIn1 = 32'd10063
; 
32'd187988: dataIn1 = 32'd10064
; 
32'd187989: dataIn1 = 32'd10065
; 
32'd187990: dataIn1 = 32'd10072
; 
32'd187991: dataIn1 = 32'd10075
; 
32'd187992: dataIn1 = 32'd2220
; 
32'd187993: dataIn1 = 32'd9579
; 
32'd187994: dataIn1 = 32'd10066
; 
32'd187995: dataIn1 = 32'd10067
; 
32'd187996: dataIn1 = 32'd10068
; 
32'd187997: dataIn1 = 32'd10078
; 
32'd187998: dataIn1 = 32'd10080
; 
32'd187999: dataIn1 = 32'd9577
; 
32'd188000: dataIn1 = 32'd9578
; 
32'd188001: dataIn1 = 32'd9579
; 
32'd188002: dataIn1 = 32'd10066
; 
32'd188003: dataIn1 = 32'd10067
; 
32'd188004: dataIn1 = 32'd10068
; 
32'd188005: dataIn1 = 32'd2220
; 
32'd188006: dataIn1 = 32'd9577
; 
32'd188007: dataIn1 = 32'd10066
; 
32'd188008: dataIn1 = 32'd10067
; 
32'd188009: dataIn1 = 32'd10068
; 
32'd188010: dataIn1 = 32'd10086
; 
32'd188011: dataIn1 = 32'd10089
; 
32'd188012: dataIn1 = 32'd3758
; 
32'd188013: dataIn1 = 32'd9581
; 
32'd188014: dataIn1 = 32'd10069
; 
32'd188015: dataIn1 = 32'd10070
; 
32'd188016: dataIn1 = 32'd10071
; 
32'd188017: dataIn1 = 32'd10079
; 
32'd188018: dataIn1 = 32'd10081
; 
32'd188019: dataIn1 = 32'd3758
; 
32'd188020: dataIn1 = 32'd9580
; 
32'd188021: dataIn1 = 32'd10069
; 
32'd188022: dataIn1 = 32'd10070
; 
32'd188023: dataIn1 = 32'd10071
; 
32'd188024: dataIn1 = 32'd10074
; 
32'd188025: dataIn1 = 32'd10076
; 
32'd188026: dataIn1 = 32'd9580
; 
32'd188027: dataIn1 = 32'd9581
; 
32'd188028: dataIn1 = 32'd9582
; 
32'd188029: dataIn1 = 32'd10069
; 
32'd188030: dataIn1 = 32'd10070
; 
32'd188031: dataIn1 = 32'd10071
; 
32'd188032: dataIn1 = 32'd9576
; 
32'd188033: dataIn1 = 32'd9583
; 
32'd188034: dataIn1 = 32'd10065
; 
32'd188035: dataIn1 = 32'd10072
; 
32'd188036: dataIn1 = 32'd10073
; 
32'd188037: dataIn1 = 32'd10074
; 
32'd188038: dataIn1 = 32'd10075
; 
32'd188039: dataIn1 = 32'd3751
; 
32'd188040: dataIn1 = 32'd9576
; 
32'd188041: dataIn1 = 32'd9580
; 
32'd188042: dataIn1 = 32'd10072
; 
32'd188043: dataIn1 = 32'd10073
; 
32'd188044: dataIn1 = 32'd10074
; 
32'd188045: dataIn1 = 32'd9580
; 
32'd188046: dataIn1 = 32'd9583
; 
32'd188047: dataIn1 = 32'd10070
; 
32'd188048: dataIn1 = 32'd10072
; 
32'd188049: dataIn1 = 32'd10073
; 
32'd188050: dataIn1 = 32'd10074
; 
32'd188051: dataIn1 = 32'd10076
; 
32'd188052: dataIn1 = 32'd67
; 
32'd188053: dataIn1 = 32'd9583
; 
32'd188054: dataIn1 = 32'd10065
; 
32'd188055: dataIn1 = 32'd10072
; 
32'd188056: dataIn1 = 32'd10075
; 
32'd188057: dataIn1 = 32'd10208
; 
32'd188058: dataIn1 = 32'd3758
; 
32'd188059: dataIn1 = 32'd9583
; 
32'd188060: dataIn1 = 32'd10070
; 
32'd188061: dataIn1 = 32'd10074
; 
32'd188062: dataIn1 = 32'd10076
; 
32'd188063: dataIn1 = 32'd10207
; 
32'd188064: dataIn1 = 32'd3755
; 
32'd188065: dataIn1 = 32'd9579
; 
32'd188066: dataIn1 = 32'd9581
; 
32'd188067: dataIn1 = 32'd10077
; 
32'd188068: dataIn1 = 32'd10078
; 
32'd188069: dataIn1 = 32'd10079
; 
32'd188070: dataIn1 = 32'd9579
; 
32'd188071: dataIn1 = 32'd9584
; 
32'd188072: dataIn1 = 32'd10066
; 
32'd188073: dataIn1 = 32'd10077
; 
32'd188074: dataIn1 = 32'd10078
; 
32'd188075: dataIn1 = 32'd10079
; 
32'd188076: dataIn1 = 32'd10080
; 
32'd188077: dataIn1 = 32'd9581
; 
32'd188078: dataIn1 = 32'd9584
; 
32'd188079: dataIn1 = 32'd10069
; 
32'd188080: dataIn1 = 32'd10077
; 
32'd188081: dataIn1 = 32'd10078
; 
32'd188082: dataIn1 = 32'd10079
; 
32'd188083: dataIn1 = 32'd10081
; 
32'd188084: dataIn1 = 32'd2220
; 
32'd188085: dataIn1 = 32'd9584
; 
32'd188086: dataIn1 = 32'd10066
; 
32'd188087: dataIn1 = 32'd10078
; 
32'd188088: dataIn1 = 32'd10080
; 
32'd188089: dataIn1 = 32'd10210
; 
32'd188090: dataIn1 = 32'd3758
; 
32'd188091: dataIn1 = 32'd9584
; 
32'd188092: dataIn1 = 32'd10069
; 
32'd188093: dataIn1 = 32'd10079
; 
32'd188094: dataIn1 = 32'd10081
; 
32'd188095: dataIn1 = 32'd10209
; 
32'd188096: dataIn1 = 32'd9585
; 
32'd188097: dataIn1 = 32'd9586
; 
32'd188098: dataIn1 = 32'd9587
; 
32'd188099: dataIn1 = 32'd10082
; 
32'd188100: dataIn1 = 32'd10083
; 
32'd188101: dataIn1 = 32'd10084
; 
32'd188102: dataIn1 = 32'd3660
; 
32'd188103: dataIn1 = 32'd9587
; 
32'd188104: dataIn1 = 32'd10082
; 
32'd188105: dataIn1 = 32'd10083
; 
32'd188106: dataIn1 = 32'd10084
; 
32'd188107: dataIn1 = 32'd10090
; 
32'd188108: dataIn1 = 32'd10093
; 
32'd188109: dataIn1 = 32'd3660
; 
32'd188110: dataIn1 = 32'd9586
; 
32'd188111: dataIn1 = 32'd10082
; 
32'd188112: dataIn1 = 32'd10083
; 
32'd188113: dataIn1 = 32'd10084
; 
32'd188114: dataIn1 = 32'd10085
; 
32'd188115: dataIn1 = 32'd10088
; 
32'd188116: dataIn1 = 32'd9586
; 
32'd188117: dataIn1 = 32'd9588
; 
32'd188118: dataIn1 = 32'd10084
; 
32'd188119: dataIn1 = 32'd10085
; 
32'd188120: dataIn1 = 32'd10086
; 
32'd188121: dataIn1 = 32'd10087
; 
32'd188122: dataIn1 = 32'd10088
; 
32'd188123: dataIn1 = 32'd9577
; 
32'd188124: dataIn1 = 32'd9588
; 
32'd188125: dataIn1 = 32'd10068
; 
32'd188126: dataIn1 = 32'd10085
; 
32'd188127: dataIn1 = 32'd10086
; 
32'd188128: dataIn1 = 32'd10087
; 
32'd188129: dataIn1 = 32'd10089
; 
32'd188130: dataIn1 = 32'd3757
; 
32'd188131: dataIn1 = 32'd9577
; 
32'd188132: dataIn1 = 32'd9586
; 
32'd188133: dataIn1 = 32'd10085
; 
32'd188134: dataIn1 = 32'd10086
; 
32'd188135: dataIn1 = 32'd10087
; 
32'd188136: dataIn1 = 32'd3660
; 
32'd188137: dataIn1 = 32'd9588
; 
32'd188138: dataIn1 = 32'd10084
; 
32'd188139: dataIn1 = 32'd10085
; 
32'd188140: dataIn1 = 32'd10088
; 
32'd188141: dataIn1 = 32'd10211
; 
32'd188142: dataIn1 = 32'd2220
; 
32'd188143: dataIn1 = 32'd9588
; 
32'd188144: dataIn1 = 32'd10068
; 
32'd188145: dataIn1 = 32'd10086
; 
32'd188146: dataIn1 = 32'd10089
; 
32'd188147: dataIn1 = 32'd10212
; 
32'd188148: dataIn1 = 32'd9587
; 
32'd188149: dataIn1 = 32'd9590
; 
32'd188150: dataIn1 = 32'd10083
; 
32'd188151: dataIn1 = 32'd10090
; 
32'd188152: dataIn1 = 32'd10091
; 
32'd188153: dataIn1 = 32'd10092
; 
32'd188154: dataIn1 = 32'd10093
; 
32'd188155: dataIn1 = 32'd3760
; 
32'd188156: dataIn1 = 32'd9587
; 
32'd188157: dataIn1 = 32'd9589
; 
32'd188158: dataIn1 = 32'd10090
; 
32'd188159: dataIn1 = 32'd10091
; 
32'd188160: dataIn1 = 32'd10092
; 
32'd188161: dataIn1 = 32'd9589
; 
32'd188162: dataIn1 = 32'd9590
; 
32'd188163: dataIn1 = 32'd10090
; 
32'd188164: dataIn1 = 32'd10091
; 
32'd188165: dataIn1 = 32'd10092
; 
32'd188166: dataIn1 = 32'd10094
; 
32'd188167: dataIn1 = 32'd10095
; 
32'd188168: dataIn1 = 32'd3660
; 
32'd188169: dataIn1 = 32'd9590
; 
32'd188170: dataIn1 = 32'd10083
; 
32'd188171: dataIn1 = 32'd10090
; 
32'd188172: dataIn1 = 32'd10093
; 
32'd188173: dataIn1 = 32'd10214
; 
32'd188174: dataIn1 = 32'd68
; 
32'd188175: dataIn1 = 32'd9590
; 
32'd188176: dataIn1 = 32'd10092
; 
32'd188177: dataIn1 = 32'd10094
; 
32'd188178: dataIn1 = 32'd10095
; 
32'd188179: dataIn1 = 32'd10213
; 
32'd188180: dataIn1 = 32'd68
; 
32'd188181: dataIn1 = 32'd9589
; 
32'd188182: dataIn1 = 32'd10092
; 
32'd188183: dataIn1 = 32'd10094
; 
32'd188184: dataIn1 = 32'd10095
; 
32'd188185: dataIn1 = 32'd10096
; 
32'd188186: dataIn1 = 32'd10097
; 
32'd188187: dataIn1 = 32'd9589
; 
32'd188188: dataIn1 = 32'd9591
; 
32'd188189: dataIn1 = 32'd9592
; 
32'd188190: dataIn1 = 32'd10095
; 
32'd188191: dataIn1 = 32'd10096
; 
32'd188192: dataIn1 = 32'd10097
; 
32'd188193: dataIn1 = 32'd68
; 
32'd188194: dataIn1 = 32'd9592
; 
32'd188195: dataIn1 = 32'd10095
; 
32'd188196: dataIn1 = 32'd10096
; 
32'd188197: dataIn1 = 32'd10097
; 
32'd188198: dataIn1 = 32'd10104
; 
32'd188199: dataIn1 = 32'd10107
; 
32'd188200: dataIn1 = 32'd2223
; 
32'd188201: dataIn1 = 32'd9595
; 
32'd188202: dataIn1 = 32'd10098
; 
32'd188203: dataIn1 = 32'd10099
; 
32'd188204: dataIn1 = 32'd10100
; 
32'd188205: dataIn1 = 32'd10110
; 
32'd188206: dataIn1 = 32'd10112
; 
32'd188207: dataIn1 = 32'd9593
; 
32'd188208: dataIn1 = 32'd9594
; 
32'd188209: dataIn1 = 32'd9595
; 
32'd188210: dataIn1 = 32'd10098
; 
32'd188211: dataIn1 = 32'd10099
; 
32'd188212: dataIn1 = 32'd10100
; 
32'd188213: dataIn1 = 32'd2223
; 
32'd188214: dataIn1 = 32'd9593
; 
32'd188215: dataIn1 = 32'd10098
; 
32'd188216: dataIn1 = 32'd10099
; 
32'd188217: dataIn1 = 32'd10100
; 
32'd188218: dataIn1 = 32'd10115
; 
32'd188219: dataIn1 = 32'd10118
; 
32'd188220: dataIn1 = 32'd3667
; 
32'd188221: dataIn1 = 32'd9597
; 
32'd188222: dataIn1 = 32'd10101
; 
32'd188223: dataIn1 = 32'd10102
; 
32'd188224: dataIn1 = 32'd10103
; 
32'd188225: dataIn1 = 32'd10111
; 
32'd188226: dataIn1 = 32'd10113
; 
32'd188227: dataIn1 = 32'd3667
; 
32'd188228: dataIn1 = 32'd9596
; 
32'd188229: dataIn1 = 32'd10101
; 
32'd188230: dataIn1 = 32'd10102
; 
32'd188231: dataIn1 = 32'd10103
; 
32'd188232: dataIn1 = 32'd10106
; 
32'd188233: dataIn1 = 32'd10108
; 
32'd188234: dataIn1 = 32'd9596
; 
32'd188235: dataIn1 = 32'd9597
; 
32'd188236: dataIn1 = 32'd9598
; 
32'd188237: dataIn1 = 32'd10101
; 
32'd188238: dataIn1 = 32'd10102
; 
32'd188239: dataIn1 = 32'd10103
; 
32'd188240: dataIn1 = 32'd9592
; 
32'd188241: dataIn1 = 32'd9599
; 
32'd188242: dataIn1 = 32'd10097
; 
32'd188243: dataIn1 = 32'd10104
; 
32'd188244: dataIn1 = 32'd10105
; 
32'd188245: dataIn1 = 32'd10106
; 
32'd188246: dataIn1 = 32'd10107
; 
32'd188247: dataIn1 = 32'd3764
; 
32'd188248: dataIn1 = 32'd9592
; 
32'd188249: dataIn1 = 32'd9596
; 
32'd188250: dataIn1 = 32'd10104
; 
32'd188251: dataIn1 = 32'd10105
; 
32'd188252: dataIn1 = 32'd10106
; 
32'd188253: dataIn1 = 32'd9596
; 
32'd188254: dataIn1 = 32'd9599
; 
32'd188255: dataIn1 = 32'd10102
; 
32'd188256: dataIn1 = 32'd10104
; 
32'd188257: dataIn1 = 32'd10105
; 
32'd188258: dataIn1 = 32'd10106
; 
32'd188259: dataIn1 = 32'd10108
; 
32'd188260: dataIn1 = 32'd68
; 
32'd188261: dataIn1 = 32'd9599
; 
32'd188262: dataIn1 = 32'd10097
; 
32'd188263: dataIn1 = 32'd10104
; 
32'd188264: dataIn1 = 32'd10107
; 
32'd188265: dataIn1 = 32'd10216
; 
32'd188266: dataIn1 = 32'd3667
; 
32'd188267: dataIn1 = 32'd9599
; 
32'd188268: dataIn1 = 32'd10102
; 
32'd188269: dataIn1 = 32'd10106
; 
32'd188270: dataIn1 = 32'd10108
; 
32'd188271: dataIn1 = 32'd10215
; 
32'd188272: dataIn1 = 32'd3768
; 
32'd188273: dataIn1 = 32'd9595
; 
32'd188274: dataIn1 = 32'd9597
; 
32'd188275: dataIn1 = 32'd10109
; 
32'd188276: dataIn1 = 32'd10110
; 
32'd188277: dataIn1 = 32'd10111
; 
32'd188278: dataIn1 = 32'd9595
; 
32'd188279: dataIn1 = 32'd9600
; 
32'd188280: dataIn1 = 32'd10098
; 
32'd188281: dataIn1 = 32'd10109
; 
32'd188282: dataIn1 = 32'd10110
; 
32'd188283: dataIn1 = 32'd10111
; 
32'd188284: dataIn1 = 32'd10112
; 
32'd188285: dataIn1 = 32'd9597
; 
32'd188286: dataIn1 = 32'd9600
; 
32'd188287: dataIn1 = 32'd10101
; 
32'd188288: dataIn1 = 32'd10109
; 
32'd188289: dataIn1 = 32'd10110
; 
32'd188290: dataIn1 = 32'd10111
; 
32'd188291: dataIn1 = 32'd10113
; 
32'd188292: dataIn1 = 32'd2223
; 
32'd188293: dataIn1 = 32'd9600
; 
32'd188294: dataIn1 = 32'd10098
; 
32'd188295: dataIn1 = 32'd10110
; 
32'd188296: dataIn1 = 32'd10112
; 
32'd188297: dataIn1 = 32'd10218
; 
32'd188298: dataIn1 = 32'd3667
; 
32'd188299: dataIn1 = 32'd9600
; 
32'd188300: dataIn1 = 32'd10101
; 
32'd188301: dataIn1 = 32'd10111
; 
32'd188302: dataIn1 = 32'd10113
; 
32'd188303: dataIn1 = 32'd10217
; 
32'd188304: dataIn1 = 32'd9502
; 
32'd188305: dataIn1 = 32'd9601
; 
32'd188306: dataIn1 = 32'd9914
; 
32'd188307: dataIn1 = 32'd10114
; 
32'd188308: dataIn1 = 32'd10115
; 
32'd188309: dataIn1 = 32'd10116
; 
32'd188310: dataIn1 = 32'd10117
; 
32'd188311: dataIn1 = 32'd9502
; 
32'd188312: dataIn1 = 32'd9593
; 
32'd188313: dataIn1 = 32'd10100
; 
32'd188314: dataIn1 = 32'd10114
; 
32'd188315: dataIn1 = 32'd10115
; 
32'd188316: dataIn1 = 32'd10116
; 
32'd188317: dataIn1 = 32'd10118
; 
32'd188318: dataIn1 = 32'd3770
; 
32'd188319: dataIn1 = 32'd9593
; 
32'd188320: dataIn1 = 32'd9601
; 
32'd188321: dataIn1 = 32'd10114
; 
32'd188322: dataIn1 = 32'd10115
; 
32'd188323: dataIn1 = 32'd10116
; 
32'd188324: dataIn1 = 32'd3669
; 
32'd188325: dataIn1 = 32'd9601
; 
32'd188326: dataIn1 = 32'd9914
; 
32'd188327: dataIn1 = 32'd10114
; 
32'd188328: dataIn1 = 32'd10117
; 
32'd188329: dataIn1 = 32'd10174
; 
32'd188330: dataIn1 = 32'd2223
; 
32'd188331: dataIn1 = 32'd9501
; 
32'd188332: dataIn1 = 32'd9502
; 
32'd188333: dataIn1 = 32'd10100
; 
32'd188334: dataIn1 = 32'd10115
; 
32'd188335: dataIn1 = 32'd10118
; 
32'd188336: dataIn1 = 32'd6162
; 
32'd188337: dataIn1 = 32'd9669
; 
32'd188338: dataIn1 = 32'd10119
; 
32'd188339: dataIn1 = 32'd10120
; 
32'd188340: dataIn1 = 32'd10121
; 
32'd188341: dataIn1 = 32'd10122
; 
32'd188342: dataIn1 = 32'd10123
; 
32'd188343: dataIn1 = 32'd2700
; 
32'd188344: dataIn1 = 32'd9669
; 
32'd188345: dataIn1 = 32'd9670
; 
32'd188346: dataIn1 = 32'd10119
; 
32'd188347: dataIn1 = 32'd10120
; 
32'd188348: dataIn1 = 32'd10121
; 
32'd188349: dataIn1 = 32'd6162
; 
32'd188350: dataIn1 = 32'd9670
; 
32'd188351: dataIn1 = 32'd10119
; 
32'd188352: dataIn1 = 32'd10120
; 
32'd188353: dataIn1 = 32'd10121
; 
32'd188354: dataIn1 = 32'd10124
; 
32'd188355: dataIn1 = 32'd10125
; 
32'd188356: dataIn1 = 32'd5140
; 
32'd188357: dataIn1 = 32'd9669
; 
32'd188358: dataIn1 = 32'd9760
; 
32'd188359: dataIn1 = 32'd10119
; 
32'd188360: dataIn1 = 32'd10122
; 
32'd188361: dataIn1 = 32'd10123
; 
32'd188362: dataIn1 = 32'd10150
; 
32'd188363: dataIn1 = 32'd5140
; 
32'd188364: dataIn1 = 32'd6162
; 
32'd188365: dataIn1 = 32'd7262
; 
32'd188366: dataIn1 = 32'd10119
; 
32'd188367: dataIn1 = 32'd10122
; 
32'd188368: dataIn1 = 32'd10123
; 
32'd188369: dataIn1 = 32'd10220
; 
32'd188370: dataIn1 = 32'd5143
; 
32'd188371: dataIn1 = 32'd6162
; 
32'd188372: dataIn1 = 32'd9778
; 
32'd188373: dataIn1 = 32'd10121
; 
32'd188374: dataIn1 = 32'd10124
; 
32'd188375: dataIn1 = 32'd10125
; 
32'd188376: dataIn1 = 32'd10151
; 
32'd188377: dataIn1 = 32'd5143
; 
32'd188378: dataIn1 = 32'd9670
; 
32'd188379: dataIn1 = 32'd9745
; 
32'd188380: dataIn1 = 32'd10121
; 
32'd188381: dataIn1 = 32'd10124
; 
32'd188382: dataIn1 = 32'd10125
; 
32'd188383: dataIn1 = 32'd10134
; 
32'd188384: dataIn1 = 32'd6738
; 
32'd188385: dataIn1 = 32'd9672
; 
32'd188386: dataIn1 = 32'd9673
; 
32'd188387: dataIn1 = 32'd9754
; 
32'd188388: dataIn1 = 32'd10126
; 
32'd188389: dataIn1 = 32'd10127
; 
32'd188390: dataIn1 = 32'd5440
; 
32'd188391: dataIn1 = 32'd9673
; 
32'd188392: dataIn1 = 32'd9754
; 
32'd188393: dataIn1 = 32'd10126
; 
32'd188394: dataIn1 = 32'd10127
; 
32'd188395: dataIn1 = 32'd10128
; 
32'd188396: dataIn1 = 32'd10131
; 
32'd188397: dataIn1 = 32'd10148
; 
32'd188398: dataIn1 = 32'd9673
; 
32'd188399: dataIn1 = 32'd9675
; 
32'd188400: dataIn1 = 32'd10127
; 
32'd188401: dataIn1 = 32'd10128
; 
32'd188402: dataIn1 = 32'd10129
; 
32'd188403: dataIn1 = 32'd10130
; 
32'd188404: dataIn1 = 32'd10131
; 
32'd188405: dataIn1 = 32'd20
; 
32'd188406: dataIn1 = 32'd9674
; 
32'd188407: dataIn1 = 32'd9675
; 
32'd188408: dataIn1 = 32'd10128
; 
32'd188409: dataIn1 = 32'd10129
; 
32'd188410: dataIn1 = 32'd10130
; 
32'd188411: dataIn1 = 32'd9673
; 
32'd188412: dataIn1 = 32'd9674
; 
32'd188413: dataIn1 = 32'd10128
; 
32'd188414: dataIn1 = 32'd10129
; 
32'd188415: dataIn1 = 32'd10130
; 
32'd188416: dataIn1 = 32'd10132
; 
32'd188417: dataIn1 = 32'd10133
; 
32'd188418: dataIn1 = 32'd5440
; 
32'd188419: dataIn1 = 32'd6739
; 
32'd188420: dataIn1 = 32'd9675
; 
32'd188421: dataIn1 = 32'd10127
; 
32'd188422: dataIn1 = 32'd10128
; 
32'd188423: dataIn1 = 32'd10131
; 
32'd188424: dataIn1 = 32'd5520
; 
32'd188425: dataIn1 = 32'd9672
; 
32'd188426: dataIn1 = 32'd9673
; 
32'd188427: dataIn1 = 32'd10130
; 
32'd188428: dataIn1 = 32'd10132
; 
32'd188429: dataIn1 = 32'd10133
; 
32'd188430: dataIn1 = 32'd5520
; 
32'd188431: dataIn1 = 32'd9674
; 
32'd188432: dataIn1 = 32'd9822
; 
32'd188433: dataIn1 = 32'd10130
; 
32'd188434: dataIn1 = 32'd10132
; 
32'd188435: dataIn1 = 32'd10133
; 
32'd188436: dataIn1 = 32'd6597
; 
32'd188437: dataIn1 = 32'd9670
; 
32'd188438: dataIn1 = 32'd9671
; 
32'd188439: dataIn1 = 32'd9745
; 
32'd188440: dataIn1 = 32'd10125
; 
32'd188441: dataIn1 = 32'd10134
; 
32'd188442: dataIn1 = 32'd6713
; 
32'd188443: dataIn1 = 32'd9749
; 
32'd188444: dataIn1 = 32'd10135
; 
32'd188445: dataIn1 = 32'd10136
; 
32'd188446: dataIn1 = 32'd10137
; 
32'd188447: dataIn1 = 32'd10142
; 
32'd188448: dataIn1 = 32'd10143
; 
32'd188449: dataIn1 = 32'd9747
; 
32'd188450: dataIn1 = 32'd9748
; 
32'd188451: dataIn1 = 32'd9749
; 
32'd188452: dataIn1 = 32'd10135
; 
32'd188453: dataIn1 = 32'd10136
; 
32'd188454: dataIn1 = 32'd10137
; 
32'd188455: dataIn1 = 32'd6713
; 
32'd188456: dataIn1 = 32'd9747
; 
32'd188457: dataIn1 = 32'd10135
; 
32'd188458: dataIn1 = 32'd10136
; 
32'd188459: dataIn1 = 32'd10137
; 
32'd188460: dataIn1 = 32'd10139
; 
32'd188461: dataIn1 = 32'd10141
; 
32'd188462: dataIn1 = 32'd1129
; 
32'd188463: dataIn1 = 32'd6395
; 
32'd188464: dataIn1 = 32'd9750
; 
32'd188465: dataIn1 = 32'd10138
; 
32'd188466: dataIn1 = 32'd10139
; 
32'd188467: dataIn1 = 32'd10140
; 
32'd188468: dataIn1 = 32'd9747
; 
32'd188469: dataIn1 = 32'd9750
; 
32'd188470: dataIn1 = 32'd10137
; 
32'd188471: dataIn1 = 32'd10138
; 
32'd188472: dataIn1 = 32'd10139
; 
32'd188473: dataIn1 = 32'd10140
; 
32'd188474: dataIn1 = 32'd10141
; 
32'd188475: dataIn1 = 32'd6395
; 
32'd188476: dataIn1 = 32'd9740
; 
32'd188477: dataIn1 = 32'd9747
; 
32'd188478: dataIn1 = 32'd10138
; 
32'd188479: dataIn1 = 32'd10139
; 
32'd188480: dataIn1 = 32'd10140
; 
32'd188481: dataIn1 = 32'd10221
; 
32'd188482: dataIn1 = 32'd6713
; 
32'd188483: dataIn1 = 32'd9750
; 
32'd188484: dataIn1 = 32'd10137
; 
32'd188485: dataIn1 = 32'd10139
; 
32'd188486: dataIn1 = 32'd10141
; 
32'd188487: dataIn1 = 32'd10223
; 
32'd188488: dataIn1 = 32'd9749
; 
32'd188489: dataIn1 = 32'd9751
; 
32'd188490: dataIn1 = 32'd9752
; 
32'd188491: dataIn1 = 32'd10135
; 
32'd188492: dataIn1 = 32'd10142
; 
32'd188493: dataIn1 = 32'd10143
; 
32'd188494: dataIn1 = 32'd6713
; 
32'd188495: dataIn1 = 32'd9751
; 
32'd188496: dataIn1 = 32'd10135
; 
32'd188497: dataIn1 = 32'd10142
; 
32'd188498: dataIn1 = 32'd10143
; 
32'd188499: dataIn1 = 32'd10145
; 
32'd188500: dataIn1 = 32'd10149
; 
32'd188501: dataIn1 = 32'd9751
; 
32'd188502: dataIn1 = 32'd9754
; 
32'd188503: dataIn1 = 32'd10144
; 
32'd188504: dataIn1 = 32'd10145
; 
32'd188505: dataIn1 = 32'd10146
; 
32'd188506: dataIn1 = 32'd10147
; 
32'd188507: dataIn1 = 32'd10148
; 
32'd188508: dataIn1 = 32'd9751
; 
32'd188509: dataIn1 = 32'd9753
; 
32'd188510: dataIn1 = 32'd10143
; 
32'd188511: dataIn1 = 32'd10144
; 
32'd188512: dataIn1 = 32'd10145
; 
32'd188513: dataIn1 = 32'd10146
; 
32'd188514: dataIn1 = 32'd10149
; 
32'd188515: dataIn1 = 32'd6738
; 
32'd188516: dataIn1 = 32'd9753
; 
32'd188517: dataIn1 = 32'd9754
; 
32'd188518: dataIn1 = 32'd10144
; 
32'd188519: dataIn1 = 32'd10145
; 
32'd188520: dataIn1 = 32'd10146
; 
32'd188521: dataIn1 = 32'd5440
; 
32'd188522: dataIn1 = 32'd9751
; 
32'd188523: dataIn1 = 32'd9752
; 
32'd188524: dataIn1 = 32'd10144
; 
32'd188525: dataIn1 = 32'd10147
; 
32'd188526: dataIn1 = 32'd10148
; 
32'd188527: dataIn1 = 32'd5440
; 
32'd188528: dataIn1 = 32'd9754
; 
32'd188529: dataIn1 = 32'd10127
; 
32'd188530: dataIn1 = 32'd10144
; 
32'd188531: dataIn1 = 32'd10147
; 
32'd188532: dataIn1 = 32'd10148
; 
32'd188533: dataIn1 = 32'd6713
; 
32'd188534: dataIn1 = 32'd9753
; 
32'd188535: dataIn1 = 32'd10143
; 
32'd188536: dataIn1 = 32'd10145
; 
32'd188537: dataIn1 = 32'd10149
; 
32'd188538: dataIn1 = 32'd10223
; 
32'd188539: dataIn1 = 32'd6155
; 
32'd188540: dataIn1 = 32'd9668
; 
32'd188541: dataIn1 = 32'd9669
; 
32'd188542: dataIn1 = 32'd9760
; 
32'd188543: dataIn1 = 32'd10122
; 
32'd188544: dataIn1 = 32'd10150
; 
32'd188545: dataIn1 = 32'd6161
; 
32'd188546: dataIn1 = 32'd6162
; 
32'd188547: dataIn1 = 32'd9286
; 
32'd188548: dataIn1 = 32'd9778
; 
32'd188549: dataIn1 = 32'd10124
; 
32'd188550: dataIn1 = 32'd10151
; 
32'd188551: dataIn1 = 32'd10220
; 
32'd188552: dataIn1 = 32'd2114
; 
32'd188553: dataIn1 = 32'd2115
; 
32'd188554: dataIn1 = 32'd9454
; 
32'd188555: dataIn1 = 32'd9456
; 
32'd188556: dataIn1 = 32'd9821
; 
32'd188557: dataIn1 = 32'd9826
; 
32'd188558: dataIn1 = 32'd10152
; 
32'd188559: dataIn1 = 32'd10153
; 
32'd188560: dataIn1 = 32'd10154
; 
32'd188561: dataIn1 = 32'd31
; 
32'd188562: dataIn1 = 32'd2115
; 
32'd188563: dataIn1 = 32'd2116
; 
32'd188564: dataIn1 = 32'd9454
; 
32'd188565: dataIn1 = 32'd10152
; 
32'd188566: dataIn1 = 32'd10153
; 
32'd188567: dataIn1 = 32'd1141
; 
32'd188568: dataIn1 = 32'd2115
; 
32'd188569: dataIn1 = 32'd5523
; 
32'd188570: dataIn1 = 32'd9456
; 
32'd188571: dataIn1 = 32'd10152
; 
32'd188572: dataIn1 = 32'd10154
; 
32'd188573: dataIn1 = 32'd10225
; 
32'd188574: dataIn1 = 32'd10283
; 
32'd188575: dataIn1 = 32'd30
; 
32'd188576: dataIn1 = 32'd2113
; 
32'd188577: dataIn1 = 32'd2146
; 
32'd188578: dataIn1 = 32'd9458
; 
32'd188579: dataIn1 = 32'd9832
; 
32'd188580: dataIn1 = 32'd10155
; 
32'd188581: dataIn1 = 32'd10156
; 
32'd188582: dataIn1 = 32'd2146
; 
32'd188583: dataIn1 = 32'd2147
; 
32'd188584: dataIn1 = 32'd9458
; 
32'd188585: dataIn1 = 32'd9463
; 
32'd188586: dataIn1 = 32'd9830
; 
32'd188587: dataIn1 = 32'd9842
; 
32'd188588: dataIn1 = 32'd10155
; 
32'd188589: dataIn1 = 32'd10156
; 
32'd188590: dataIn1 = 32'd10157
; 
32'd188591: dataIn1 = 32'd41
; 
32'd188592: dataIn1 = 32'd2145
; 
32'd188593: dataIn1 = 32'd2146
; 
32'd188594: dataIn1 = 32'd9463
; 
32'd188595: dataIn1 = 32'd10156
; 
32'd188596: dataIn1 = 32'd10157
; 
32'd188597: dataIn1 = 32'd52
; 
32'd188598: dataIn1 = 32'd3588
; 
32'd188599: dataIn1 = 32'd9470
; 
32'd188600: dataIn1 = 32'd9853
; 
32'd188601: dataIn1 = 32'd10158
; 
32'd188602: dataIn1 = 32'd10159
; 
32'd188603: dataIn1 = 32'd10172
; 
32'd188604: dataIn1 = 32'd10226
; 
32'd188605: dataIn1 = 32'd52
; 
32'd188606: dataIn1 = 32'd3587
; 
32'd188607: dataIn1 = 32'd3591
; 
32'd188608: dataIn1 = 32'd9470
; 
32'd188609: dataIn1 = 32'd10158
; 
32'd188610: dataIn1 = 32'd10159
; 
32'd188611: dataIn1 = 32'd3589
; 
32'd188612: dataIn1 = 32'd9473
; 
32'd188613: dataIn1 = 32'd9770
; 
32'd188614: dataIn1 = 32'd9771
; 
32'd188615: dataIn1 = 32'd9864
; 
32'd188616: dataIn1 = 32'd10160
; 
32'd188617: dataIn1 = 32'd10161
; 
32'd188618: dataIn1 = 32'd2177
; 
32'd188619: dataIn1 = 32'd9473
; 
32'd188620: dataIn1 = 32'd9770
; 
32'd188621: dataIn1 = 32'd9849
; 
32'd188622: dataIn1 = 32'd9863
; 
32'd188623: dataIn1 = 32'd10160
; 
32'd188624: dataIn1 = 32'd10161
; 
32'd188625: dataIn1 = 32'd10227
; 
32'd188626: dataIn1 = 32'd3622
; 
32'd188627: dataIn1 = 32'd3627
; 
32'd188628: dataIn1 = 32'd9481
; 
32'd188629: dataIn1 = 32'd9487
; 
32'd188630: dataIn1 = 32'd9875
; 
32'd188631: dataIn1 = 32'd9889
; 
32'd188632: dataIn1 = 32'd10162
; 
32'd188633: dataIn1 = 32'd10163
; 
32'd188634: dataIn1 = 32'd10166
; 
32'd188635: dataIn1 = 32'd2204
; 
32'd188636: dataIn1 = 32'd3627
; 
32'd188637: dataIn1 = 32'd3708
; 
32'd188638: dataIn1 = 32'd9481
; 
32'd188639: dataIn1 = 32'd10162
; 
32'd188640: dataIn1 = 32'd10163
; 
32'd188641: dataIn1 = 32'd3619
; 
32'd188642: dataIn1 = 32'd3625
; 
32'd188643: dataIn1 = 32'd9485
; 
32'd188644: dataIn1 = 32'd9556
; 
32'd188645: dataIn1 = 32'd9883
; 
32'd188646: dataIn1 = 32'd10025
; 
32'd188647: dataIn1 = 32'd10164
; 
32'd188648: dataIn1 = 32'd10165
; 
32'd188649: dataIn1 = 32'd10196
; 
32'd188650: dataIn1 = 32'd2203
; 
32'd188651: dataIn1 = 32'd3619
; 
32'd188652: dataIn1 = 32'd3621
; 
32'd188653: dataIn1 = 32'd9485
; 
32'd188654: dataIn1 = 32'd9881
; 
32'd188655: dataIn1 = 32'd10164
; 
32'd188656: dataIn1 = 32'd10165
; 
32'd188657: dataIn1 = 32'd62
; 
32'd188658: dataIn1 = 32'd3626
; 
32'd188659: dataIn1 = 32'd3627
; 
32'd188660: dataIn1 = 32'd9487
; 
32'd188661: dataIn1 = 32'd10162
; 
32'd188662: dataIn1 = 32'd10166
; 
32'd188663: dataIn1 = 32'd2206
; 
32'd188664: dataIn1 = 32'd3630
; 
32'd188665: dataIn1 = 32'd9489
; 
32'd188666: dataIn1 = 32'd9896
; 
32'd188667: dataIn1 = 32'd10167
; 
32'd188668: dataIn1 = 32'd10168
; 
32'd188669: dataIn1 = 32'd10171
; 
32'd188670: dataIn1 = 32'd10228
; 
32'd188671: dataIn1 = 32'd2206
; 
32'd188672: dataIn1 = 32'd3629
; 
32'd188673: dataIn1 = 32'd3632
; 
32'd188674: dataIn1 = 32'd9489
; 
32'd188675: dataIn1 = 32'd10167
; 
32'd188676: dataIn1 = 32'd10168
; 
32'd188677: dataIn1 = 32'd2205
; 
32'd188678: dataIn1 = 32'd3624
; 
32'd188679: dataIn1 = 32'd9484
; 
32'd188680: dataIn1 = 32'd9495
; 
32'd188681: dataIn1 = 32'd9903
; 
32'd188682: dataIn1 = 32'd10169
; 
32'd188683: dataIn1 = 32'd10170
; 
32'd188684: dataIn1 = 32'd10229
; 
32'd188685: dataIn1 = 32'd3624
; 
32'd188686: dataIn1 = 32'd3628
; 
32'd188687: dataIn1 = 32'd3631
; 
32'd188688: dataIn1 = 32'd9495
; 
32'd188689: dataIn1 = 32'd9902
; 
32'd188690: dataIn1 = 32'd10169
; 
32'd188691: dataIn1 = 32'd10170
; 
32'd188692: dataIn1 = 32'd3630
; 
32'd188693: dataIn1 = 32'd3633
; 
32'd188694: dataIn1 = 32'd9497
; 
32'd188695: dataIn1 = 32'd9910
; 
32'd188696: dataIn1 = 32'd10167
; 
32'd188697: dataIn1 = 32'd10171
; 
32'd188698: dataIn1 = 32'd10172
; 
32'd188699: dataIn1 = 32'd10228
; 
32'd188700: dataIn1 = 32'd3588
; 
32'd188701: dataIn1 = 32'd3633
; 
32'd188702: dataIn1 = 32'd9497
; 
32'd188703: dataIn1 = 32'd9909
; 
32'd188704: dataIn1 = 32'd10158
; 
32'd188705: dataIn1 = 32'd10171
; 
32'd188706: dataIn1 = 32'd10172
; 
32'd188707: dataIn1 = 32'd10226
; 
32'd188708: dataIn1 = 32'd69
; 
32'd188709: dataIn1 = 32'd3772
; 
32'd188710: dataIn1 = 32'd9503
; 
32'd188711: dataIn1 = 32'd9921
; 
32'd188712: dataIn1 = 32'd10173
; 
32'd188713: dataIn1 = 32'd10174
; 
32'd188714: dataIn1 = 32'd10180
; 
32'd188715: dataIn1 = 32'd10230
; 
32'd188716: dataIn1 = 32'd3669
; 
32'd188717: dataIn1 = 32'd3772
; 
32'd188718: dataIn1 = 32'd9503
; 
32'd188719: dataIn1 = 32'd9601
; 
32'd188720: dataIn1 = 32'd9919
; 
32'd188721: dataIn1 = 32'd10117
; 
32'd188722: dataIn1 = 32'd10173
; 
32'd188723: dataIn1 = 32'd10174
; 
32'd188724: dataIn1 = 32'd10219
; 
32'd188725: dataIn1 = 32'd3672
; 
32'd188726: dataIn1 = 32'd3674
; 
32'd188727: dataIn1 = 32'd9507
; 
32'd188728: dataIn1 = 32'd9930
; 
32'd188729: dataIn1 = 32'd10175
; 
32'd188730: dataIn1 = 32'd10176
; 
32'd188731: dataIn1 = 32'd10181
; 
32'd188732: dataIn1 = 32'd10231
; 
32'd188733: dataIn1 = 32'd2225
; 
32'd188734: dataIn1 = 32'd3672
; 
32'd188735: dataIn1 = 32'd3673
; 
32'd188736: dataIn1 = 32'd9507
; 
32'd188737: dataIn1 = 32'd10175
; 
32'd188738: dataIn1 = 32'd10176
; 
32'd188739: dataIn1 = 32'd3677
; 
32'd188740: dataIn1 = 32'd3780
; 
32'd188741: dataIn1 = 32'd9513
; 
32'd188742: dataIn1 = 32'd9938
; 
32'd188743: dataIn1 = 32'd10177
; 
32'd188744: dataIn1 = 32'd10178
; 
32'd188745: dataIn1 = 32'd10179
; 
32'd188746: dataIn1 = 32'd10232
; 
32'd188747: dataIn1 = 32'd2226
; 
32'd188748: dataIn1 = 32'd3780
; 
32'd188749: dataIn1 = 32'd3782
; 
32'd188750: dataIn1 = 32'd9513
; 
32'd188751: dataIn1 = 32'd9937
; 
32'd188752: dataIn1 = 32'd10177
; 
32'd188753: dataIn1 = 32'd10178
; 
32'd188754: dataIn1 = 32'd3677
; 
32'd188755: dataIn1 = 32'd3776
; 
32'd188756: dataIn1 = 32'd9514
; 
32'd188757: dataIn1 = 32'd9943
; 
32'd188758: dataIn1 = 32'd10177
; 
32'd188759: dataIn1 = 32'd10179
; 
32'd188760: dataIn1 = 32'd10180
; 
32'd188761: dataIn1 = 32'd10232
; 
32'd188762: dataIn1 = 32'd69
; 
32'd188763: dataIn1 = 32'd3776
; 
32'd188764: dataIn1 = 32'd9514
; 
32'd188765: dataIn1 = 32'd9942
; 
32'd188766: dataIn1 = 32'd10173
; 
32'd188767: dataIn1 = 32'd10179
; 
32'd188768: dataIn1 = 32'd10180
; 
32'd188769: dataIn1 = 32'd10230
; 
32'd188770: dataIn1 = 32'd2227
; 
32'd188771: dataIn1 = 32'd3674
; 
32'd188772: dataIn1 = 32'd9516
; 
32'd188773: dataIn1 = 32'd9949
; 
32'd188774: dataIn1 = 32'd10175
; 
32'd188775: dataIn1 = 32'd10181
; 
32'd188776: dataIn1 = 32'd10182
; 
32'd188777: dataIn1 = 32'd10231
; 
32'd188778: dataIn1 = 32'd2227
; 
32'd188779: dataIn1 = 32'd3678
; 
32'd188780: dataIn1 = 32'd9516
; 
32'd188781: dataIn1 = 32'd9523
; 
32'd188782: dataIn1 = 32'd9948
; 
32'd188783: dataIn1 = 32'd10181
; 
32'd188784: dataIn1 = 32'd10182
; 
32'd188785: dataIn1 = 32'd10233
; 
32'd188786: dataIn1 = 32'd70
; 
32'd188787: dataIn1 = 32'd3691
; 
32'd188788: dataIn1 = 32'd3788
; 
32'd188789: dataIn1 = 32'd9526
; 
32'd188790: dataIn1 = 32'd10183
; 
32'd188791: dataIn1 = 32'd10184
; 
32'd188792: dataIn1 = 32'd3684
; 
32'd188793: dataIn1 = 32'd3691
; 
32'd188794: dataIn1 = 32'd9526
; 
32'd188795: dataIn1 = 32'd9534
; 
32'd188796: dataIn1 = 32'd9963
; 
32'd188797: dataIn1 = 32'd9982
; 
32'd188798: dataIn1 = 32'd10183
; 
32'd188799: dataIn1 = 32'd10184
; 
32'd188800: dataIn1 = 32'd10189
; 
32'd188801: dataIn1 = 32'd2229
; 
32'd188802: dataIn1 = 32'd3689
; 
32'd188803: dataIn1 = 32'd3693
; 
32'd188804: dataIn1 = 32'd9527
; 
32'd188805: dataIn1 = 32'd10185
; 
32'd188806: dataIn1 = 32'd10186
; 
32'd188807: dataIn1 = 32'd2229
; 
32'd188808: dataIn1 = 32'd3688
; 
32'd188809: dataIn1 = 32'd9527
; 
32'd188810: dataIn1 = 32'd9970
; 
32'd188811: dataIn1 = 32'd10185
; 
32'd188812: dataIn1 = 32'd10186
; 
32'd188813: dataIn1 = 32'd10189
; 
32'd188814: dataIn1 = 32'd10234
; 
32'd188815: dataIn1 = 32'd2230
; 
32'd188816: dataIn1 = 32'd3690
; 
32'd188817: dataIn1 = 32'd9531
; 
32'd188818: dataIn1 = 32'd9543
; 
32'd188819: dataIn1 = 32'd9975
; 
32'd188820: dataIn1 = 32'd9999
; 
32'd188821: dataIn1 = 32'd10187
; 
32'd188822: dataIn1 = 32'd10188
; 
32'd188823: dataIn1 = 32'd10192
; 
32'd188824: dataIn1 = 32'd3686
; 
32'd188825: dataIn1 = 32'd3687
; 
32'd188826: dataIn1 = 32'd3690
; 
32'd188827: dataIn1 = 32'd9531
; 
32'd188828: dataIn1 = 32'd9974
; 
32'd188829: dataIn1 = 32'd10187
; 
32'd188830: dataIn1 = 32'd10188
; 
32'd188831: dataIn1 = 32'd3688
; 
32'd188832: dataIn1 = 32'd3691
; 
32'd188833: dataIn1 = 32'd9534
; 
32'd188834: dataIn1 = 32'd9983
; 
32'd188835: dataIn1 = 32'd10184
; 
32'd188836: dataIn1 = 32'd10186
; 
32'd188837: dataIn1 = 32'd10189
; 
32'd188838: dataIn1 = 32'd10234
; 
32'd188839: dataIn1 = 32'd3695
; 
32'd188840: dataIn1 = 32'd3697
; 
32'd188841: dataIn1 = 32'd9541
; 
32'd188842: dataIn1 = 32'd9544
; 
32'd188843: dataIn1 = 32'd9992
; 
32'd188844: dataIn1 = 32'd10190
; 
32'd188845: dataIn1 = 32'd10191
; 
32'd188846: dataIn1 = 32'd10235
; 
32'd188847: dataIn1 = 32'd2231
; 
32'd188848: dataIn1 = 32'd3697
; 
32'd188849: dataIn1 = 32'd3700
; 
32'd188850: dataIn1 = 32'd9541
; 
32'd188851: dataIn1 = 32'd10190
; 
32'd188852: dataIn1 = 32'd10191
; 
32'd188853: dataIn1 = 32'd3615
; 
32'd188854: dataIn1 = 32'd3690
; 
32'd188855: dataIn1 = 32'd3694
; 
32'd188856: dataIn1 = 32'd9543
; 
32'd188857: dataIn1 = 32'd10187
; 
32'd188858: dataIn1 = 32'd10192
; 
32'd188859: dataIn1 = 32'd2231
; 
32'd188860: dataIn1 = 32'd3699
; 
32'd188861: dataIn1 = 32'd3700
; 
32'd188862: dataIn1 = 32'd9548
; 
32'd188863: dataIn1 = 32'd10193
; 
32'd188864: dataIn1 = 32'd10194
; 
32'd188865: dataIn1 = 32'd3698
; 
32'd188866: dataIn1 = 32'd3699
; 
32'd188867: dataIn1 = 32'd9548
; 
32'd188868: dataIn1 = 32'd9551
; 
32'd188869: dataIn1 = 32'd10008
; 
32'd188870: dataIn1 = 32'd10015
; 
32'd188871: dataIn1 = 32'd10193
; 
32'd188872: dataIn1 = 32'd10194
; 
32'd188873: dataIn1 = 32'd10195
; 
32'd188874: dataIn1 = 32'd2233
; 
32'd188875: dataIn1 = 32'd3699
; 
32'd188876: dataIn1 = 32'd3702
; 
32'd188877: dataIn1 = 32'd9551
; 
32'd188878: dataIn1 = 32'd10017
; 
32'd188879: dataIn1 = 32'd10194
; 
32'd188880: dataIn1 = 32'd10195
; 
32'd188881: dataIn1 = 32'd61
; 
32'd188882: dataIn1 = 32'd3616
; 
32'd188883: dataIn1 = 32'd3619
; 
32'd188884: dataIn1 = 32'd9556
; 
32'd188885: dataIn1 = 32'd10164
; 
32'd188886: dataIn1 = 32'd10196
; 
32'd188887: dataIn1 = 32'd3732
; 
32'd188888: dataIn1 = 32'd3736
; 
32'd188889: dataIn1 = 32'd10033
; 
32'd188890: dataIn1 = 32'd10197
; 
32'd188891: dataIn1 = 32'd10198
; 
32'd188892: dataIn1 = 32'd10201
; 
32'd188893: dataIn1 = 32'd10236
; 
32'd188894: dataIn1 = 32'd2243
; 
32'd188895: dataIn1 = 32'd3732
; 
32'd188896: dataIn1 = 32'd9558
; 
32'd188897: dataIn1 = 32'd10031
; 
32'd188898: dataIn1 = 32'd10033
; 
32'd188899: dataIn1 = 32'd10197
; 
32'd188900: dataIn1 = 32'd10198
; 
32'd188901: dataIn1 = 32'd10287
; 
32'd188902: dataIn1 = 32'd2244
; 
32'd188903: dataIn1 = 32'd3742
; 
32'd188904: dataIn1 = 32'd3743
; 
32'd188905: dataIn1 = 32'd9562
; 
32'd188906: dataIn1 = 32'd10199
; 
32'd188907: dataIn1 = 32'd10200
; 
32'd188908: dataIn1 = 32'd3741
; 
32'd188909: dataIn1 = 32'd3742
; 
32'd188910: dataIn1 = 32'd9562
; 
32'd188911: dataIn1 = 32'd10038
; 
32'd188912: dataIn1 = 32'd10199
; 
32'd188913: dataIn1 = 32'd10200
; 
32'd188914: dataIn1 = 32'd10202
; 
32'd188915: dataIn1 = 32'd10237
; 
32'd188916: dataIn1 = 32'd2242
; 
32'd188917: dataIn1 = 32'd3736
; 
32'd188918: dataIn1 = 32'd9566
; 
32'd188919: dataIn1 = 32'd10046
; 
32'd188920: dataIn1 = 32'd10197
; 
32'd188921: dataIn1 = 32'd10201
; 
32'd188922: dataIn1 = 32'd10202
; 
32'd188923: dataIn1 = 32'd10236
; 
32'd188924: dataIn1 = 32'd2242
; 
32'd188925: dataIn1 = 32'd3741
; 
32'd188926: dataIn1 = 32'd9566
; 
32'd188927: dataIn1 = 32'd10044
; 
32'd188928: dataIn1 = 32'd10200
; 
32'd188929: dataIn1 = 32'd10201
; 
32'd188930: dataIn1 = 32'd10202
; 
32'd188931: dataIn1 = 32'd10237
; 
32'd188932: dataIn1 = 32'd3746
; 
32'd188933: dataIn1 = 32'd9572
; 
32'd188934: dataIn1 = 32'd9773
; 
32'd188935: dataIn1 = 32'd10056
; 
32'd188936: dataIn1 = 32'd10203
; 
32'd188937: dataIn1 = 32'd10204
; 
32'd188938: dataIn1 = 32'd10206
; 
32'd188939: dataIn1 = 32'd10238
; 
32'd188940: dataIn1 = 32'd2217
; 
32'd188941: dataIn1 = 32'd5310
; 
32'd188942: dataIn1 = 32'd9572
; 
32'd188943: dataIn1 = 32'd9773
; 
32'd188944: dataIn1 = 32'd10057
; 
32'd188945: dataIn1 = 32'd10203
; 
32'd188946: dataIn1 = 32'd10204
; 
32'd188947: dataIn1 = 32'd67
; 
32'd188948: dataIn1 = 32'd9574
; 
32'd188949: dataIn1 = 32'd9772
; 
32'd188950: dataIn1 = 32'd10062
; 
32'd188951: dataIn1 = 32'd10205
; 
32'd188952: dataIn1 = 32'd10206
; 
32'd188953: dataIn1 = 32'd10208
; 
32'd188954: dataIn1 = 32'd10239
; 
32'd188955: dataIn1 = 32'd3746
; 
32'd188956: dataIn1 = 32'd9574
; 
32'd188957: dataIn1 = 32'd9772
; 
32'd188958: dataIn1 = 32'd10061
; 
32'd188959: dataIn1 = 32'd10203
; 
32'd188960: dataIn1 = 32'd10205
; 
32'd188961: dataIn1 = 32'd10206
; 
32'd188962: dataIn1 = 32'd10238
; 
32'd188963: dataIn1 = 32'd3758
; 
32'd188964: dataIn1 = 32'd9583
; 
32'd188965: dataIn1 = 32'd9774
; 
32'd188966: dataIn1 = 32'd10076
; 
32'd188967: dataIn1 = 32'd10207
; 
32'd188968: dataIn1 = 32'd10208
; 
32'd188969: dataIn1 = 32'd10209
; 
32'd188970: dataIn1 = 32'd10240
; 
32'd188971: dataIn1 = 32'd67
; 
32'd188972: dataIn1 = 32'd9583
; 
32'd188973: dataIn1 = 32'd9774
; 
32'd188974: dataIn1 = 32'd10075
; 
32'd188975: dataIn1 = 32'd10205
; 
32'd188976: dataIn1 = 32'd10207
; 
32'd188977: dataIn1 = 32'd10208
; 
32'd188978: dataIn1 = 32'd10239
; 
32'd188979: dataIn1 = 32'd3758
; 
32'd188980: dataIn1 = 32'd9584
; 
32'd188981: dataIn1 = 32'd9775
; 
32'd188982: dataIn1 = 32'd10081
; 
32'd188983: dataIn1 = 32'd10207
; 
32'd188984: dataIn1 = 32'd10209
; 
32'd188985: dataIn1 = 32'd10210
; 
32'd188986: dataIn1 = 32'd10240
; 
32'd188987: dataIn1 = 32'd2220
; 
32'd188988: dataIn1 = 32'd9584
; 
32'd188989: dataIn1 = 32'd9775
; 
32'd188990: dataIn1 = 32'd10080
; 
32'd188991: dataIn1 = 32'd10209
; 
32'd188992: dataIn1 = 32'd10210
; 
32'd188993: dataIn1 = 32'd10212
; 
32'd188994: dataIn1 = 32'd10241
; 
32'd188995: dataIn1 = 32'd3660
; 
32'd188996: dataIn1 = 32'd3661
; 
32'd188997: dataIn1 = 32'd9588
; 
32'd188998: dataIn1 = 32'd10088
; 
32'd188999: dataIn1 = 32'd10211
; 
32'd189000: dataIn1 = 32'd10212
; 
32'd189001: dataIn1 = 32'd10214
; 
32'd189002: dataIn1 = 32'd10242
; 
32'd189003: dataIn1 = 32'd2220
; 
32'd189004: dataIn1 = 32'd3661
; 
32'd189005: dataIn1 = 32'd9588
; 
32'd189006: dataIn1 = 32'd10089
; 
32'd189007: dataIn1 = 32'd10210
; 
32'd189008: dataIn1 = 32'd10211
; 
32'd189009: dataIn1 = 32'd10212
; 
32'd189010: dataIn1 = 32'd10241
; 
32'd189011: dataIn1 = 32'd68
; 
32'd189012: dataIn1 = 32'd3659
; 
32'd189013: dataIn1 = 32'd9590
; 
32'd189014: dataIn1 = 32'd10094
; 
32'd189015: dataIn1 = 32'd10213
; 
32'd189016: dataIn1 = 32'd10214
; 
32'd189017: dataIn1 = 32'd10216
; 
32'd189018: dataIn1 = 32'd10243
; 
32'd189019: dataIn1 = 32'd3659
; 
32'd189020: dataIn1 = 32'd3660
; 
32'd189021: dataIn1 = 32'd9590
; 
32'd189022: dataIn1 = 32'd10093
; 
32'd189023: dataIn1 = 32'd10211
; 
32'd189024: dataIn1 = 32'd10213
; 
32'd189025: dataIn1 = 32'd10214
; 
32'd189026: dataIn1 = 32'd10242
; 
32'd189027: dataIn1 = 32'd3663
; 
32'd189028: dataIn1 = 32'd3667
; 
32'd189029: dataIn1 = 32'd9599
; 
32'd189030: dataIn1 = 32'd10108
; 
32'd189031: dataIn1 = 32'd10215
; 
32'd189032: dataIn1 = 32'd10216
; 
32'd189033: dataIn1 = 32'd10217
; 
32'd189034: dataIn1 = 32'd10244
; 
32'd189035: dataIn1 = 32'd68
; 
32'd189036: dataIn1 = 32'd3663
; 
32'd189037: dataIn1 = 32'd9599
; 
32'd189038: dataIn1 = 32'd10107
; 
32'd189039: dataIn1 = 32'd10213
; 
32'd189040: dataIn1 = 32'd10215
; 
32'd189041: dataIn1 = 32'd10216
; 
32'd189042: dataIn1 = 32'd10243
; 
32'd189043: dataIn1 = 32'd3665
; 
32'd189044: dataIn1 = 32'd3667
; 
32'd189045: dataIn1 = 32'd9600
; 
32'd189046: dataIn1 = 32'd10113
; 
32'd189047: dataIn1 = 32'd10215
; 
32'd189048: dataIn1 = 32'd10217
; 
32'd189049: dataIn1 = 32'd10218
; 
32'd189050: dataIn1 = 32'd10244
; 
32'd189051: dataIn1 = 32'd2223
; 
32'd189052: dataIn1 = 32'd3665
; 
32'd189053: dataIn1 = 32'd9501
; 
32'd189054: dataIn1 = 32'd9600
; 
32'd189055: dataIn1 = 32'd10112
; 
32'd189056: dataIn1 = 32'd10217
; 
32'd189057: dataIn1 = 32'd10218
; 
32'd189058: dataIn1 = 32'd10245
; 
32'd189059: dataIn1 = 32'd2250
; 
32'd189060: dataIn1 = 32'd3770
; 
32'd189061: dataIn1 = 32'd3772
; 
32'd189062: dataIn1 = 32'd9601
; 
32'd189063: dataIn1 = 32'd10174
; 
32'd189064: dataIn1 = 32'd10219
; 
32'd189065: dataIn1 = 32'd6162
; 
32'd189066: dataIn1 = 32'd6163
; 
32'd189067: dataIn1 = 32'd7262
; 
32'd189068: dataIn1 = 32'd9286
; 
32'd189069: dataIn1 = 32'd10123
; 
32'd189070: dataIn1 = 32'd10151
; 
32'd189071: dataIn1 = 32'd10220
; 
32'd189072: dataIn1 = 32'd5211
; 
32'd189073: dataIn1 = 32'd9740
; 
32'd189074: dataIn1 = 32'd9747
; 
32'd189075: dataIn1 = 32'd9748
; 
32'd189076: dataIn1 = 32'd10140
; 
32'd189077: dataIn1 = 32'd10221
; 
32'd189078: dataIn1 = 32'd1129
; 
32'd189079: dataIn1 = 32'd6678
; 
32'd189080: dataIn1 = 32'd6728
; 
32'd189081: dataIn1 = 32'd9750
; 
32'd189082: dataIn1 = 32'd10222
; 
32'd189083: dataIn1 = 32'd10223
; 
32'd189084: dataIn1 = 32'd10246
; 
32'd189085: dataIn1 = 32'd6713
; 
32'd189086: dataIn1 = 32'd6728
; 
32'd189087: dataIn1 = 32'd9750
; 
32'd189088: dataIn1 = 32'd9753
; 
32'd189089: dataIn1 = 32'd10141
; 
32'd189090: dataIn1 = 32'd10149
; 
32'd189091: dataIn1 = 32'd10222
; 
32'd189092: dataIn1 = 32'd10223
; 
32'd189093: dataIn1 = 32'd10224
; 
32'd189094: dataIn1 = 32'd5451
; 
32'd189095: dataIn1 = 32'd6728
; 
32'd189096: dataIn1 = 32'd6738
; 
32'd189097: dataIn1 = 32'd9753
; 
32'd189098: dataIn1 = 32'd10223
; 
32'd189099: dataIn1 = 32'd10224
; 
32'd189100: dataIn1 = 32'd21
; 
32'd189101: dataIn1 = 32'd2115
; 
32'd189102: dataIn1 = 32'd2117
; 
32'd189103: dataIn1 = 32'd5523
; 
32'd189104: dataIn1 = 32'd10154
; 
32'd189105: dataIn1 = 32'd10225
; 
32'd189106: dataIn1 = 32'd52
; 
32'd189107: dataIn1 = 32'd3633
; 
32'd189108: dataIn1 = 32'd3637
; 
32'd189109: dataIn1 = 32'd10158
; 
32'd189110: dataIn1 = 32'd10172
; 
32'd189111: dataIn1 = 32'd10226
; 
32'd189112: dataIn1 = 32'd9467
; 
32'd189113: dataIn1 = 32'd9770
; 
32'd189114: dataIn1 = 32'd9781
; 
32'd189115: dataIn1 = 32'd9849
; 
32'd189116: dataIn1 = 32'd10161
; 
32'd189117: dataIn1 = 32'd10227
; 
32'd189118: dataIn1 = 32'd2206
; 
32'd189119: dataIn1 = 32'd3633
; 
32'd189120: dataIn1 = 32'd3634
; 
32'd189121: dataIn1 = 32'd10167
; 
32'd189122: dataIn1 = 32'd10171
; 
32'd189123: dataIn1 = 32'd10228
; 
32'd189124: dataIn1 = 32'd3620
; 
32'd189125: dataIn1 = 32'd3623
; 
32'd189126: dataIn1 = 32'd3624
; 
32'd189127: dataIn1 = 32'd9484
; 
32'd189128: dataIn1 = 32'd10169
; 
32'd189129: dataIn1 = 32'd10229
; 
32'd189130: dataIn1 = 32'd3772
; 
32'd189131: dataIn1 = 32'd3773
; 
32'd189132: dataIn1 = 32'd3776
; 
32'd189133: dataIn1 = 32'd10173
; 
32'd189134: dataIn1 = 32'd10180
; 
32'd189135: dataIn1 = 32'd10230
; 
32'd189136: dataIn1 = 32'd2227
; 
32'd189137: dataIn1 = 32'd3672
; 
32'd189138: dataIn1 = 32'd3676
; 
32'd189139: dataIn1 = 32'd10175
; 
32'd189140: dataIn1 = 32'd10181
; 
32'd189141: dataIn1 = 32'd10231
; 
32'd189142: dataIn1 = 32'd2252
; 
32'd189143: dataIn1 = 32'd3776
; 
32'd189144: dataIn1 = 32'd3780
; 
32'd189145: dataIn1 = 32'd10177
; 
32'd189146: dataIn1 = 32'd10179
; 
32'd189147: dataIn1 = 32'd10232
; 
32'd189148: dataIn1 = 32'd2227
; 
32'd189149: dataIn1 = 32'd3680
; 
32'd189150: dataIn1 = 32'd3681
; 
32'd189151: dataIn1 = 32'd9523
; 
32'd189152: dataIn1 = 32'd10182
; 
32'd189153: dataIn1 = 32'd10233
; 
32'd189154: dataIn1 = 32'd2229
; 
32'd189155: dataIn1 = 32'd3691
; 
32'd189156: dataIn1 = 32'd3792
; 
32'd189157: dataIn1 = 32'd10186
; 
32'd189158: dataIn1 = 32'd10189
; 
32'd189159: dataIn1 = 32'd10234
; 
32'd189160: dataIn1 = 32'd71
; 
32'd189161: dataIn1 = 32'd3692
; 
32'd189162: dataIn1 = 32'd3697
; 
32'd189163: dataIn1 = 32'd9544
; 
32'd189164: dataIn1 = 32'd10190
; 
32'd189165: dataIn1 = 32'd10235
; 
32'd189166: dataIn1 = 32'd2242
; 
32'd189167: dataIn1 = 32'd3732
; 
32'd189168: dataIn1 = 32'd3733
; 
32'd189169: dataIn1 = 32'd3734
; 
32'd189170: dataIn1 = 32'd10197
; 
32'd189171: dataIn1 = 32'd10201
; 
32'd189172: dataIn1 = 32'd10236
; 
32'd189173: dataIn1 = 32'd2242
; 
32'd189174: dataIn1 = 32'd3739
; 
32'd189175: dataIn1 = 32'd3742
; 
32'd189176: dataIn1 = 32'd10200
; 
32'd189177: dataIn1 = 32'd10202
; 
32'd189178: dataIn1 = 32'd10237
; 
32'd189179: dataIn1 = 32'd2218
; 
32'd189180: dataIn1 = 32'd9772
; 
32'd189181: dataIn1 = 32'd9773
; 
32'd189182: dataIn1 = 32'd10203
; 
32'd189183: dataIn1 = 32'd10206
; 
32'd189184: dataIn1 = 32'd10238
; 
32'd189185: dataIn1 = 32'd9772
; 
32'd189186: dataIn1 = 32'd9774
; 
32'd189187: dataIn1 = 32'd9783
; 
32'd189188: dataIn1 = 32'd10205
; 
32'd189189: dataIn1 = 32'd10208
; 
32'd189190: dataIn1 = 32'd10239
; 
32'd189191: dataIn1 = 32'd2219
; 
32'd189192: dataIn1 = 32'd9774
; 
32'd189193: dataIn1 = 32'd9775
; 
32'd189194: dataIn1 = 32'd10207
; 
32'd189195: dataIn1 = 32'd10209
; 
32'd189196: dataIn1 = 32'd10240
; 
32'd189197: dataIn1 = 32'd3661
; 
32'd189198: dataIn1 = 32'd9775
; 
32'd189199: dataIn1 = 32'd9784
; 
32'd189200: dataIn1 = 32'd10210
; 
32'd189201: dataIn1 = 32'd10212
; 
32'd189202: dataIn1 = 32'd10241
; 
32'd189203: dataIn1 = 32'd2221
; 
32'd189204: dataIn1 = 32'd3659
; 
32'd189205: dataIn1 = 32'd3661
; 
32'd189206: dataIn1 = 32'd10211
; 
32'd189207: dataIn1 = 32'd10214
; 
32'd189208: dataIn1 = 32'd10242
; 
32'd189209: dataIn1 = 32'd3659
; 
32'd189210: dataIn1 = 32'd3662
; 
32'd189211: dataIn1 = 32'd3663
; 
32'd189212: dataIn1 = 32'd10213
; 
32'd189213: dataIn1 = 32'd10216
; 
32'd189214: dataIn1 = 32'd10243
; 
32'd189215: dataIn1 = 32'd2222
; 
32'd189216: dataIn1 = 32'd3663
; 
32'd189217: dataIn1 = 32'd3665
; 
32'd189218: dataIn1 = 32'd10215
; 
32'd189219: dataIn1 = 32'd10217
; 
32'd189220: dataIn1 = 32'd10244
; 
32'd189221: dataIn1 = 32'd3664
; 
32'd189222: dataIn1 = 32'd3665
; 
32'd189223: dataIn1 = 32'd3666
; 
32'd189224: dataIn1 = 32'd9501
; 
32'd189225: dataIn1 = 32'd10218
; 
32'd189226: dataIn1 = 32'd10245
; 
32'd189227: dataIn1 = 32'd5298
; 
32'd189228: dataIn1 = 32'd6678
; 
32'd189229: dataIn1 = 32'd6728
; 
32'd189230: dataIn1 = 32'd6729
; 
32'd189231: dataIn1 = 32'd10222
; 
32'd189232: dataIn1 = 32'd10246
; 
32'd189233: dataIn1 = 32'd558
; 
32'd189234: dataIn1 = 32'd1272
; 
32'd189235: dataIn1 = 32'd2101
; 
32'd189236: dataIn1 = 32'd10247
; 
32'd189237: dataIn1 = 32'd10248
; 
32'd189238: dataIn1 = 32'd10254
; 
32'd189239: dataIn1 = 32'd11656
; 
32'd189240: dataIn1 = 32'd11657
; 
32'd189241: dataIn1 = 32'd557
; 
32'd189242: dataIn1 = 32'd558
; 
32'd189243: dataIn1 = 32'd1273
; 
32'd189244: dataIn1 = 32'd2101
; 
32'd189245: dataIn1 = 32'd10247
; 
32'd189246: dataIn1 = 32'd10248
; 
32'd189247: dataIn1 = 32'd10255
; 
32'd189248: dataIn1 = 32'd267
; 
32'd189249: dataIn1 = 32'd958
; 
32'd189250: dataIn1 = 32'd1259
; 
32'd189251: dataIn1 = 32'd1266
; 
32'd189252: dataIn1 = 32'd10249
; 
32'd189253: dataIn1 = 32'd10250
; 
32'd189254: dataIn1 = 32'd10253
; 
32'd189255: dataIn1 = 32'd547
; 
32'd189256: dataIn1 = 32'd958
; 
32'd189257: dataIn1 = 32'd1259
; 
32'd189258: dataIn1 = 32'd2755
; 
32'd189259: dataIn1 = 32'd10249
; 
32'd189260: dataIn1 = 32'd10250
; 
32'd189261: dataIn1 = 32'd10269
; 
32'd189262: dataIn1 = 32'd800
; 
32'd189263: dataIn1 = 32'd981
; 
32'd189264: dataIn1 = 32'd2513
; 
32'd189265: dataIn1 = 32'd3445
; 
32'd189266: dataIn1 = 32'd10251
; 
32'd189267: dataIn1 = 32'd10252
; 
32'd189268: dataIn1 = 32'd10264
; 
32'd189269: dataIn1 = 32'd806
; 
32'd189270: dataIn1 = 32'd981
; 
32'd189271: dataIn1 = 32'd2521
; 
32'd189272: dataIn1 = 32'd3445
; 
32'd189273: dataIn1 = 32'd10251
; 
32'd189274: dataIn1 = 32'd10252
; 
32'd189275: dataIn1 = 32'd10265
; 
32'd189276: dataIn1 = 32'd550
; 
32'd189277: dataIn1 = 32'd958
; 
32'd189278: dataIn1 = 32'd959
; 
32'd189279: dataIn1 = 32'd1266
; 
32'd189280: dataIn1 = 32'd10249
; 
32'd189281: dataIn1 = 32'd10253
; 
32'd189282: dataIn1 = 32'd556
; 
32'd189283: dataIn1 = 32'd558
; 
32'd189284: dataIn1 = 32'd960
; 
32'd189285: dataIn1 = 32'd1272
; 
32'd189286: dataIn1 = 32'd10247
; 
32'd189287: dataIn1 = 32'd10254
; 
32'd189288: dataIn1 = 32'd268
; 
32'd189289: dataIn1 = 32'd555
; 
32'd189290: dataIn1 = 32'd558
; 
32'd189291: dataIn1 = 32'd1273
; 
32'd189292: dataIn1 = 32'd10248
; 
32'd189293: dataIn1 = 32'd10255
; 
32'd189294: dataIn1 = 32'd1854
; 
32'd189295: dataIn1 = 32'd1855
; 
32'd189296: dataIn1 = 32'd3030
; 
32'd189297: dataIn1 = 32'd3460
; 
32'd189298: dataIn1 = 32'd10256
; 
32'd189299: dataIn1 = 32'd10257
; 
32'd189300: dataIn1 = 32'd10271
; 
32'd189301: dataIn1 = 32'd391
; 
32'd189302: dataIn1 = 32'd1855
; 
32'd189303: dataIn1 = 32'd3030
; 
32'd189304: dataIn1 = 32'd4611
; 
32'd189305: dataIn1 = 32'd10256
; 
32'd189306: dataIn1 = 32'd10257
; 
32'd189307: dataIn1 = 32'd10263
; 
32'd189308: dataIn1 = 32'd758
; 
32'd189309: dataIn1 = 32'd1858
; 
32'd189310: dataIn1 = 32'd3411
; 
32'd189311: dataIn1 = 32'd3469
; 
32'd189312: dataIn1 = 32'd10258
; 
32'd189313: dataIn1 = 32'd10259
; 
32'd189314: dataIn1 = 32'd10270
; 
32'd189315: dataIn1 = 32'd397
; 
32'd189316: dataIn1 = 32'd1470
; 
32'd189317: dataIn1 = 32'd1858
; 
32'd189318: dataIn1 = 32'd3469
; 
32'd189319: dataIn1 = 32'd10258
; 
32'd189320: dataIn1 = 32'd10259
; 
32'd189321: dataIn1 = 32'd10284
; 
32'd189322: dataIn1 = 32'd1869
; 
32'd189323: dataIn1 = 32'd1874
; 
32'd189324: dataIn1 = 32'd3418
; 
32'd189325: dataIn1 = 32'd3444
; 
32'd189326: dataIn1 = 32'd10260
; 
32'd189327: dataIn1 = 32'd10261
; 
32'd189328: dataIn1 = 32'd10262
; 
32'd189329: dataIn1 = 32'd1874
; 
32'd189330: dataIn1 = 32'd2048
; 
32'd189331: dataIn1 = 32'd3418
; 
32'd189332: dataIn1 = 32'd4629
; 
32'd189333: dataIn1 = 32'd10260
; 
32'd189334: dataIn1 = 32'd10261
; 
32'd189335: dataIn1 = 32'd10273
; 
32'd189336: dataIn1 = 32'd211
; 
32'd189337: dataIn1 = 32'd1508
; 
32'd189338: dataIn1 = 32'd1874
; 
32'd189339: dataIn1 = 32'd3444
; 
32'd189340: dataIn1 = 32'd10260
; 
32'd189341: dataIn1 = 32'd10262
; 
32'd189342: dataIn1 = 32'd10285
; 
32'd189343: dataIn1 = 32'd1855
; 
32'd189344: dataIn1 = 32'd2287
; 
32'd189345: dataIn1 = 32'd3863
; 
32'd189346: dataIn1 = 32'd4611
; 
32'd189347: dataIn1 = 32'd10257
; 
32'd189348: dataIn1 = 32'd10263
; 
32'd189349: dataIn1 = 32'd10272
; 
32'd189350: dataIn1 = 32'd413
; 
32'd189351: dataIn1 = 32'd981
; 
32'd189352: dataIn1 = 32'd2513
; 
32'd189353: dataIn1 = 32'd3429
; 
32'd189354: dataIn1 = 32'd10251
; 
32'd189355: dataIn1 = 32'd10264
; 
32'd189356: dataIn1 = 32'd156
; 
32'd189357: dataIn1 = 32'd981
; 
32'd189358: dataIn1 = 32'd2521
; 
32'd189359: dataIn1 = 32'd3454
; 
32'd189360: dataIn1 = 32'd10252
; 
32'd189361: dataIn1 = 32'd10265
; 
32'd189362: dataIn1 = 32'd2567
; 
32'd189363: dataIn1 = 32'd2570
; 
32'd189364: dataIn1 = 32'd4683
; 
32'd189365: dataIn1 = 32'd4856
; 
32'd189366: dataIn1 = 32'd10266
; 
32'd189367: dataIn1 = 32'd10267
; 
32'd189368: dataIn1 = 32'd10268
; 
32'd189369: dataIn1 = 32'd1042
; 
32'd189370: dataIn1 = 32'd2567
; 
32'd189371: dataIn1 = 32'd4683
; 
32'd189372: dataIn1 = 32'd5429
; 
32'd189373: dataIn1 = 32'd10266
; 
32'd189374: dataIn1 = 32'd10267
; 
32'd189375: dataIn1 = 32'd10275
; 
32'd189376: dataIn1 = 32'd1076
; 
32'd189377: dataIn1 = 32'd2567
; 
32'd189378: dataIn1 = 32'd4677
; 
32'd189379: dataIn1 = 32'd4856
; 
32'd189380: dataIn1 = 32'd10266
; 
32'd189381: dataIn1 = 32'd10268
; 
32'd189382: dataIn1 = 32'd10274
; 
32'd189383: dataIn1 = 32'd266
; 
32'd189384: dataIn1 = 32'd548
; 
32'd189385: dataIn1 = 32'd958
; 
32'd189386: dataIn1 = 32'd2755
; 
32'd189387: dataIn1 = 32'd10250
; 
32'd189388: dataIn1 = 32'd10269
; 
32'd189389: dataIn1 = 32'd393
; 
32'd189390: dataIn1 = 32'd1857
; 
32'd189391: dataIn1 = 32'd1858
; 
32'd189392: dataIn1 = 32'd3411
; 
32'd189393: dataIn1 = 32'd10258
; 
32'd189394: dataIn1 = 32'd10270
; 
32'd189395: dataIn1 = 32'd392
; 
32'd189396: dataIn1 = 32'd749
; 
32'd189397: dataIn1 = 32'd1855
; 
32'd189398: dataIn1 = 32'd3460
; 
32'd189399: dataIn1 = 32'd10256
; 
32'd189400: dataIn1 = 32'd10271
; 
32'd189401: dataIn1 = 32'd392
; 
32'd189402: dataIn1 = 32'd1855
; 
32'd189403: dataIn1 = 32'd2286
; 
32'd189404: dataIn1 = 32'd3863
; 
32'd189405: dataIn1 = 32'd10263
; 
32'd189406: dataIn1 = 32'd10272
; 
32'd189407: dataIn1 = 32'd983
; 
32'd189408: dataIn1 = 32'd1873
; 
32'd189409: dataIn1 = 32'd1874
; 
32'd189410: dataIn1 = 32'd4629
; 
32'd189411: dataIn1 = 32'd10261
; 
32'd189412: dataIn1 = 32'd10273
; 
32'd189413: dataIn1 = 32'd2565
; 
32'd189414: dataIn1 = 32'd2566
; 
32'd189415: dataIn1 = 32'd2567
; 
32'd189416: dataIn1 = 32'd4677
; 
32'd189417: dataIn1 = 32'd10268
; 
32'd189418: dataIn1 = 32'd10274
; 
32'd189419: dataIn1 = 32'd212
; 
32'd189420: dataIn1 = 32'd2565
; 
32'd189421: dataIn1 = 32'd2567
; 
32'd189422: dataIn1 = 32'd5429
; 
32'd189423: dataIn1 = 32'd10267
; 
32'd189424: dataIn1 = 32'd10275
; 
32'd189425: dataIn1 = 32'd1141
; 
32'd189426: dataIn1 = 32'd5520
; 
32'd189427: dataIn1 = 32'd9672
; 
32'd189428: dataIn1 = 32'd9823
; 
32'd189429: dataIn1 = 32'd10276
; 
32'd189430: dataIn1 = 32'd10277
; 
32'd189431: dataIn1 = 32'd10283
; 
32'd189432: dataIn1 = 32'd1141
; 
32'd189433: dataIn1 = 32'd5451
; 
32'd189434: dataIn1 = 32'd9325
; 
32'd189435: dataIn1 = 32'd9672
; 
32'd189436: dataIn1 = 32'd10276
; 
32'd189437: dataIn1 = 32'd10277
; 
32'd189438: dataIn1 = 32'd10281
; 
32'd189439: dataIn1 = 32'd5210
; 
32'd189440: dataIn1 = 32'd6396
; 
32'd189441: dataIn1 = 32'd8307
; 
32'd189442: dataIn1 = 32'd9766
; 
32'd189443: dataIn1 = 32'd10278
; 
32'd189444: dataIn1 = 32'd10279
; 
32'd189445: dataIn1 = 32'd10280
; 
32'd189446: dataIn1 = 32'd6392
; 
32'd189447: dataIn1 = 32'd6396
; 
32'd189448: dataIn1 = 32'd9741
; 
32'd189449: dataIn1 = 32'd9766
; 
32'd189450: dataIn1 = 32'd10278
; 
32'd189451: dataIn1 = 32'd10279
; 
32'd189452: dataIn1 = 32'd10282
; 
32'd189453: dataIn1 = 32'd6396
; 
32'd189454: dataIn1 = 32'd6440
; 
32'd189455: dataIn1 = 32'd6443
; 
32'd189456: dataIn1 = 32'd8307
; 
32'd189457: dataIn1 = 32'd10278
; 
32'd189458: dataIn1 = 32'd10280
; 
32'd189459: dataIn1 = 32'd1141
; 
32'd189460: dataIn1 = 32'd5452
; 
32'd189461: dataIn1 = 32'd5523
; 
32'd189462: dataIn1 = 32'd9325
; 
32'd189463: dataIn1 = 32'd10277
; 
32'd189464: dataIn1 = 32'd10281
; 
32'd189465: dataIn1 = 32'd1129
; 
32'd189466: dataIn1 = 32'd6395
; 
32'd189467: dataIn1 = 32'd6396
; 
32'd189468: dataIn1 = 32'd9741
; 
32'd189469: dataIn1 = 32'd10279
; 
32'd189470: dataIn1 = 32'd10282
; 
32'd189471: dataIn1 = 32'd1141
; 
32'd189472: dataIn1 = 32'd9456
; 
32'd189473: dataIn1 = 32'd9823
; 
32'd189474: dataIn1 = 32'd10154
; 
32'd189475: dataIn1 = 32'd10276
; 
32'd189476: dataIn1 = 32'd10283
; 
32'd189477: dataIn1 = 32'd771
; 
32'd189478: dataIn1 = 32'd1470
; 
32'd189479: dataIn1 = 32'd1858
; 
32'd189480: dataIn1 = 32'd1859
; 
32'd189481: dataIn1 = 32'd10259
; 
32'd189482: dataIn1 = 32'd10284
; 
32'd189483: dataIn1 = 32'd801
; 
32'd189484: dataIn1 = 32'd1508
; 
32'd189485: dataIn1 = 32'd1873
; 
32'd189486: dataIn1 = 32'd1874
; 
32'd189487: dataIn1 = 32'd10262
; 
32'd189488: dataIn1 = 32'd10285
; 
32'd189489: dataIn1 = 32'd2103
; 
32'd189490: dataIn1 = 32'd6826
; 
32'd189491: dataIn1 = 32'd9264
; 
32'd189492: dataIn1 = 32'd9313
; 
32'd189493: dataIn1 = 32'd10286
; 
32'd189494: dataIn1 = 32'd2243
; 
32'd189495: dataIn1 = 32'd3735
; 
32'd189496: dataIn1 = 32'd10031
; 
32'd189497: dataIn1 = 32'd10198
; 
32'd189498: dataIn1 = 32'd10287
; 
32'd189499: dataIn1 = 32'd87
; 
32'd189500: dataIn1 = 32'd97
; 
32'd189501: dataIn1 = 32'd5315
; 
32'd189502: dataIn1 = 32'd10288
; 
32'd189503: dataIn1 = 32'd99
; 
32'd189504: dataIn1 = 32'd100
; 
32'd189505: dataIn1 = 32'd5316
; 
32'd189506: dataIn1 = 32'd10289
; 
32'd189507: dataIn1 = 32'd2105
; 
32'd189508: dataIn1 = 32'd9266
; 
32'd189509: dataIn1 = 32'd9316
; 
32'd189510: dataIn1 = 32'd10290
; 
32'd189511: dataIn1 = 32'd2105
; 
32'd189512: dataIn1 = 32'd5646
; 
32'd189513: dataIn1 = 32'd6843
; 
32'd189514: dataIn1 = 32'd9438
; 
32'd189515: dataIn1 = 32'd10291
; 
32'd189516: dataIn1 = 32'd250
; 
32'd189517: dataIn1 = 32'd957
; 
32'd189518: dataIn1 = 32'd10292
; 
32'd189519: dataIn1 = 32'd10293
; 
32'd189520: dataIn1 = 32'd250
; 
32'd189521: dataIn1 = 32'd954
; 
32'd189522: dataIn1 = 32'd957
; 
32'd189523: dataIn1 = 32'd1714
; 
32'd189524: dataIn1 = 32'd1719
; 
32'd189525: dataIn1 = 32'd10292
; 
32'd189526: dataIn1 = 32'd10293
; 
32'd189527: dataIn1 = 32'd10294
; 
32'd189528: dataIn1 = 32'd953
; 
32'd189529: dataIn1 = 32'd954
; 
32'd189530: dataIn1 = 32'd1712
; 
32'd189531: dataIn1 = 32'd1719
; 
32'd189532: dataIn1 = 32'd10293
; 
32'd189533: dataIn1 = 32'd10294
; 
32'd189534: dataIn1 = 32'd10295
; 
32'd189535: dataIn1 = 32'd951
; 
32'd189536: dataIn1 = 32'd954
; 
32'd189537: dataIn1 = 32'd1712
; 
32'd189538: dataIn1 = 32'd1713
; 
32'd189539: dataIn1 = 32'd10294
; 
32'd189540: dataIn1 = 32'd10295
; 
32'd189541: dataIn1 = 32'd10296
; 
32'd189542: dataIn1 = 32'd441
; 
32'd189543: dataIn1 = 32'd951
; 
32'd189544: dataIn1 = 32'd1711
; 
32'd189545: dataIn1 = 32'd1713
; 
32'd189546: dataIn1 = 32'd10295
; 
32'd189547: dataIn1 = 32'd10296
; 
32'd189548: dataIn1 = 32'd10297
; 
32'd189549: dataIn1 = 32'd441
; 
32'd189550: dataIn1 = 32'd952
; 
32'd189551: dataIn1 = 32'd1711
; 
32'd189552: dataIn1 = 32'd1716
; 
32'd189553: dataIn1 = 32'd10296
; 
32'd189554: dataIn1 = 32'd10297
; 
32'd189555: dataIn1 = 32'd10298
; 
32'd189556: dataIn1 = 32'd952
; 
32'd189557: dataIn1 = 32'd956
; 
32'd189558: dataIn1 = 32'd1715
; 
32'd189559: dataIn1 = 32'd1716
; 
32'd189560: dataIn1 = 32'd10297
; 
32'd189561: dataIn1 = 32'd10298
; 
32'd189562: dataIn1 = 32'd10299
; 
32'd189563: dataIn1 = 32'd955
; 
32'd189564: dataIn1 = 32'd956
; 
32'd189565: dataIn1 = 32'd1715
; 
32'd189566: dataIn1 = 32'd1717
; 
32'd189567: dataIn1 = 32'd10298
; 
32'd189568: dataIn1 = 32'd10299
; 
32'd189569: dataIn1 = 32'd10300
; 
32'd189570: dataIn1 = 32'd249
; 
32'd189571: dataIn1 = 32'd955
; 
32'd189572: dataIn1 = 32'd1717
; 
32'd189573: dataIn1 = 32'd1718
; 
32'd189574: dataIn1 = 32'd10299
; 
32'd189575: dataIn1 = 32'd10300
; 
32'd189576: dataIn1 = 32'd10301
; 
32'd189577: dataIn1 = 32'd249
; 
32'd189578: dataIn1 = 32'd944
; 
32'd189579: dataIn1 = 32'd1701
; 
32'd189580: dataIn1 = 32'd1718
; 
32'd189581: dataIn1 = 32'd10300
; 
32'd189582: dataIn1 = 32'd10301
; 
32'd189583: dataIn1 = 32'd10302
; 
32'd189584: dataIn1 = 32'd943
; 
32'd189585: dataIn1 = 32'd944
; 
32'd189586: dataIn1 = 32'd1699
; 
32'd189587: dataIn1 = 32'd1701
; 
32'd189588: dataIn1 = 32'd10301
; 
32'd189589: dataIn1 = 32'd10302
; 
32'd189590: dataIn1 = 32'd10303
; 
32'd189591: dataIn1 = 32'd940
; 
32'd189592: dataIn1 = 32'd943
; 
32'd189593: dataIn1 = 32'd1699
; 
32'd189594: dataIn1 = 32'd1700
; 
32'd189595: dataIn1 = 32'd10302
; 
32'd189596: dataIn1 = 32'd10303
; 
32'd189597: dataIn1 = 32'd10304
; 
32'd189598: dataIn1 = 32'd439
; 
32'd189599: dataIn1 = 32'd940
; 
32'd189600: dataIn1 = 32'd1695
; 
32'd189601: dataIn1 = 32'd1700
; 
32'd189602: dataIn1 = 32'd10303
; 
32'd189603: dataIn1 = 32'd10304
; 
32'd189604: dataIn1 = 32'd10305
; 
32'd189605: dataIn1 = 32'd439
; 
32'd189606: dataIn1 = 32'd939
; 
32'd189607: dataIn1 = 32'd1695
; 
32'd189608: dataIn1 = 32'd1698
; 
32'd189609: dataIn1 = 32'd10304
; 
32'd189610: dataIn1 = 32'd10305
; 
32'd189611: dataIn1 = 32'd10306
; 
32'd189612: dataIn1 = 32'd939
; 
32'd189613: dataIn1 = 32'd942
; 
32'd189614: dataIn1 = 32'd1696
; 
32'd189615: dataIn1 = 32'd1698
; 
32'd189616: dataIn1 = 32'd10305
; 
32'd189617: dataIn1 = 32'd10306
; 
32'd189618: dataIn1 = 32'd10307
; 
32'd189619: dataIn1 = 32'd247
; 
32'd189620: dataIn1 = 32'd942
; 
32'd189621: dataIn1 = 32'd1696
; 
32'd189622: dataIn1 = 32'd1697
; 
32'd189623: dataIn1 = 32'd10306
; 
32'd189624: dataIn1 = 32'd10307
; 
32'd189625: dataIn1 = 32'd10308
; 
32'd189626: dataIn1 = 32'd247
; 
32'd189627: dataIn1 = 32'd941
; 
32'd189628: dataIn1 = 32'd1696
; 
32'd189629: dataIn1 = 32'd1704
; 
32'd189630: dataIn1 = 32'd10307
; 
32'd189631: dataIn1 = 32'd10308
; 
32'd189632: dataIn1 = 32'd10309
; 
32'd189633: dataIn1 = 32'd941
; 
32'd189634: dataIn1 = 32'd948
; 
32'd189635: dataIn1 = 32'd1704
; 
32'd189636: dataIn1 = 32'd1710
; 
32'd189637: dataIn1 = 32'd10308
; 
32'd189638: dataIn1 = 32'd10309
; 
32'd189639: dataIn1 = 32'd10310
; 
32'd189640: dataIn1 = 32'd947
; 
32'd189641: dataIn1 = 32'd948
; 
32'd189642: dataIn1 = 32'd1703
; 
32'd189643: dataIn1 = 32'd1704
; 
32'd189644: dataIn1 = 32'd10309
; 
32'd189645: dataIn1 = 32'd10310
; 
32'd189646: dataIn1 = 32'd10311
; 
32'd189647: dataIn1 = 32'd945
; 
32'd189648: dataIn1 = 32'd947
; 
32'd189649: dataIn1 = 32'd1703
; 
32'd189650: dataIn1 = 32'd1705
; 
32'd189651: dataIn1 = 32'd10310
; 
32'd189652: dataIn1 = 32'd10311
; 
32'd189653: dataIn1 = 32'd10312
; 
32'd189654: dataIn1 = 32'd440
; 
32'd189655: dataIn1 = 32'd945
; 
32'd189656: dataIn1 = 32'd1705
; 
32'd189657: dataIn1 = 32'd1708
; 
32'd189658: dataIn1 = 32'd10311
; 
32'd189659: dataIn1 = 32'd10312
; 
32'd189660: dataIn1 = 32'd10313
; 
32'd189661: dataIn1 = 32'd945
; 
32'd189662: dataIn1 = 32'd949
; 
32'd189663: dataIn1 = 32'd1702
; 
32'd189664: dataIn1 = 32'd1708
; 
32'd189665: dataIn1 = 32'd10312
; 
32'd189666: dataIn1 = 32'd10313
; 
32'd189667: dataIn1 = 32'd10314
; 
32'd189668: dataIn1 = 32'd946
; 
32'd189669: dataIn1 = 32'd949
; 
32'd189670: dataIn1 = 32'd1702
; 
32'd189671: dataIn1 = 32'd1707
; 
32'd189672: dataIn1 = 32'd10313
; 
32'd189673: dataIn1 = 32'd10314
; 
32'd189674: dataIn1 = 32'd10315
; 
32'd189675: dataIn1 = 32'd246
; 
32'd189676: dataIn1 = 32'd946
; 
32'd189677: dataIn1 = 32'd1706
; 
32'd189678: dataIn1 = 32'd1707
; 
32'd189679: dataIn1 = 32'd10314
; 
32'd189680: dataIn1 = 32'd10315
; 
32'd189681: dataIn1 = 32'd10316
; 
32'd189682: dataIn1 = 32'd246
; 
32'd189683: dataIn1 = 32'd950
; 
32'd189684: dataIn1 = 32'd1706
; 
32'd189685: dataIn1 = 32'd1709
; 
32'd189686: dataIn1 = 32'd10315
; 
32'd189687: dataIn1 = 32'd10316
; 
32'd189688: dataIn1 = 32'd10317
; 
32'd189689: dataIn1 = 32'd246
; 
32'd189690: dataIn1 = 32'd937
; 
32'd189691: dataIn1 = 32'd1694
; 
32'd189692: dataIn1 = 32'd1709
; 
32'd189693: dataIn1 = 32'd10316
; 
32'd189694: dataIn1 = 32'd10317
; 
32'd189695: dataIn1 = 32'd10318
; 
32'd189696: dataIn1 = 32'd937
; 
32'd189697: dataIn1 = 32'd938
; 
32'd189698: dataIn1 = 32'd1692
; 
32'd189699: dataIn1 = 32'd1694
; 
32'd189700: dataIn1 = 32'd10317
; 
32'd189701: dataIn1 = 32'd10318
; 
32'd189702: dataIn1 = 32'd10319
; 
32'd189703: dataIn1 = 32'd935
; 
32'd189704: dataIn1 = 32'd938
; 
32'd189705: dataIn1 = 32'd1692
; 
32'd189706: dataIn1 = 32'd1693
; 
32'd189707: dataIn1 = 32'd10318
; 
32'd189708: dataIn1 = 32'd10319
; 
32'd189709: dataIn1 = 32'd10320
; 
32'd189710: dataIn1 = 32'd438
; 
32'd189711: dataIn1 = 32'd935
; 
32'd189712: dataIn1 = 32'd1688
; 
32'd189713: dataIn1 = 32'd1693
; 
32'd189714: dataIn1 = 32'd10319
; 
32'd189715: dataIn1 = 32'd10320
; 
32'd189716: dataIn1 = 32'd10321
; 
32'd189717: dataIn1 = 32'd438
; 
32'd189718: dataIn1 = 32'd934
; 
32'd189719: dataIn1 = 32'd1688
; 
32'd189720: dataIn1 = 32'd1690
; 
32'd189721: dataIn1 = 32'd10320
; 
32'd189722: dataIn1 = 32'd10321
; 
32'd189723: dataIn1 = 32'd10322
; 
32'd189724: dataIn1 = 32'd934
; 
32'd189725: dataIn1 = 32'd936
; 
32'd189726: dataIn1 = 32'd1689
; 
32'd189727: dataIn1 = 32'd1690
; 
32'd189728: dataIn1 = 32'd10321
; 
32'd189729: dataIn1 = 32'd10322
; 
32'd189730: dataIn1 = 32'd10323
; 
32'd189731: dataIn1 = 32'd933
; 
32'd189732: dataIn1 = 32'd936
; 
32'd189733: dataIn1 = 32'd1689
; 
32'd189734: dataIn1 = 32'd1691
; 
32'd189735: dataIn1 = 32'd10322
; 
32'd189736: dataIn1 = 32'd10323
; 
32'd189737: dataIn1 = 32'd10324
; 
32'd189738: dataIn1 = 32'd244
; 
32'd189739: dataIn1 = 32'd933
; 
32'd189740: dataIn1 = 32'd1687
; 
32'd189741: dataIn1 = 32'd1691
; 
32'd189742: dataIn1 = 32'd10323
; 
32'd189743: dataIn1 = 32'd10324
; 
32'd189744: dataIn1 = 32'd10325
; 
32'd189745: dataIn1 = 32'd244
; 
32'd189746: dataIn1 = 32'd929
; 
32'd189747: dataIn1 = 32'd1682
; 
32'd189748: dataIn1 = 32'd1687
; 
32'd189749: dataIn1 = 32'd10324
; 
32'd189750: dataIn1 = 32'd10325
; 
32'd189751: dataIn1 = 32'd10326
; 
32'd189752: dataIn1 = 32'd929
; 
32'd189753: dataIn1 = 32'd930
; 
32'd189754: dataIn1 = 32'd1680
; 
32'd189755: dataIn1 = 32'd1682
; 
32'd189756: dataIn1 = 32'd10325
; 
32'd189757: dataIn1 = 32'd10326
; 
32'd189758: dataIn1 = 32'd10327
; 
32'd189759: dataIn1 = 32'd927
; 
32'd189760: dataIn1 = 32'd930
; 
32'd189761: dataIn1 = 32'd1680
; 
32'd189762: dataIn1 = 32'd1681
; 
32'd189763: dataIn1 = 32'd10326
; 
32'd189764: dataIn1 = 32'd10327
; 
32'd189765: dataIn1 = 32'd10328
; 
32'd189766: dataIn1 = 32'd437
; 
32'd189767: dataIn1 = 32'd927
; 
32'd189768: dataIn1 = 32'd1679
; 
32'd189769: dataIn1 = 32'd1681
; 
32'd189770: dataIn1 = 32'd10327
; 
32'd189771: dataIn1 = 32'd10328
; 
32'd189772: dataIn1 = 32'd10329
; 
32'd189773: dataIn1 = 32'd437
; 
32'd189774: dataIn1 = 32'd928
; 
32'd189775: dataIn1 = 32'd1679
; 
32'd189776: dataIn1 = 32'd1684
; 
32'd189777: dataIn1 = 32'd10328
; 
32'd189778: dataIn1 = 32'd10329
; 
32'd189779: dataIn1 = 32'd10330
; 
32'd189780: dataIn1 = 32'd928
; 
32'd189781: dataIn1 = 32'd932
; 
32'd189782: dataIn1 = 32'd1683
; 
32'd189783: dataIn1 = 32'd1684
; 
32'd189784: dataIn1 = 32'd10329
; 
32'd189785: dataIn1 = 32'd10330
; 
32'd189786: dataIn1 = 32'd10331
; 
32'd189787: dataIn1 = 32'd931
; 
32'd189788: dataIn1 = 32'd932
; 
32'd189789: dataIn1 = 32'd1683
; 
32'd189790: dataIn1 = 32'd1685
; 
32'd189791: dataIn1 = 32'd10330
; 
32'd189792: dataIn1 = 32'd10331
; 
32'd189793: dataIn1 = 32'd10332
; 
32'd189794: dataIn1 = 32'd243
; 
32'd189795: dataIn1 = 32'd931
; 
32'd189796: dataIn1 = 32'd1685
; 
32'd189797: dataIn1 = 32'd1686
; 
32'd189798: dataIn1 = 32'd10331
; 
32'd189799: dataIn1 = 32'd10332
; 
32'd189800: dataIn1 = 32'd10333
; 
32'd189801: dataIn1 = 32'd243
; 
32'd189802: dataIn1 = 32'd920
; 
32'd189803: dataIn1 = 32'd1669
; 
32'd189804: dataIn1 = 32'd1686
; 
32'd189805: dataIn1 = 32'd10332
; 
32'd189806: dataIn1 = 32'd10333
; 
32'd189807: dataIn1 = 32'd10334
; 
32'd189808: dataIn1 = 32'd919
; 
32'd189809: dataIn1 = 32'd920
; 
32'd189810: dataIn1 = 32'd1667
; 
32'd189811: dataIn1 = 32'd1669
; 
32'd189812: dataIn1 = 32'd10333
; 
32'd189813: dataIn1 = 32'd10334
; 
32'd189814: dataIn1 = 32'd10335
; 
32'd189815: dataIn1 = 32'd916
; 
32'd189816: dataIn1 = 32'd919
; 
32'd189817: dataIn1 = 32'd1667
; 
32'd189818: dataIn1 = 32'd1668
; 
32'd189819: dataIn1 = 32'd10334
; 
32'd189820: dataIn1 = 32'd10335
; 
32'd189821: dataIn1 = 32'd10336
; 
32'd189822: dataIn1 = 32'd435
; 
32'd189823: dataIn1 = 32'd916
; 
32'd189824: dataIn1 = 32'd1663
; 
32'd189825: dataIn1 = 32'd1668
; 
32'd189826: dataIn1 = 32'd10335
; 
32'd189827: dataIn1 = 32'd10336
; 
32'd189828: dataIn1 = 32'd10337
; 
32'd189829: dataIn1 = 32'd435
; 
32'd189830: dataIn1 = 32'd915
; 
32'd189831: dataIn1 = 32'd1663
; 
32'd189832: dataIn1 = 32'd1666
; 
32'd189833: dataIn1 = 32'd10336
; 
32'd189834: dataIn1 = 32'd10337
; 
32'd189835: dataIn1 = 32'd10338
; 
32'd189836: dataIn1 = 32'd915
; 
32'd189837: dataIn1 = 32'd918
; 
32'd189838: dataIn1 = 32'd1664
; 
32'd189839: dataIn1 = 32'd1666
; 
32'd189840: dataIn1 = 32'd10337
; 
32'd189841: dataIn1 = 32'd10338
; 
32'd189842: dataIn1 = 32'd10339
; 
32'd189843: dataIn1 = 32'd917
; 
32'd189844: dataIn1 = 32'd918
; 
32'd189845: dataIn1 = 32'd1664
; 
32'd189846: dataIn1 = 32'd1665
; 
32'd189847: dataIn1 = 32'd10338
; 
32'd189848: dataIn1 = 32'd10339
; 
32'd189849: dataIn1 = 32'd10340
; 
32'd189850: dataIn1 = 32'd241
; 
32'd189851: dataIn1 = 32'd917
; 
32'd189852: dataIn1 = 32'd1665
; 
32'd189853: dataIn1 = 32'd1678
; 
32'd189854: dataIn1 = 32'd10339
; 
32'd189855: dataIn1 = 32'd10340
; 
32'd189856: dataIn1 = 32'd10341
; 
32'd189857: dataIn1 = 32'd241
; 
32'd189858: dataIn1 = 32'd924
; 
32'd189859: dataIn1 = 32'd1672
; 
32'd189860: dataIn1 = 32'd1678
; 
32'd189861: dataIn1 = 32'd10340
; 
32'd189862: dataIn1 = 32'd10341
; 
32'd189863: dataIn1 = 32'd10342
; 
32'd189864: dataIn1 = 32'd923
; 
32'd189865: dataIn1 = 32'd924
; 
32'd189866: dataIn1 = 32'd1671
; 
32'd189867: dataIn1 = 32'd1672
; 
32'd189868: dataIn1 = 32'd10341
; 
32'd189869: dataIn1 = 32'd10342
; 
32'd189870: dataIn1 = 32'd10343
; 
32'd189871: dataIn1 = 32'd921
; 
32'd189872: dataIn1 = 32'd923
; 
32'd189873: dataIn1 = 32'd1671
; 
32'd189874: dataIn1 = 32'd1673
; 
32'd189875: dataIn1 = 32'd10342
; 
32'd189876: dataIn1 = 32'd10343
; 
32'd189877: dataIn1 = 32'd10344
; 
32'd189878: dataIn1 = 32'd436
; 
32'd189879: dataIn1 = 32'd921
; 
32'd189880: dataIn1 = 32'd1670
; 
32'd189881: dataIn1 = 32'd1673
; 
32'd189882: dataIn1 = 32'd10343
; 
32'd189883: dataIn1 = 32'd10344
; 
32'd189884: dataIn1 = 32'd10345
; 
32'd189885: dataIn1 = 32'd436
; 
32'd189886: dataIn1 = 32'd922
; 
32'd189887: dataIn1 = 32'd1670
; 
32'd189888: dataIn1 = 32'd1676
; 
32'd189889: dataIn1 = 32'd10344
; 
32'd189890: dataIn1 = 32'd10345
; 
32'd189891: dataIn1 = 32'd10346
; 
32'd189892: dataIn1 = 32'd922
; 
32'd189893: dataIn1 = 32'd925
; 
32'd189894: dataIn1 = 32'd1674
; 
32'd189895: dataIn1 = 32'd1676
; 
32'd189896: dataIn1 = 32'd10345
; 
32'd189897: dataIn1 = 32'd10346
; 
32'd189898: dataIn1 = 32'd10347
; 
32'd189899: dataIn1 = 32'd925
; 
32'd189900: dataIn1 = 32'd926
; 
32'd189901: dataIn1 = 32'd1674
; 
32'd189902: dataIn1 = 32'd1675
; 
32'd189903: dataIn1 = 32'd10346
; 
32'd189904: dataIn1 = 32'd10347
; 
32'd189905: dataIn1 = 32'd10348
; 
32'd189906: dataIn1 = 32'd240
; 
32'd189907: dataIn1 = 32'd926
; 
32'd189908: dataIn1 = 32'd1675
; 
32'd189909: dataIn1 = 32'd1677
; 
32'd189910: dataIn1 = 32'd10347
; 
32'd189911: dataIn1 = 32'd10348
; 
32'd189912: dataIn1 = 32'd10349
; 
32'd189913: dataIn1 = 32'd240
; 
32'd189914: dataIn1 = 32'd913
; 
32'd189915: dataIn1 = 32'd1662
; 
32'd189916: dataIn1 = 32'd1677
; 
32'd189917: dataIn1 = 32'd10348
; 
32'd189918: dataIn1 = 32'd10349
; 
32'd189919: dataIn1 = 32'd10350
; 
32'd189920: dataIn1 = 32'd913
; 
32'd189921: dataIn1 = 32'd914
; 
32'd189922: dataIn1 = 32'd1660
; 
32'd189923: dataIn1 = 32'd1662
; 
32'd189924: dataIn1 = 32'd10349
; 
32'd189925: dataIn1 = 32'd10350
; 
32'd189926: dataIn1 = 32'd10351
; 
32'd189927: dataIn1 = 32'd911
; 
32'd189928: dataIn1 = 32'd914
; 
32'd189929: dataIn1 = 32'd1660
; 
32'd189930: dataIn1 = 32'd1661
; 
32'd189931: dataIn1 = 32'd10350
; 
32'd189932: dataIn1 = 32'd10351
; 
32'd189933: dataIn1 = 32'd10352
; 
32'd189934: dataIn1 = 32'd434
; 
32'd189935: dataIn1 = 32'd911
; 
32'd189936: dataIn1 = 32'd1656
; 
32'd189937: dataIn1 = 32'd1661
; 
32'd189938: dataIn1 = 32'd10351
; 
32'd189939: dataIn1 = 32'd10352
; 
32'd189940: dataIn1 = 32'd10353
; 
32'd189941: dataIn1 = 32'd434
; 
32'd189942: dataIn1 = 32'd910
; 
32'd189943: dataIn1 = 32'd1656
; 
32'd189944: dataIn1 = 32'd1658
; 
32'd189945: dataIn1 = 32'd10352
; 
32'd189946: dataIn1 = 32'd10353
; 
32'd189947: dataIn1 = 32'd10354
; 
32'd189948: dataIn1 = 32'd910
; 
32'd189949: dataIn1 = 32'd912
; 
32'd189950: dataIn1 = 32'd1657
; 
32'd189951: dataIn1 = 32'd1658
; 
32'd189952: dataIn1 = 32'd10353
; 
32'd189953: dataIn1 = 32'd10354
; 
32'd189954: dataIn1 = 32'd10355
; 
32'd189955: dataIn1 = 32'd909
; 
32'd189956: dataIn1 = 32'd912
; 
32'd189957: dataIn1 = 32'd1657
; 
32'd189958: dataIn1 = 32'd1659
; 
32'd189959: dataIn1 = 32'd10354
; 
32'd189960: dataIn1 = 32'd10355
; 
32'd189961: dataIn1 = 32'd10356
; 
32'd189962: dataIn1 = 32'd238
; 
32'd189963: dataIn1 = 32'd909
; 
32'd189964: dataIn1 = 32'd1655
; 
32'd189965: dataIn1 = 32'd1659
; 
32'd189966: dataIn1 = 32'd10355
; 
32'd189967: dataIn1 = 32'd10356
; 
32'd189968: dataIn1 = 32'd10357
; 
32'd189969: dataIn1 = 32'd238
; 
32'd189970: dataIn1 = 32'd905
; 
32'd189971: dataIn1 = 32'd1650
; 
32'd189972: dataIn1 = 32'd1655
; 
32'd189973: dataIn1 = 32'd10356
; 
32'd189974: dataIn1 = 32'd10357
; 
32'd189975: dataIn1 = 32'd10358
; 
32'd189976: dataIn1 = 32'd905
; 
32'd189977: dataIn1 = 32'd906
; 
32'd189978: dataIn1 = 32'd1648
; 
32'd189979: dataIn1 = 32'd1650
; 
32'd189980: dataIn1 = 32'd10357
; 
32'd189981: dataIn1 = 32'd10358
; 
32'd189982: dataIn1 = 32'd10359
; 
32'd189983: dataIn1 = 32'd903
; 
32'd189984: dataIn1 = 32'd906
; 
32'd189985: dataIn1 = 32'd1648
; 
32'd189986: dataIn1 = 32'd1649
; 
32'd189987: dataIn1 = 32'd10358
; 
32'd189988: dataIn1 = 32'd10359
; 
32'd189989: dataIn1 = 32'd10360
; 
32'd189990: dataIn1 = 32'd433
; 
32'd189991: dataIn1 = 32'd903
; 
32'd189992: dataIn1 = 32'd1647
; 
32'd189993: dataIn1 = 32'd1649
; 
32'd189994: dataIn1 = 32'd10359
; 
32'd189995: dataIn1 = 32'd10360
; 
32'd189996: dataIn1 = 32'd10361
; 
32'd189997: dataIn1 = 32'd433
; 
32'd189998: dataIn1 = 32'd904
; 
32'd189999: dataIn1 = 32'd1647
; 
32'd190000: dataIn1 = 32'd1652
; 
32'd190001: dataIn1 = 32'd10360
; 
32'd190002: dataIn1 = 32'd10361
; 
32'd190003: dataIn1 = 32'd10362
; 
32'd190004: dataIn1 = 32'd904
; 
32'd190005: dataIn1 = 32'd908
; 
32'd190006: dataIn1 = 32'd1651
; 
32'd190007: dataIn1 = 32'd1652
; 
32'd190008: dataIn1 = 32'd10361
; 
32'd190009: dataIn1 = 32'd10362
; 
32'd190010: dataIn1 = 32'd10363
; 
32'd190011: dataIn1 = 32'd907
; 
32'd190012: dataIn1 = 32'd908
; 
32'd190013: dataIn1 = 32'd1651
; 
32'd190014: dataIn1 = 32'd1653
; 
32'd190015: dataIn1 = 32'd10362
; 
32'd190016: dataIn1 = 32'd10363
; 
32'd190017: dataIn1 = 32'd10364
; 
32'd190018: dataIn1 = 32'd237
; 
32'd190019: dataIn1 = 32'd907
; 
32'd190020: dataIn1 = 32'd1653
; 
32'd190021: dataIn1 = 32'd1654
; 
32'd190022: dataIn1 = 32'd10363
; 
32'd190023: dataIn1 = 32'd10364
; 
32'd190024: dataIn1 = 32'd10365
; 
32'd190025: dataIn1 = 32'd237
; 
32'd190026: dataIn1 = 32'd896
; 
32'd190027: dataIn1 = 32'd1637
; 
32'd190028: dataIn1 = 32'd1654
; 
32'd190029: dataIn1 = 32'd10364
; 
32'd190030: dataIn1 = 32'd10365
; 
32'd190031: dataIn1 = 32'd10366
; 
32'd190032: dataIn1 = 32'd895
; 
32'd190033: dataIn1 = 32'd896
; 
32'd190034: dataIn1 = 32'd1635
; 
32'd190035: dataIn1 = 32'd1637
; 
32'd190036: dataIn1 = 32'd10365
; 
32'd190037: dataIn1 = 32'd10366
; 
32'd190038: dataIn1 = 32'd10367
; 
32'd190039: dataIn1 = 32'd892
; 
32'd190040: dataIn1 = 32'd895
; 
32'd190041: dataIn1 = 32'd1635
; 
32'd190042: dataIn1 = 32'd1636
; 
32'd190043: dataIn1 = 32'd10366
; 
32'd190044: dataIn1 = 32'd10367
; 
32'd190045: dataIn1 = 32'd10368
; 
32'd190046: dataIn1 = 32'd431
; 
32'd190047: dataIn1 = 32'd892
; 
32'd190048: dataIn1 = 32'd1631
; 
32'd190049: dataIn1 = 32'd1636
; 
32'd190050: dataIn1 = 32'd10367
; 
32'd190051: dataIn1 = 32'd10368
; 
32'd190052: dataIn1 = 32'd10369
; 
32'd190053: dataIn1 = 32'd431
; 
32'd190054: dataIn1 = 32'd891
; 
32'd190055: dataIn1 = 32'd1631
; 
32'd190056: dataIn1 = 32'd1634
; 
32'd190057: dataIn1 = 32'd10368
; 
32'd190058: dataIn1 = 32'd10369
; 
32'd190059: dataIn1 = 32'd10370
; 
32'd190060: dataIn1 = 32'd891
; 
32'd190061: dataIn1 = 32'd894
; 
32'd190062: dataIn1 = 32'd1632
; 
32'd190063: dataIn1 = 32'd1634
; 
32'd190064: dataIn1 = 32'd10369
; 
32'd190065: dataIn1 = 32'd10370
; 
32'd190066: dataIn1 = 32'd10371
; 
32'd190067: dataIn1 = 32'd893
; 
32'd190068: dataIn1 = 32'd894
; 
32'd190069: dataIn1 = 32'd1632
; 
32'd190070: dataIn1 = 32'd1633
; 
32'd190071: dataIn1 = 32'd10370
; 
32'd190072: dataIn1 = 32'd10371
; 
32'd190073: dataIn1 = 32'd10372
; 
32'd190074: dataIn1 = 32'd235
; 
32'd190075: dataIn1 = 32'd893
; 
32'd190076: dataIn1 = 32'd1633
; 
32'd190077: dataIn1 = 32'd1646
; 
32'd190078: dataIn1 = 32'd10371
; 
32'd190079: dataIn1 = 32'd10372
; 
32'd190080: dataIn1 = 32'd10373
; 
32'd190081: dataIn1 = 32'd235
; 
32'd190082: dataIn1 = 32'd900
; 
32'd190083: dataIn1 = 32'd1640
; 
32'd190084: dataIn1 = 32'd1646
; 
32'd190085: dataIn1 = 32'd10372
; 
32'd190086: dataIn1 = 32'd10373
; 
32'd190087: dataIn1 = 32'd10374
; 
32'd190088: dataIn1 = 32'd899
; 
32'd190089: dataIn1 = 32'd900
; 
32'd190090: dataIn1 = 32'd1639
; 
32'd190091: dataIn1 = 32'd1640
; 
32'd190092: dataIn1 = 32'd10373
; 
32'd190093: dataIn1 = 32'd10374
; 
32'd190094: dataIn1 = 32'd10375
; 
32'd190095: dataIn1 = 32'd897
; 
32'd190096: dataIn1 = 32'd899
; 
32'd190097: dataIn1 = 32'd1639
; 
32'd190098: dataIn1 = 32'd1641
; 
32'd190099: dataIn1 = 32'd10374
; 
32'd190100: dataIn1 = 32'd10375
; 
32'd190101: dataIn1 = 32'd10376
; 
32'd190102: dataIn1 = 32'd432
; 
32'd190103: dataIn1 = 32'd897
; 
32'd190104: dataIn1 = 32'd1638
; 
32'd190105: dataIn1 = 32'd1641
; 
32'd190106: dataIn1 = 32'd10375
; 
32'd190107: dataIn1 = 32'd10376
; 
32'd190108: dataIn1 = 32'd10377
; 
32'd190109: dataIn1 = 32'd432
; 
32'd190110: dataIn1 = 32'd898
; 
32'd190111: dataIn1 = 32'd1638
; 
32'd190112: dataIn1 = 32'd1644
; 
32'd190113: dataIn1 = 32'd10376
; 
32'd190114: dataIn1 = 32'd10377
; 
32'd190115: dataIn1 = 32'd10378
; 
32'd190116: dataIn1 = 32'd898
; 
32'd190117: dataIn1 = 32'd901
; 
32'd190118: dataIn1 = 32'd1642
; 
32'd190119: dataIn1 = 32'd1644
; 
32'd190120: dataIn1 = 32'd10377
; 
32'd190121: dataIn1 = 32'd10378
; 
32'd190122: dataIn1 = 32'd10379
; 
32'd190123: dataIn1 = 32'd901
; 
32'd190124: dataIn1 = 32'd902
; 
32'd190125: dataIn1 = 32'd1642
; 
32'd190126: dataIn1 = 32'd1643
; 
32'd190127: dataIn1 = 32'd10378
; 
32'd190128: dataIn1 = 32'd10379
; 
32'd190129: dataIn1 = 32'd10380
; 
32'd190130: dataIn1 = 32'd234
; 
32'd190131: dataIn1 = 32'd902
; 
32'd190132: dataIn1 = 32'd1643
; 
32'd190133: dataIn1 = 32'd1645
; 
32'd190134: dataIn1 = 32'd10379
; 
32'd190135: dataIn1 = 32'd10380
; 
32'd190136: dataIn1 = 32'd10381
; 
32'd190137: dataIn1 = 32'd234
; 
32'd190138: dataIn1 = 32'd889
; 
32'd190139: dataIn1 = 32'd1630
; 
32'd190140: dataIn1 = 32'd1645
; 
32'd190141: dataIn1 = 32'd10380
; 
32'd190142: dataIn1 = 32'd10381
; 
32'd190143: dataIn1 = 32'd10382
; 
32'd190144: dataIn1 = 32'd889
; 
32'd190145: dataIn1 = 32'd890
; 
32'd190146: dataIn1 = 32'd1628
; 
32'd190147: dataIn1 = 32'd1630
; 
32'd190148: dataIn1 = 32'd10381
; 
32'd190149: dataIn1 = 32'd10382
; 
32'd190150: dataIn1 = 32'd10383
; 
32'd190151: dataIn1 = 32'd887
; 
32'd190152: dataIn1 = 32'd890
; 
32'd190153: dataIn1 = 32'd1628
; 
32'd190154: dataIn1 = 32'd1629
; 
32'd190155: dataIn1 = 32'd10382
; 
32'd190156: dataIn1 = 32'd10383
; 
32'd190157: dataIn1 = 32'd10384
; 
32'd190158: dataIn1 = 32'd430
; 
32'd190159: dataIn1 = 32'd887
; 
32'd190160: dataIn1 = 32'd1624
; 
32'd190161: dataIn1 = 32'd1629
; 
32'd190162: dataIn1 = 32'd10383
; 
32'd190163: dataIn1 = 32'd10384
; 
32'd190164: dataIn1 = 32'd10385
; 
32'd190165: dataIn1 = 32'd430
; 
32'd190166: dataIn1 = 32'd886
; 
32'd190167: dataIn1 = 32'd1624
; 
32'd190168: dataIn1 = 32'd1626
; 
32'd190169: dataIn1 = 32'd10384
; 
32'd190170: dataIn1 = 32'd10385
; 
32'd190171: dataIn1 = 32'd10386
; 
32'd190172: dataIn1 = 32'd886
; 
32'd190173: dataIn1 = 32'd888
; 
32'd190174: dataIn1 = 32'd1625
; 
32'd190175: dataIn1 = 32'd1626
; 
32'd190176: dataIn1 = 32'd10385
; 
32'd190177: dataIn1 = 32'd10386
; 
32'd190178: dataIn1 = 32'd10387
; 
32'd190179: dataIn1 = 32'd885
; 
32'd190180: dataIn1 = 32'd888
; 
32'd190181: dataIn1 = 32'd1625
; 
32'd190182: dataIn1 = 32'd1627
; 
32'd190183: dataIn1 = 32'd10386
; 
32'd190184: dataIn1 = 32'd10387
; 
32'd190185: dataIn1 = 32'd10388
; 
32'd190186: dataIn1 = 32'd232
; 
32'd190187: dataIn1 = 32'd885
; 
32'd190188: dataIn1 = 32'd1623
; 
32'd190189: dataIn1 = 32'd1627
; 
32'd190190: dataIn1 = 32'd10387
; 
32'd190191: dataIn1 = 32'd10388
; 
32'd190192: dataIn1 = 32'd10389
; 
32'd190193: dataIn1 = 32'd232
; 
32'd190194: dataIn1 = 32'd881
; 
32'd190195: dataIn1 = 32'd1618
; 
32'd190196: dataIn1 = 32'd1623
; 
32'd190197: dataIn1 = 32'd10388
; 
32'd190198: dataIn1 = 32'd10389
; 
32'd190199: dataIn1 = 32'd10390
; 
32'd190200: dataIn1 = 32'd881
; 
32'd190201: dataIn1 = 32'd882
; 
32'd190202: dataIn1 = 32'd1616
; 
32'd190203: dataIn1 = 32'd1618
; 
32'd190204: dataIn1 = 32'd10389
; 
32'd190205: dataIn1 = 32'd10390
; 
32'd190206: dataIn1 = 32'd10391
; 
32'd190207: dataIn1 = 32'd879
; 
32'd190208: dataIn1 = 32'd882
; 
32'd190209: dataIn1 = 32'd1616
; 
32'd190210: dataIn1 = 32'd1617
; 
32'd190211: dataIn1 = 32'd10390
; 
32'd190212: dataIn1 = 32'd10391
; 
32'd190213: dataIn1 = 32'd10392
; 
32'd190214: dataIn1 = 32'd429
; 
32'd190215: dataIn1 = 32'd879
; 
32'd190216: dataIn1 = 32'd1615
; 
32'd190217: dataIn1 = 32'd1617
; 
32'd190218: dataIn1 = 32'd10391
; 
32'd190219: dataIn1 = 32'd10392
; 
32'd190220: dataIn1 = 32'd10393
; 
32'd190221: dataIn1 = 32'd429
; 
32'd190222: dataIn1 = 32'd880
; 
32'd190223: dataIn1 = 32'd1615
; 
32'd190224: dataIn1 = 32'd1620
; 
32'd190225: dataIn1 = 32'd10392
; 
32'd190226: dataIn1 = 32'd10393
; 
32'd190227: dataIn1 = 32'd10394
; 
32'd190228: dataIn1 = 32'd880
; 
32'd190229: dataIn1 = 32'd884
; 
32'd190230: dataIn1 = 32'd1619
; 
32'd190231: dataIn1 = 32'd1620
; 
32'd190232: dataIn1 = 32'd10393
; 
32'd190233: dataIn1 = 32'd10394
; 
32'd190234: dataIn1 = 32'd10395
; 
32'd190235: dataIn1 = 32'd883
; 
32'd190236: dataIn1 = 32'd884
; 
32'd190237: dataIn1 = 32'd1619
; 
32'd190238: dataIn1 = 32'd1621
; 
32'd190239: dataIn1 = 32'd10394
; 
32'd190240: dataIn1 = 32'd10395
; 
32'd190241: dataIn1 = 32'd10396
; 
32'd190242: dataIn1 = 32'd231
; 
32'd190243: dataIn1 = 32'd883
; 
32'd190244: dataIn1 = 32'd1621
; 
32'd190245: dataIn1 = 32'd1622
; 
32'd190246: dataIn1 = 32'd10395
; 
32'd190247: dataIn1 = 32'd10396
; 
32'd190248: dataIn1 = 32'd10397
; 
32'd190249: dataIn1 = 32'd231
; 
32'd190250: dataIn1 = 32'd872
; 
32'd190251: dataIn1 = 32'd1605
; 
32'd190252: dataIn1 = 32'd1622
; 
32'd190253: dataIn1 = 32'd10396
; 
32'd190254: dataIn1 = 32'd10397
; 
32'd190255: dataIn1 = 32'd10398
; 
32'd190256: dataIn1 = 32'd871
; 
32'd190257: dataIn1 = 32'd872
; 
32'd190258: dataIn1 = 32'd1603
; 
32'd190259: dataIn1 = 32'd1605
; 
32'd190260: dataIn1 = 32'd10397
; 
32'd190261: dataIn1 = 32'd10398
; 
32'd190262: dataIn1 = 32'd10399
; 
32'd190263: dataIn1 = 32'd868
; 
32'd190264: dataIn1 = 32'd871
; 
32'd190265: dataIn1 = 32'd1603
; 
32'd190266: dataIn1 = 32'd1604
; 
32'd190267: dataIn1 = 32'd10398
; 
32'd190268: dataIn1 = 32'd10399
; 
32'd190269: dataIn1 = 32'd10400
; 
32'd190270: dataIn1 = 32'd427
; 
32'd190271: dataIn1 = 32'd868
; 
32'd190272: dataIn1 = 32'd1599
; 
32'd190273: dataIn1 = 32'd1604
; 
32'd190274: dataIn1 = 32'd10399
; 
32'd190275: dataIn1 = 32'd10400
; 
32'd190276: dataIn1 = 32'd10401
; 
32'd190277: dataIn1 = 32'd427
; 
32'd190278: dataIn1 = 32'd867
; 
32'd190279: dataIn1 = 32'd1599
; 
32'd190280: dataIn1 = 32'd1602
; 
32'd190281: dataIn1 = 32'd10400
; 
32'd190282: dataIn1 = 32'd10401
; 
32'd190283: dataIn1 = 32'd10402
; 
32'd190284: dataIn1 = 32'd867
; 
32'd190285: dataIn1 = 32'd870
; 
32'd190286: dataIn1 = 32'd1600
; 
32'd190287: dataIn1 = 32'd1602
; 
32'd190288: dataIn1 = 32'd10401
; 
32'd190289: dataIn1 = 32'd10402
; 
32'd190290: dataIn1 = 32'd10403
; 
32'd190291: dataIn1 = 32'd869
; 
32'd190292: dataIn1 = 32'd870
; 
32'd190293: dataIn1 = 32'd1600
; 
32'd190294: dataIn1 = 32'd1601
; 
32'd190295: dataIn1 = 32'd10402
; 
32'd190296: dataIn1 = 32'd10403
; 
32'd190297: dataIn1 = 32'd10404
; 
32'd190298: dataIn1 = 32'd229
; 
32'd190299: dataIn1 = 32'd869
; 
32'd190300: dataIn1 = 32'd1601
; 
32'd190301: dataIn1 = 32'd1614
; 
32'd190302: dataIn1 = 32'd10403
; 
32'd190303: dataIn1 = 32'd10404
; 
32'd190304: dataIn1 = 32'd10405
; 
32'd190305: dataIn1 = 32'd229
; 
32'd190306: dataIn1 = 32'd876
; 
32'd190307: dataIn1 = 32'd1608
; 
32'd190308: dataIn1 = 32'd1614
; 
32'd190309: dataIn1 = 32'd10404
; 
32'd190310: dataIn1 = 32'd10405
; 
32'd190311: dataIn1 = 32'd10406
; 
32'd190312: dataIn1 = 32'd875
; 
32'd190313: dataIn1 = 32'd876
; 
32'd190314: dataIn1 = 32'd1607
; 
32'd190315: dataIn1 = 32'd1608
; 
32'd190316: dataIn1 = 32'd10405
; 
32'd190317: dataIn1 = 32'd10406
; 
32'd190318: dataIn1 = 32'd10407
; 
32'd190319: dataIn1 = 32'd873
; 
32'd190320: dataIn1 = 32'd875
; 
32'd190321: dataIn1 = 32'd1607
; 
32'd190322: dataIn1 = 32'd1609
; 
32'd190323: dataIn1 = 32'd10406
; 
32'd190324: dataIn1 = 32'd10407
; 
32'd190325: dataIn1 = 32'd10408
; 
32'd190326: dataIn1 = 32'd428
; 
32'd190327: dataIn1 = 32'd873
; 
32'd190328: dataIn1 = 32'd1606
; 
32'd190329: dataIn1 = 32'd1609
; 
32'd190330: dataIn1 = 32'd10407
; 
32'd190331: dataIn1 = 32'd10408
; 
32'd190332: dataIn1 = 32'd10409
; 
32'd190333: dataIn1 = 32'd428
; 
32'd190334: dataIn1 = 32'd874
; 
32'd190335: dataIn1 = 32'd1606
; 
32'd190336: dataIn1 = 32'd1612
; 
32'd190337: dataIn1 = 32'd10408
; 
32'd190338: dataIn1 = 32'd10409
; 
32'd190339: dataIn1 = 32'd10410
; 
32'd190340: dataIn1 = 32'd874
; 
32'd190341: dataIn1 = 32'd877
; 
32'd190342: dataIn1 = 32'd1610
; 
32'd190343: dataIn1 = 32'd1612
; 
32'd190344: dataIn1 = 32'd10409
; 
32'd190345: dataIn1 = 32'd10410
; 
32'd190346: dataIn1 = 32'd10411
; 
32'd190347: dataIn1 = 32'd877
; 
32'd190348: dataIn1 = 32'd878
; 
32'd190349: dataIn1 = 32'd1610
; 
32'd190350: dataIn1 = 32'd1611
; 
32'd190351: dataIn1 = 32'd10410
; 
32'd190352: dataIn1 = 32'd10411
; 
32'd190353: dataIn1 = 32'd10412
; 
32'd190354: dataIn1 = 32'd228
; 
32'd190355: dataIn1 = 32'd878
; 
32'd190356: dataIn1 = 32'd1611
; 
32'd190357: dataIn1 = 32'd1613
; 
32'd190358: dataIn1 = 32'd10411
; 
32'd190359: dataIn1 = 32'd10412
; 
32'd190360: dataIn1 = 32'd10413
; 
32'd190361: dataIn1 = 32'd228
; 
32'd190362: dataIn1 = 32'd865
; 
32'd190363: dataIn1 = 32'd1598
; 
32'd190364: dataIn1 = 32'd1613
; 
32'd190365: dataIn1 = 32'd10412
; 
32'd190366: dataIn1 = 32'd10413
; 
32'd190367: dataIn1 = 32'd10414
; 
32'd190368: dataIn1 = 32'd865
; 
32'd190369: dataIn1 = 32'd866
; 
32'd190370: dataIn1 = 32'd1596
; 
32'd190371: dataIn1 = 32'd1598
; 
32'd190372: dataIn1 = 32'd10413
; 
32'd190373: dataIn1 = 32'd10414
; 
32'd190374: dataIn1 = 32'd10415
; 
32'd190375: dataIn1 = 32'd863
; 
32'd190376: dataIn1 = 32'd866
; 
32'd190377: dataIn1 = 32'd1596
; 
32'd190378: dataIn1 = 32'd1597
; 
32'd190379: dataIn1 = 32'd10414
; 
32'd190380: dataIn1 = 32'd10415
; 
32'd190381: dataIn1 = 32'd10416
; 
32'd190382: dataIn1 = 32'd426
; 
32'd190383: dataIn1 = 32'd863
; 
32'd190384: dataIn1 = 32'd1592
; 
32'd190385: dataIn1 = 32'd1597
; 
32'd190386: dataIn1 = 32'd10415
; 
32'd190387: dataIn1 = 32'd10416
; 
32'd190388: dataIn1 = 32'd10417
; 
32'd190389: dataIn1 = 32'd426
; 
32'd190390: dataIn1 = 32'd862
; 
32'd190391: dataIn1 = 32'd1592
; 
32'd190392: dataIn1 = 32'd1594
; 
32'd190393: dataIn1 = 32'd10416
; 
32'd190394: dataIn1 = 32'd10417
; 
32'd190395: dataIn1 = 32'd10418
; 
32'd190396: dataIn1 = 32'd862
; 
32'd190397: dataIn1 = 32'd864
; 
32'd190398: dataIn1 = 32'd1593
; 
32'd190399: dataIn1 = 32'd1594
; 
32'd190400: dataIn1 = 32'd10417
; 
32'd190401: dataIn1 = 32'd10418
; 
32'd190402: dataIn1 = 32'd10419
; 
32'd190403: dataIn1 = 32'd861
; 
32'd190404: dataIn1 = 32'd864
; 
32'd190405: dataIn1 = 32'd1593
; 
32'd190406: dataIn1 = 32'd1595
; 
32'd190407: dataIn1 = 32'd10418
; 
32'd190408: dataIn1 = 32'd10419
; 
32'd190409: dataIn1 = 32'd10420
; 
32'd190410: dataIn1 = 32'd226
; 
32'd190411: dataIn1 = 32'd861
; 
32'd190412: dataIn1 = 32'd1591
; 
32'd190413: dataIn1 = 32'd1595
; 
32'd190414: dataIn1 = 32'd10419
; 
32'd190415: dataIn1 = 32'd10420
; 
32'd190416: dataIn1 = 32'd10421
; 
32'd190417: dataIn1 = 32'd226
; 
32'd190418: dataIn1 = 32'd857
; 
32'd190419: dataIn1 = 32'd1586
; 
32'd190420: dataIn1 = 32'd1591
; 
32'd190421: dataIn1 = 32'd10420
; 
32'd190422: dataIn1 = 32'd10421
; 
32'd190423: dataIn1 = 32'd10422
; 
32'd190424: dataIn1 = 32'd857
; 
32'd190425: dataIn1 = 32'd858
; 
32'd190426: dataIn1 = 32'd1584
; 
32'd190427: dataIn1 = 32'd1586
; 
32'd190428: dataIn1 = 32'd10421
; 
32'd190429: dataIn1 = 32'd10422
; 
32'd190430: dataIn1 = 32'd10423
; 
32'd190431: dataIn1 = 32'd855
; 
32'd190432: dataIn1 = 32'd858
; 
32'd190433: dataIn1 = 32'd1584
; 
32'd190434: dataIn1 = 32'd1585
; 
32'd190435: dataIn1 = 32'd10422
; 
32'd190436: dataIn1 = 32'd10423
; 
32'd190437: dataIn1 = 32'd10424
; 
32'd190438: dataIn1 = 32'd425
; 
32'd190439: dataIn1 = 32'd855
; 
32'd190440: dataIn1 = 32'd1583
; 
32'd190441: dataIn1 = 32'd1585
; 
32'd190442: dataIn1 = 32'd10423
; 
32'd190443: dataIn1 = 32'd10424
; 
32'd190444: dataIn1 = 32'd10425
; 
32'd190445: dataIn1 = 32'd425
; 
32'd190446: dataIn1 = 32'd856
; 
32'd190447: dataIn1 = 32'd1583
; 
32'd190448: dataIn1 = 32'd1588
; 
32'd190449: dataIn1 = 32'd10424
; 
32'd190450: dataIn1 = 32'd10425
; 
32'd190451: dataIn1 = 32'd10426
; 
32'd190452: dataIn1 = 32'd856
; 
32'd190453: dataIn1 = 32'd860
; 
32'd190454: dataIn1 = 32'd1587
; 
32'd190455: dataIn1 = 32'd1588
; 
32'd190456: dataIn1 = 32'd10425
; 
32'd190457: dataIn1 = 32'd10426
; 
32'd190458: dataIn1 = 32'd10427
; 
32'd190459: dataIn1 = 32'd859
; 
32'd190460: dataIn1 = 32'd860
; 
32'd190461: dataIn1 = 32'd1587
; 
32'd190462: dataIn1 = 32'd1589
; 
32'd190463: dataIn1 = 32'd10426
; 
32'd190464: dataIn1 = 32'd10427
; 
32'd190465: dataIn1 = 32'd10428
; 
32'd190466: dataIn1 = 32'd225
; 
32'd190467: dataIn1 = 32'd859
; 
32'd190468: dataIn1 = 32'd1589
; 
32'd190469: dataIn1 = 32'd1590
; 
32'd190470: dataIn1 = 32'd10427
; 
32'd190471: dataIn1 = 32'd10428
; 
32'd190472: dataIn1 = 32'd10429
; 
32'd190473: dataIn1 = 32'd225
; 
32'd190474: dataIn1 = 32'd848
; 
32'd190475: dataIn1 = 32'd1573
; 
32'd190476: dataIn1 = 32'd1590
; 
32'd190477: dataIn1 = 32'd10428
; 
32'd190478: dataIn1 = 32'd10429
; 
32'd190479: dataIn1 = 32'd10430
; 
32'd190480: dataIn1 = 32'd847
; 
32'd190481: dataIn1 = 32'd848
; 
32'd190482: dataIn1 = 32'd1571
; 
32'd190483: dataIn1 = 32'd1573
; 
32'd190484: dataIn1 = 32'd10429
; 
32'd190485: dataIn1 = 32'd10430
; 
32'd190486: dataIn1 = 32'd10431
; 
32'd190487: dataIn1 = 32'd844
; 
32'd190488: dataIn1 = 32'd847
; 
32'd190489: dataIn1 = 32'd1571
; 
32'd190490: dataIn1 = 32'd1572
; 
32'd190491: dataIn1 = 32'd10430
; 
32'd190492: dataIn1 = 32'd10431
; 
32'd190493: dataIn1 = 32'd10432
; 
32'd190494: dataIn1 = 32'd423
; 
32'd190495: dataIn1 = 32'd844
; 
32'd190496: dataIn1 = 32'd1567
; 
32'd190497: dataIn1 = 32'd1572
; 
32'd190498: dataIn1 = 32'd10431
; 
32'd190499: dataIn1 = 32'd10432
; 
32'd190500: dataIn1 = 32'd10433
; 
32'd190501: dataIn1 = 32'd423
; 
32'd190502: dataIn1 = 32'd843
; 
32'd190503: dataIn1 = 32'd1567
; 
32'd190504: dataIn1 = 32'd1570
; 
32'd190505: dataIn1 = 32'd10432
; 
32'd190506: dataIn1 = 32'd10433
; 
32'd190507: dataIn1 = 32'd10434
; 
32'd190508: dataIn1 = 32'd843
; 
32'd190509: dataIn1 = 32'd846
; 
32'd190510: dataIn1 = 32'd1568
; 
32'd190511: dataIn1 = 32'd1570
; 
32'd190512: dataIn1 = 32'd10433
; 
32'd190513: dataIn1 = 32'd10434
; 
32'd190514: dataIn1 = 32'd10435
; 
32'd190515: dataIn1 = 32'd845
; 
32'd190516: dataIn1 = 32'd846
; 
32'd190517: dataIn1 = 32'd1568
; 
32'd190518: dataIn1 = 32'd1569
; 
32'd190519: dataIn1 = 32'd10434
; 
32'd190520: dataIn1 = 32'd10435
; 
32'd190521: dataIn1 = 32'd10436
; 
32'd190522: dataIn1 = 32'd223
; 
32'd190523: dataIn1 = 32'd845
; 
32'd190524: dataIn1 = 32'd1569
; 
32'd190525: dataIn1 = 32'd1582
; 
32'd190526: dataIn1 = 32'd10435
; 
32'd190527: dataIn1 = 32'd10436
; 
32'd190528: dataIn1 = 32'd10437
; 
32'd190529: dataIn1 = 32'd223
; 
32'd190530: dataIn1 = 32'd852
; 
32'd190531: dataIn1 = 32'd1576
; 
32'd190532: dataIn1 = 32'd1582
; 
32'd190533: dataIn1 = 32'd10436
; 
32'd190534: dataIn1 = 32'd10437
; 
32'd190535: dataIn1 = 32'd10438
; 
32'd190536: dataIn1 = 32'd851
; 
32'd190537: dataIn1 = 32'd852
; 
32'd190538: dataIn1 = 32'd1575
; 
32'd190539: dataIn1 = 32'd1576
; 
32'd190540: dataIn1 = 32'd10437
; 
32'd190541: dataIn1 = 32'd10438
; 
32'd190542: dataIn1 = 32'd10439
; 
32'd190543: dataIn1 = 32'd849
; 
32'd190544: dataIn1 = 32'd851
; 
32'd190545: dataIn1 = 32'd1575
; 
32'd190546: dataIn1 = 32'd1577
; 
32'd190547: dataIn1 = 32'd10438
; 
32'd190548: dataIn1 = 32'd10439
; 
32'd190549: dataIn1 = 32'd10440
; 
32'd190550: dataIn1 = 32'd424
; 
32'd190551: dataIn1 = 32'd849
; 
32'd190552: dataIn1 = 32'd1574
; 
32'd190553: dataIn1 = 32'd1577
; 
32'd190554: dataIn1 = 32'd10439
; 
32'd190555: dataIn1 = 32'd10440
; 
32'd190556: dataIn1 = 32'd10441
; 
32'd190557: dataIn1 = 32'd424
; 
32'd190558: dataIn1 = 32'd850
; 
32'd190559: dataIn1 = 32'd1574
; 
32'd190560: dataIn1 = 32'd1580
; 
32'd190561: dataIn1 = 32'd10440
; 
32'd190562: dataIn1 = 32'd10441
; 
32'd190563: dataIn1 = 32'd10442
; 
32'd190564: dataIn1 = 32'd850
; 
32'd190565: dataIn1 = 32'd853
; 
32'd190566: dataIn1 = 32'd1578
; 
32'd190567: dataIn1 = 32'd1580
; 
32'd190568: dataIn1 = 32'd10441
; 
32'd190569: dataIn1 = 32'd10442
; 
32'd190570: dataIn1 = 32'd10443
; 
32'd190571: dataIn1 = 32'd853
; 
32'd190572: dataIn1 = 32'd854
; 
32'd190573: dataIn1 = 32'd1578
; 
32'd190574: dataIn1 = 32'd1579
; 
32'd190575: dataIn1 = 32'd10442
; 
32'd190576: dataIn1 = 32'd10443
; 
32'd190577: dataIn1 = 32'd10444
; 
32'd190578: dataIn1 = 32'd222
; 
32'd190579: dataIn1 = 32'd854
; 
32'd190580: dataIn1 = 32'd1579
; 
32'd190581: dataIn1 = 32'd1581
; 
32'd190582: dataIn1 = 32'd10443
; 
32'd190583: dataIn1 = 32'd10444
; 
32'd190584: dataIn1 = 32'd10445
; 
32'd190585: dataIn1 = 32'd222
; 
32'd190586: dataIn1 = 32'd841
; 
32'd190587: dataIn1 = 32'd1566
; 
32'd190588: dataIn1 = 32'd1581
; 
32'd190589: dataIn1 = 32'd10444
; 
32'd190590: dataIn1 = 32'd10445
; 
32'd190591: dataIn1 = 32'd10446
; 
32'd190592: dataIn1 = 32'd841
; 
32'd190593: dataIn1 = 32'd842
; 
32'd190594: dataIn1 = 32'd1564
; 
32'd190595: dataIn1 = 32'd1566
; 
32'd190596: dataIn1 = 32'd10445
; 
32'd190597: dataIn1 = 32'd10446
; 
32'd190598: dataIn1 = 32'd10447
; 
32'd190599: dataIn1 = 32'd839
; 
32'd190600: dataIn1 = 32'd842
; 
32'd190601: dataIn1 = 32'd1564
; 
32'd190602: dataIn1 = 32'd1565
; 
32'd190603: dataIn1 = 32'd10446
; 
32'd190604: dataIn1 = 32'd10447
; 
32'd190605: dataIn1 = 32'd10448
; 
32'd190606: dataIn1 = 32'd422
; 
32'd190607: dataIn1 = 32'd839
; 
32'd190608: dataIn1 = 32'd1560
; 
32'd190609: dataIn1 = 32'd1565
; 
32'd190610: dataIn1 = 32'd10447
; 
32'd190611: dataIn1 = 32'd10448
; 
32'd190612: dataIn1 = 32'd10449
; 
32'd190613: dataIn1 = 32'd422
; 
32'd190614: dataIn1 = 32'd838
; 
32'd190615: dataIn1 = 32'd1560
; 
32'd190616: dataIn1 = 32'd1562
; 
32'd190617: dataIn1 = 32'd10448
; 
32'd190618: dataIn1 = 32'd10449
; 
32'd190619: dataIn1 = 32'd10450
; 
32'd190620: dataIn1 = 32'd838
; 
32'd190621: dataIn1 = 32'd840
; 
32'd190622: dataIn1 = 32'd1561
; 
32'd190623: dataIn1 = 32'd1562
; 
32'd190624: dataIn1 = 32'd10449
; 
32'd190625: dataIn1 = 32'd10450
; 
32'd190626: dataIn1 = 32'd10451
; 
32'd190627: dataIn1 = 32'd837
; 
32'd190628: dataIn1 = 32'd840
; 
32'd190629: dataIn1 = 32'd1561
; 
32'd190630: dataIn1 = 32'd1563
; 
32'd190631: dataIn1 = 32'd10450
; 
32'd190632: dataIn1 = 32'd10451
; 
32'd190633: dataIn1 = 32'd10452
; 
32'd190634: dataIn1 = 32'd220
; 
32'd190635: dataIn1 = 32'd837
; 
32'd190636: dataIn1 = 32'd1559
; 
32'd190637: dataIn1 = 32'd1563
; 
32'd190638: dataIn1 = 32'd10451
; 
32'd190639: dataIn1 = 32'd10452
; 
32'd190640: dataIn1 = 32'd10453
; 
32'd190641: dataIn1 = 32'd220
; 
32'd190642: dataIn1 = 32'd833
; 
32'd190643: dataIn1 = 32'd1554
; 
32'd190644: dataIn1 = 32'd1559
; 
32'd190645: dataIn1 = 32'd10452
; 
32'd190646: dataIn1 = 32'd10453
; 
32'd190647: dataIn1 = 32'd10454
; 
32'd190648: dataIn1 = 32'd833
; 
32'd190649: dataIn1 = 32'd834
; 
32'd190650: dataIn1 = 32'd1552
; 
32'd190651: dataIn1 = 32'd1554
; 
32'd190652: dataIn1 = 32'd10453
; 
32'd190653: dataIn1 = 32'd10454
; 
32'd190654: dataIn1 = 32'd10455
; 
32'd190655: dataIn1 = 32'd831
; 
32'd190656: dataIn1 = 32'd834
; 
32'd190657: dataIn1 = 32'd1552
; 
32'd190658: dataIn1 = 32'd1553
; 
32'd190659: dataIn1 = 32'd10454
; 
32'd190660: dataIn1 = 32'd10455
; 
32'd190661: dataIn1 = 32'd10456
; 
32'd190662: dataIn1 = 32'd421
; 
32'd190663: dataIn1 = 32'd831
; 
32'd190664: dataIn1 = 32'd1551
; 
32'd190665: dataIn1 = 32'd1553
; 
32'd190666: dataIn1 = 32'd10455
; 
32'd190667: dataIn1 = 32'd10456
; 
32'd190668: dataIn1 = 32'd10457
; 
32'd190669: dataIn1 = 32'd421
; 
32'd190670: dataIn1 = 32'd832
; 
32'd190671: dataIn1 = 32'd1551
; 
32'd190672: dataIn1 = 32'd1556
; 
32'd190673: dataIn1 = 32'd10456
; 
32'd190674: dataIn1 = 32'd10457
; 
32'd190675: dataIn1 = 32'd10458
; 
32'd190676: dataIn1 = 32'd832
; 
32'd190677: dataIn1 = 32'd836
; 
32'd190678: dataIn1 = 32'd1555
; 
32'd190679: dataIn1 = 32'd1556
; 
32'd190680: dataIn1 = 32'd10457
; 
32'd190681: dataIn1 = 32'd10458
; 
32'd190682: dataIn1 = 32'd10459
; 
32'd190683: dataIn1 = 32'd835
; 
32'd190684: dataIn1 = 32'd836
; 
32'd190685: dataIn1 = 32'd1555
; 
32'd190686: dataIn1 = 32'd1557
; 
32'd190687: dataIn1 = 32'd10458
; 
32'd190688: dataIn1 = 32'd10459
; 
32'd190689: dataIn1 = 32'd10460
; 
32'd190690: dataIn1 = 32'd219
; 
32'd190691: dataIn1 = 32'd835
; 
32'd190692: dataIn1 = 32'd1557
; 
32'd190693: dataIn1 = 32'd1558
; 
32'd190694: dataIn1 = 32'd10459
; 
32'd190695: dataIn1 = 32'd10460
; 
32'd190696: dataIn1 = 32'd10461
; 
32'd190697: dataIn1 = 32'd219
; 
32'd190698: dataIn1 = 32'd824
; 
32'd190699: dataIn1 = 32'd1541
; 
32'd190700: dataIn1 = 32'd1558
; 
32'd190701: dataIn1 = 32'd10460
; 
32'd190702: dataIn1 = 32'd10461
; 
32'd190703: dataIn1 = 32'd10462
; 
32'd190704: dataIn1 = 32'd823
; 
32'd190705: dataIn1 = 32'd824
; 
32'd190706: dataIn1 = 32'd1539
; 
32'd190707: dataIn1 = 32'd1541
; 
32'd190708: dataIn1 = 32'd10461
; 
32'd190709: dataIn1 = 32'd10462
; 
32'd190710: dataIn1 = 32'd10463
; 
32'd190711: dataIn1 = 32'd820
; 
32'd190712: dataIn1 = 32'd823
; 
32'd190713: dataIn1 = 32'd1539
; 
32'd190714: dataIn1 = 32'd1540
; 
32'd190715: dataIn1 = 32'd10462
; 
32'd190716: dataIn1 = 32'd10463
; 
32'd190717: dataIn1 = 32'd10464
; 
32'd190718: dataIn1 = 32'd419
; 
32'd190719: dataIn1 = 32'd820
; 
32'd190720: dataIn1 = 32'd1535
; 
32'd190721: dataIn1 = 32'd1540
; 
32'd190722: dataIn1 = 32'd10463
; 
32'd190723: dataIn1 = 32'd10464
; 
32'd190724: dataIn1 = 32'd10465
; 
32'd190725: dataIn1 = 32'd419
; 
32'd190726: dataIn1 = 32'd819
; 
32'd190727: dataIn1 = 32'd1535
; 
32'd190728: dataIn1 = 32'd1538
; 
32'd190729: dataIn1 = 32'd10464
; 
32'd190730: dataIn1 = 32'd10465
; 
32'd190731: dataIn1 = 32'd10466
; 
32'd190732: dataIn1 = 32'd819
; 
32'd190733: dataIn1 = 32'd822
; 
32'd190734: dataIn1 = 32'd1536
; 
32'd190735: dataIn1 = 32'd1538
; 
32'd190736: dataIn1 = 32'd10465
; 
32'd190737: dataIn1 = 32'd10466
; 
32'd190738: dataIn1 = 32'd10467
; 
32'd190739: dataIn1 = 32'd821
; 
32'd190740: dataIn1 = 32'd822
; 
32'd190741: dataIn1 = 32'd1536
; 
32'd190742: dataIn1 = 32'd1537
; 
32'd190743: dataIn1 = 32'd10466
; 
32'd190744: dataIn1 = 32'd10467
; 
32'd190745: dataIn1 = 32'd10468
; 
32'd190746: dataIn1 = 32'd217
; 
32'd190747: dataIn1 = 32'd821
; 
32'd190748: dataIn1 = 32'd1537
; 
32'd190749: dataIn1 = 32'd1550
; 
32'd190750: dataIn1 = 32'd10467
; 
32'd190751: dataIn1 = 32'd10468
; 
32'd190752: dataIn1 = 32'd10469
; 
32'd190753: dataIn1 = 32'd217
; 
32'd190754: dataIn1 = 32'd828
; 
32'd190755: dataIn1 = 32'd1544
; 
32'd190756: dataIn1 = 32'd1550
; 
32'd190757: dataIn1 = 32'd10468
; 
32'd190758: dataIn1 = 32'd10469
; 
32'd190759: dataIn1 = 32'd10470
; 
32'd190760: dataIn1 = 32'd827
; 
32'd190761: dataIn1 = 32'd828
; 
32'd190762: dataIn1 = 32'd1543
; 
32'd190763: dataIn1 = 32'd1544
; 
32'd190764: dataIn1 = 32'd10469
; 
32'd190765: dataIn1 = 32'd10470
; 
32'd190766: dataIn1 = 32'd10471
; 
32'd190767: dataIn1 = 32'd825
; 
32'd190768: dataIn1 = 32'd827
; 
32'd190769: dataIn1 = 32'd1543
; 
32'd190770: dataIn1 = 32'd1545
; 
32'd190771: dataIn1 = 32'd10470
; 
32'd190772: dataIn1 = 32'd10471
; 
32'd190773: dataIn1 = 32'd10472
; 
32'd190774: dataIn1 = 32'd420
; 
32'd190775: dataIn1 = 32'd825
; 
32'd190776: dataIn1 = 32'd1542
; 
32'd190777: dataIn1 = 32'd1545
; 
32'd190778: dataIn1 = 32'd10471
; 
32'd190779: dataIn1 = 32'd10472
; 
32'd190780: dataIn1 = 32'd10473
; 
32'd190781: dataIn1 = 32'd420
; 
32'd190782: dataIn1 = 32'd826
; 
32'd190783: dataIn1 = 32'd1542
; 
32'd190784: dataIn1 = 32'd1548
; 
32'd190785: dataIn1 = 32'd10472
; 
32'd190786: dataIn1 = 32'd10473
; 
32'd190787: dataIn1 = 32'd10474
; 
32'd190788: dataIn1 = 32'd826
; 
32'd190789: dataIn1 = 32'd829
; 
32'd190790: dataIn1 = 32'd1546
; 
32'd190791: dataIn1 = 32'd1548
; 
32'd190792: dataIn1 = 32'd10473
; 
32'd190793: dataIn1 = 32'd10474
; 
32'd190794: dataIn1 = 32'd10475
; 
32'd190795: dataIn1 = 32'd829
; 
32'd190796: dataIn1 = 32'd830
; 
32'd190797: dataIn1 = 32'd1546
; 
32'd190798: dataIn1 = 32'd1547
; 
32'd190799: dataIn1 = 32'd10474
; 
32'd190800: dataIn1 = 32'd10475
; 
32'd190801: dataIn1 = 32'd10476
; 
32'd190802: dataIn1 = 32'd216
; 
32'd190803: dataIn1 = 32'd830
; 
32'd190804: dataIn1 = 32'd1547
; 
32'd190805: dataIn1 = 32'd1549
; 
32'd190806: dataIn1 = 32'd10475
; 
32'd190807: dataIn1 = 32'd10476
; 
32'd190808: dataIn1 = 32'd10477
; 
32'd190809: dataIn1 = 32'd216
; 
32'd190810: dataIn1 = 32'd817
; 
32'd190811: dataIn1 = 32'd1534
; 
32'd190812: dataIn1 = 32'd1549
; 
32'd190813: dataIn1 = 32'd10476
; 
32'd190814: dataIn1 = 32'd10477
; 
32'd190815: dataIn1 = 32'd10478
; 
32'd190816: dataIn1 = 32'd817
; 
32'd190817: dataIn1 = 32'd818
; 
32'd190818: dataIn1 = 32'd1532
; 
32'd190819: dataIn1 = 32'd1534
; 
32'd190820: dataIn1 = 32'd10477
; 
32'd190821: dataIn1 = 32'd10478
; 
32'd190822: dataIn1 = 32'd10479
; 
32'd190823: dataIn1 = 32'd815
; 
32'd190824: dataIn1 = 32'd818
; 
32'd190825: dataIn1 = 32'd1532
; 
32'd190826: dataIn1 = 32'd1533
; 
32'd190827: dataIn1 = 32'd10478
; 
32'd190828: dataIn1 = 32'd10479
; 
32'd190829: dataIn1 = 32'd10480
; 
32'd190830: dataIn1 = 32'd418
; 
32'd190831: dataIn1 = 32'd815
; 
32'd190832: dataIn1 = 32'd1528
; 
32'd190833: dataIn1 = 32'd1533
; 
32'd190834: dataIn1 = 32'd10479
; 
32'd190835: dataIn1 = 32'd10480
; 
32'd190836: dataIn1 = 32'd10481
; 
32'd190837: dataIn1 = 32'd418
; 
32'd190838: dataIn1 = 32'd814
; 
32'd190839: dataIn1 = 32'd1528
; 
32'd190840: dataIn1 = 32'd1530
; 
32'd190841: dataIn1 = 32'd10480
; 
32'd190842: dataIn1 = 32'd10481
; 
32'd190843: dataIn1 = 32'd10482
; 
32'd190844: dataIn1 = 32'd814
; 
32'd190845: dataIn1 = 32'd816
; 
32'd190846: dataIn1 = 32'd1529
; 
32'd190847: dataIn1 = 32'd1530
; 
32'd190848: dataIn1 = 32'd10481
; 
32'd190849: dataIn1 = 32'd10482
; 
32'd190850: dataIn1 = 32'd10483
; 
32'd190851: dataIn1 = 32'd813
; 
32'd190852: dataIn1 = 32'd816
; 
32'd190853: dataIn1 = 32'd1529
; 
32'd190854: dataIn1 = 32'd1531
; 
32'd190855: dataIn1 = 32'd10482
; 
32'd190856: dataIn1 = 32'd10483
; 
32'd190857: dataIn1 = 32'd10484
; 
32'd190858: dataIn1 = 32'd214
; 
32'd190859: dataIn1 = 32'd813
; 
32'd190860: dataIn1 = 32'd1527
; 
32'd190861: dataIn1 = 32'd1531
; 
32'd190862: dataIn1 = 32'd10483
; 
32'd190863: dataIn1 = 32'd10484
; 
32'd190864: dataIn1 = 32'd10485
; 
32'd190865: dataIn1 = 32'd214
; 
32'd190866: dataIn1 = 32'd809
; 
32'd190867: dataIn1 = 32'd1522
; 
32'd190868: dataIn1 = 32'd1527
; 
32'd190869: dataIn1 = 32'd10484
; 
32'd190870: dataIn1 = 32'd10485
; 
32'd190871: dataIn1 = 32'd10486
; 
32'd190872: dataIn1 = 32'd809
; 
32'd190873: dataIn1 = 32'd810
; 
32'd190874: dataIn1 = 32'd1520
; 
32'd190875: dataIn1 = 32'd1522
; 
32'd190876: dataIn1 = 32'd10485
; 
32'd190877: dataIn1 = 32'd10486
; 
32'd190878: dataIn1 = 32'd10487
; 
32'd190879: dataIn1 = 32'd807
; 
32'd190880: dataIn1 = 32'd810
; 
32'd190881: dataIn1 = 32'd1520
; 
32'd190882: dataIn1 = 32'd1521
; 
32'd190883: dataIn1 = 32'd10486
; 
32'd190884: dataIn1 = 32'd10487
; 
32'd190885: dataIn1 = 32'd10488
; 
32'd190886: dataIn1 = 32'd417
; 
32'd190887: dataIn1 = 32'd807
; 
32'd190888: dataIn1 = 32'd1519
; 
32'd190889: dataIn1 = 32'd1521
; 
32'd190890: dataIn1 = 32'd10487
; 
32'd190891: dataIn1 = 32'd10488
; 
32'd190892: dataIn1 = 32'd10489
; 
32'd190893: dataIn1 = 32'd417
; 
32'd190894: dataIn1 = 32'd808
; 
32'd190895: dataIn1 = 32'd1519
; 
32'd190896: dataIn1 = 32'd1524
; 
32'd190897: dataIn1 = 32'd10488
; 
32'd190898: dataIn1 = 32'd10489
; 
32'd190899: dataIn1 = 32'd10490
; 
32'd190900: dataIn1 = 32'd808
; 
32'd190901: dataIn1 = 32'd812
; 
32'd190902: dataIn1 = 32'd1523
; 
32'd190903: dataIn1 = 32'd1524
; 
32'd190904: dataIn1 = 32'd10489
; 
32'd190905: dataIn1 = 32'd10490
; 
32'd190906: dataIn1 = 32'd10491
; 
32'd190907: dataIn1 = 32'd811
; 
32'd190908: dataIn1 = 32'd812
; 
32'd190909: dataIn1 = 32'd1523
; 
32'd190910: dataIn1 = 32'd1525
; 
32'd190911: dataIn1 = 32'd10490
; 
32'd190912: dataIn1 = 32'd10491
; 
32'd190913: dataIn1 = 32'd10492
; 
32'd190914: dataIn1 = 32'd213
; 
32'd190915: dataIn1 = 32'd811
; 
32'd190916: dataIn1 = 32'd1525
; 
32'd190917: dataIn1 = 32'd1526
; 
32'd190918: dataIn1 = 32'd10491
; 
32'd190919: dataIn1 = 32'd10492
; 
32'd190920: dataIn1 = 32'd10493
; 
32'd190921: dataIn1 = 32'd213
; 
32'd190922: dataIn1 = 32'd797
; 
32'd190923: dataIn1 = 32'd1505
; 
32'd190924: dataIn1 = 32'd1526
; 
32'd190925: dataIn1 = 32'd10492
; 
32'd190926: dataIn1 = 32'd10493
; 
32'd190927: dataIn1 = 32'd10494
; 
32'd190928: dataIn1 = 32'd796
; 
32'd190929: dataIn1 = 32'd797
; 
32'd190930: dataIn1 = 32'd1503
; 
32'd190931: dataIn1 = 32'd1505
; 
32'd190932: dataIn1 = 32'd10493
; 
32'd190933: dataIn1 = 32'd10494
; 
32'd190934: dataIn1 = 32'd10495
; 
32'd190935: dataIn1 = 32'd793
; 
32'd190936: dataIn1 = 32'd796
; 
32'd190937: dataIn1 = 32'd1503
; 
32'd190938: dataIn1 = 32'd1504
; 
32'd190939: dataIn1 = 32'd10494
; 
32'd190940: dataIn1 = 32'd10495
; 
32'd190941: dataIn1 = 32'd10496
; 
32'd190942: dataIn1 = 32'd412
; 
32'd190943: dataIn1 = 32'd793
; 
32'd190944: dataIn1 = 32'd1499
; 
32'd190945: dataIn1 = 32'd1504
; 
32'd190946: dataIn1 = 32'd10495
; 
32'd190947: dataIn1 = 32'd10496
; 
32'd190948: dataIn1 = 32'd10497
; 
32'd190949: dataIn1 = 32'd412
; 
32'd190950: dataIn1 = 32'd792
; 
32'd190951: dataIn1 = 32'd1499
; 
32'd190952: dataIn1 = 32'd1502
; 
32'd190953: dataIn1 = 32'd10496
; 
32'd190954: dataIn1 = 32'd10497
; 
32'd190955: dataIn1 = 32'd10498
; 
32'd190956: dataIn1 = 32'd792
; 
32'd190957: dataIn1 = 32'd795
; 
32'd190958: dataIn1 = 32'd1500
; 
32'd190959: dataIn1 = 32'd1502
; 
32'd190960: dataIn1 = 32'd10497
; 
32'd190961: dataIn1 = 32'd10498
; 
32'd190962: dataIn1 = 32'd10499
; 
32'd190963: dataIn1 = 32'd794
; 
32'd190964: dataIn1 = 32'd795
; 
32'd190965: dataIn1 = 32'd1500
; 
32'd190966: dataIn1 = 32'd1501
; 
32'd190967: dataIn1 = 32'd10498
; 
32'd190968: dataIn1 = 32'd10499
; 
32'd190969: dataIn1 = 32'd10500
; 
32'd190970: dataIn1 = 32'd211
; 
32'd190971: dataIn1 = 32'd794
; 
32'd190972: dataIn1 = 32'd1501
; 
32'd190973: dataIn1 = 32'd1515
; 
32'd190974: dataIn1 = 32'd10499
; 
32'd190975: dataIn1 = 32'd10500
; 
32'd190976: dataIn1 = 32'd10501
; 
32'd190977: dataIn1 = 32'd211
; 
32'd190978: dataIn1 = 32'd802
; 
32'd190979: dataIn1 = 32'd1508
; 
32'd190980: dataIn1 = 32'd1515
; 
32'd190981: dataIn1 = 32'd10500
; 
32'd190982: dataIn1 = 32'd10501
; 
32'd190983: dataIn1 = 32'd10502
; 
32'd190984: dataIn1 = 32'd801
; 
32'd190985: dataIn1 = 32'd802
; 
32'd190986: dataIn1 = 32'd1507
; 
32'd190987: dataIn1 = 32'd1508
; 
32'd190988: dataIn1 = 32'd10501
; 
32'd190989: dataIn1 = 32'd10502
; 
32'd190990: dataIn1 = 32'd10503
; 
32'd190991: dataIn1 = 32'd798
; 
32'd190992: dataIn1 = 32'd801
; 
32'd190993: dataIn1 = 32'd1507
; 
32'd190994: dataIn1 = 32'd1509
; 
32'd190995: dataIn1 = 32'd10502
; 
32'd190996: dataIn1 = 32'd10503
; 
32'd190997: dataIn1 = 32'd10504
; 
32'd190998: dataIn1 = 32'd415
; 
32'd190999: dataIn1 = 32'd798
; 
32'd191000: dataIn1 = 32'd1506
; 
32'd191001: dataIn1 = 32'd1509
; 
32'd191002: dataIn1 = 32'd10503
; 
32'd191003: dataIn1 = 32'd10504
; 
32'd191004: dataIn1 = 32'd10505
; 
32'd191005: dataIn1 = 32'd415
; 
32'd191006: dataIn1 = 32'd799
; 
32'd191007: dataIn1 = 32'd1506
; 
32'd191008: dataIn1 = 32'd1512
; 
32'd191009: dataIn1 = 32'd10504
; 
32'd191010: dataIn1 = 32'd10505
; 
32'd191011: dataIn1 = 32'd10506
; 
32'd191012: dataIn1 = 32'd799
; 
32'd191013: dataIn1 = 32'd803
; 
32'd191014: dataIn1 = 32'd1510
; 
32'd191015: dataIn1 = 32'd1512
; 
32'd191016: dataIn1 = 32'd10505
; 
32'd191017: dataIn1 = 32'd10506
; 
32'd191018: dataIn1 = 32'd10507
; 
32'd191019: dataIn1 = 32'd803
; 
32'd191020: dataIn1 = 32'd804
; 
32'd191021: dataIn1 = 32'd1510
; 
32'd191022: dataIn1 = 32'd1511
; 
32'd191023: dataIn1 = 32'd10506
; 
32'd191024: dataIn1 = 32'd10507
; 
32'd191025: dataIn1 = 32'd10508
; 
32'd191026: dataIn1 = 32'd210
; 
32'd191027: dataIn1 = 32'd804
; 
32'd191028: dataIn1 = 32'd1511
; 
32'd191029: dataIn1 = 32'd1513
; 
32'd191030: dataIn1 = 32'd10507
; 
32'd191031: dataIn1 = 32'd10508
; 
32'd191032: dataIn1 = 32'd10509
; 
32'd191033: dataIn1 = 32'd210
; 
32'd191034: dataIn1 = 32'd790
; 
32'd191035: dataIn1 = 32'd1498
; 
32'd191036: dataIn1 = 32'd1513
; 
32'd191037: dataIn1 = 32'd10508
; 
32'd191038: dataIn1 = 32'd10509
; 
32'd191039: dataIn1 = 32'd10510
; 
32'd191040: dataIn1 = 32'd790
; 
32'd191041: dataIn1 = 32'd791
; 
32'd191042: dataIn1 = 32'd1496
; 
32'd191043: dataIn1 = 32'd1498
; 
32'd191044: dataIn1 = 32'd10509
; 
32'd191045: dataIn1 = 32'd10510
; 
32'd191046: dataIn1 = 32'd10511
; 
32'd191047: dataIn1 = 32'd788
; 
32'd191048: dataIn1 = 32'd791
; 
32'd191049: dataIn1 = 32'd1496
; 
32'd191050: dataIn1 = 32'd1497
; 
32'd191051: dataIn1 = 32'd10510
; 
32'd191052: dataIn1 = 32'd10511
; 
32'd191053: dataIn1 = 32'd10512
; 
32'd191054: dataIn1 = 32'd410
; 
32'd191055: dataIn1 = 32'd788
; 
32'd191056: dataIn1 = 32'd1492
; 
32'd191057: dataIn1 = 32'd1497
; 
32'd191058: dataIn1 = 32'd10511
; 
32'd191059: dataIn1 = 32'd10512
; 
32'd191060: dataIn1 = 32'd10513
; 
32'd191061: dataIn1 = 32'd410
; 
32'd191062: dataIn1 = 32'd787
; 
32'd191063: dataIn1 = 32'd1492
; 
32'd191064: dataIn1 = 32'd1494
; 
32'd191065: dataIn1 = 32'd10512
; 
32'd191066: dataIn1 = 32'd10513
; 
32'd191067: dataIn1 = 32'd10514
; 
32'd191068: dataIn1 = 32'd787
; 
32'd191069: dataIn1 = 32'd789
; 
32'd191070: dataIn1 = 32'd1493
; 
32'd191071: dataIn1 = 32'd1494
; 
32'd191072: dataIn1 = 32'd10513
; 
32'd191073: dataIn1 = 32'd10514
; 
32'd191074: dataIn1 = 32'd10515
; 
32'd191075: dataIn1 = 32'd785
; 
32'd191076: dataIn1 = 32'd789
; 
32'd191077: dataIn1 = 32'd1493
; 
32'd191078: dataIn1 = 32'd1495
; 
32'd191079: dataIn1 = 32'd10514
; 
32'd191080: dataIn1 = 32'd10515
; 
32'd191081: dataIn1 = 32'd10516
; 
32'd191082: dataIn1 = 32'd208
; 
32'd191083: dataIn1 = 32'd785
; 
32'd191084: dataIn1 = 32'd1491
; 
32'd191085: dataIn1 = 32'd1495
; 
32'd191086: dataIn1 = 32'd10515
; 
32'd191087: dataIn1 = 32'd10516
; 
32'd191088: dataIn1 = 32'd10517
; 
32'd191089: dataIn1 = 32'd208
; 
32'd191090: dataIn1 = 32'd778
; 
32'd191091: dataIn1 = 32'd1484
; 
32'd191092: dataIn1 = 32'd1491
; 
32'd191093: dataIn1 = 32'd10516
; 
32'd191094: dataIn1 = 32'd10517
; 
32'd191095: dataIn1 = 32'd10518
; 
32'd191096: dataIn1 = 32'd778
; 
32'd191097: dataIn1 = 32'd779
; 
32'd191098: dataIn1 = 32'd1482
; 
32'd191099: dataIn1 = 32'd1484
; 
32'd191100: dataIn1 = 32'd10517
; 
32'd191101: dataIn1 = 32'd10518
; 
32'd191102: dataIn1 = 32'd10519
; 
32'd191103: dataIn1 = 32'd776
; 
32'd191104: dataIn1 = 32'd779
; 
32'd191105: dataIn1 = 32'd1482
; 
32'd191106: dataIn1 = 32'd1483
; 
32'd191107: dataIn1 = 32'd10518
; 
32'd191108: dataIn1 = 32'd10519
; 
32'd191109: dataIn1 = 32'd10520
; 
32'd191110: dataIn1 = 32'd406
; 
32'd191111: dataIn1 = 32'd776
; 
32'd191112: dataIn1 = 32'd1481
; 
32'd191113: dataIn1 = 32'd1483
; 
32'd191114: dataIn1 = 32'd10519
; 
32'd191115: dataIn1 = 32'd10520
; 
32'd191116: dataIn1 = 32'd10521
; 
32'd191117: dataIn1 = 32'd406
; 
32'd191118: dataIn1 = 32'd777
; 
32'd191119: dataIn1 = 32'd1481
; 
32'd191120: dataIn1 = 32'd1486
; 
32'd191121: dataIn1 = 32'd10520
; 
32'd191122: dataIn1 = 32'd10521
; 
32'd191123: dataIn1 = 32'd10522
; 
32'd191124: dataIn1 = 32'd777
; 
32'd191125: dataIn1 = 32'd781
; 
32'd191126: dataIn1 = 32'd1485
; 
32'd191127: dataIn1 = 32'd1486
; 
32'd191128: dataIn1 = 32'd10521
; 
32'd191129: dataIn1 = 32'd10522
; 
32'd191130: dataIn1 = 32'd10523
; 
32'd191131: dataIn1 = 32'd780
; 
32'd191132: dataIn1 = 32'd781
; 
32'd191133: dataIn1 = 32'd1485
; 
32'd191134: dataIn1 = 32'd1487
; 
32'd191135: dataIn1 = 32'd10522
; 
32'd191136: dataIn1 = 32'd10523
; 
32'd191137: dataIn1 = 32'd10524
; 
32'd191138: dataIn1 = 32'd207
; 
32'd191139: dataIn1 = 32'd780
; 
32'd191140: dataIn1 = 32'd1487
; 
32'd191141: dataIn1 = 32'd1490
; 
32'd191142: dataIn1 = 32'd10523
; 
32'd191143: dataIn1 = 32'd10524
; 
32'd191144: dataIn1 = 32'd10525
; 
32'd191145: dataIn1 = 32'd207
; 
32'd191146: dataIn1 = 32'd768
; 
32'd191147: dataIn1 = 32'd1463
; 
32'd191148: dataIn1 = 32'd1490
; 
32'd191149: dataIn1 = 32'd10524
; 
32'd191150: dataIn1 = 32'd10525
; 
32'd191151: dataIn1 = 32'd10526
; 
32'd191152: dataIn1 = 32'd766
; 
32'd191153: dataIn1 = 32'd768
; 
32'd191154: dataIn1 = 32'd1461
; 
32'd191155: dataIn1 = 32'd1463
; 
32'd191156: dataIn1 = 32'd10525
; 
32'd191157: dataIn1 = 32'd10526
; 
32'd191158: dataIn1 = 32'd10684
; 
32'd191159: dataIn1 = 32'd766
; 
32'd191160: dataIn1 = 32'd1460
; 
32'd191161: dataIn1 = 32'd10527
; 
32'd191162: dataIn1 = 32'd10528
; 
32'd191163: dataIn1 = 32'd10682
; 
32'd191164: dataIn1 = 32'd10684
; 
32'd191165: dataIn1 = 32'd10685
; 
32'd191166: dataIn1 = 32'd766
; 
32'd191167: dataIn1 = 32'd1460
; 
32'd191168: dataIn1 = 32'd10527
; 
32'd191169: dataIn1 = 32'd10528
; 
32'd191170: dataIn1 = 32'd10529
; 
32'd191171: dataIn1 = 32'd766
; 
32'd191172: dataIn1 = 32'd1459
; 
32'd191173: dataIn1 = 32'd1460
; 
32'd191174: dataIn1 = 32'd10528
; 
32'd191175: dataIn1 = 32'd10529
; 
32'd191176: dataIn1 = 32'd10530
; 
32'd191177: dataIn1 = 32'd402
; 
32'd191178: dataIn1 = 32'd1451
; 
32'd191179: dataIn1 = 32'd1459
; 
32'd191180: dataIn1 = 32'd1460
; 
32'd191181: dataIn1 = 32'd10529
; 
32'd191182: dataIn1 = 32'd10530
; 
32'd191183: dataIn1 = 32'd10531
; 
32'd191184: dataIn1 = 32'd402
; 
32'd191185: dataIn1 = 32'd1451
; 
32'd191186: dataIn1 = 32'd10530
; 
32'd191187: dataIn1 = 32'd10531
; 
32'd191188: dataIn1 = 32'd10532
; 
32'd191189: dataIn1 = 32'd402
; 
32'd191190: dataIn1 = 32'd1451
; 
32'd191191: dataIn1 = 32'd1453
; 
32'd191192: dataIn1 = 32'd1458
; 
32'd191193: dataIn1 = 32'd10531
; 
32'd191194: dataIn1 = 32'd10532
; 
32'd191195: dataIn1 = 32'd10533
; 
32'd191196: dataIn1 = 32'd1453
; 
32'd191197: dataIn1 = 32'd1458
; 
32'd191198: dataIn1 = 32'd10532
; 
32'd191199: dataIn1 = 32'd10533
; 
32'd191200: dataIn1 = 32'd10534
; 
32'd191201: dataIn1 = 32'd1453
; 
32'd191202: dataIn1 = 32'd1455
; 
32'd191203: dataIn1 = 32'd1458
; 
32'd191204: dataIn1 = 32'd10533
; 
32'd191205: dataIn1 = 32'd10534
; 
32'd191206: dataIn1 = 32'd10535
; 
32'd191207: dataIn1 = 32'd10678
; 
32'd191208: dataIn1 = 32'd1455
; 
32'd191209: dataIn1 = 32'd10534
; 
32'd191210: dataIn1 = 32'd10535
; 
32'd191211: dataIn1 = 32'd10536
; 
32'd191212: dataIn1 = 32'd10677
; 
32'd191213: dataIn1 = 32'd10678
; 
32'd191214: dataIn1 = 32'd1454
; 
32'd191215: dataIn1 = 32'd1455
; 
32'd191216: dataIn1 = 32'd10535
; 
32'd191217: dataIn1 = 32'd10536
; 
32'd191218: dataIn1 = 32'd10537
; 
32'd191219: dataIn1 = 32'd10676
; 
32'd191220: dataIn1 = 32'd10677
; 
32'd191221: dataIn1 = 32'd1454
; 
32'd191222: dataIn1 = 32'd10536
; 
32'd191223: dataIn1 = 32'd10537
; 
32'd191224: dataIn1 = 32'd10676
; 
32'd191225: dataIn1 = 32'd10686
; 
32'd191226: dataIn1 = 32'd1444
; 
32'd191227: dataIn1 = 32'd1446
; 
32'd191228: dataIn1 = 32'd10538
; 
32'd191229: dataIn1 = 32'd10539
; 
32'd191230: dataIn1 = 32'd10675
; 
32'd191231: dataIn1 = 32'd10706
; 
32'd191232: dataIn1 = 32'd757
; 
32'd191233: dataIn1 = 32'd1444
; 
32'd191234: dataIn1 = 32'd10538
; 
32'd191235: dataIn1 = 32'd10539
; 
32'd191236: dataIn1 = 32'd10540
; 
32'd191237: dataIn1 = 32'd10675
; 
32'd191238: dataIn1 = 32'd757
; 
32'd191239: dataIn1 = 32'd1442
; 
32'd191240: dataIn1 = 32'd1444
; 
32'd191241: dataIn1 = 32'd10539
; 
32'd191242: dataIn1 = 32'd10540
; 
32'd191243: dataIn1 = 32'd10541
; 
32'd191244: dataIn1 = 32'd757
; 
32'd191245: dataIn1 = 32'd1442
; 
32'd191246: dataIn1 = 32'd10540
; 
32'd191247: dataIn1 = 32'd10541
; 
32'd191248: dataIn1 = 32'd10542
; 
32'd191249: dataIn1 = 32'd757
; 
32'd191250: dataIn1 = 32'd1434
; 
32'd191251: dataIn1 = 32'd1442
; 
32'd191252: dataIn1 = 32'd1445
; 
32'd191253: dataIn1 = 32'd10541
; 
32'd191254: dataIn1 = 32'd10542
; 
32'd191255: dataIn1 = 32'd10543
; 
32'd191256: dataIn1 = 32'd1434
; 
32'd191257: dataIn1 = 32'd1445
; 
32'd191258: dataIn1 = 32'd10542
; 
32'd191259: dataIn1 = 32'd10543
; 
32'd191260: dataIn1 = 32'd10544
; 
32'd191261: dataIn1 = 32'd394
; 
32'd191262: dataIn1 = 32'd1434
; 
32'd191263: dataIn1 = 32'd1435
; 
32'd191264: dataIn1 = 32'd1445
; 
32'd191265: dataIn1 = 32'd10543
; 
32'd191266: dataIn1 = 32'd10544
; 
32'd191267: dataIn1 = 32'd10545
; 
32'd191268: dataIn1 = 32'd394
; 
32'd191269: dataIn1 = 32'd1435
; 
32'd191270: dataIn1 = 32'd10544
; 
32'd191271: dataIn1 = 32'd10545
; 
32'd191272: dataIn1 = 32'd10546
; 
32'd191273: dataIn1 = 32'd394
; 
32'd191274: dataIn1 = 32'd1435
; 
32'd191275: dataIn1 = 32'd1436
; 
32'd191276: dataIn1 = 32'd1439
; 
32'd191277: dataIn1 = 32'd10545
; 
32'd191278: dataIn1 = 32'd10546
; 
32'd191279: dataIn1 = 32'd10547
; 
32'd191280: dataIn1 = 32'd1436
; 
32'd191281: dataIn1 = 32'd1439
; 
32'd191282: dataIn1 = 32'd10546
; 
32'd191283: dataIn1 = 32'd10547
; 
32'd191284: dataIn1 = 32'd10548
; 
32'd191285: dataIn1 = 32'd755
; 
32'd191286: dataIn1 = 32'd1436
; 
32'd191287: dataIn1 = 32'd1437
; 
32'd191288: dataIn1 = 32'd1439
; 
32'd191289: dataIn1 = 32'd10547
; 
32'd191290: dataIn1 = 32'd10548
; 
32'd191291: dataIn1 = 32'd10549
; 
32'd191292: dataIn1 = 32'd755
; 
32'd191293: dataIn1 = 32'd1437
; 
32'd191294: dataIn1 = 32'd10548
; 
32'd191295: dataIn1 = 32'd10549
; 
32'd191296: dataIn1 = 32'd10550
; 
32'd191297: dataIn1 = 32'd755
; 
32'd191298: dataIn1 = 32'd1437
; 
32'd191299: dataIn1 = 32'd1440
; 
32'd191300: dataIn1 = 32'd10549
; 
32'd191301: dataIn1 = 32'd10550
; 
32'd191302: dataIn1 = 32'd10551
; 
32'd191303: dataIn1 = 32'd204
; 
32'd191304: dataIn1 = 32'd1437
; 
32'd191305: dataIn1 = 32'd1440
; 
32'd191306: dataIn1 = 32'd1441
; 
32'd191307: dataIn1 = 32'd10550
; 
32'd191308: dataIn1 = 32'd10551
; 
32'd191309: dataIn1 = 32'd10552
; 
32'd191310: dataIn1 = 32'd204
; 
32'd191311: dataIn1 = 32'd1441
; 
32'd191312: dataIn1 = 32'd10551
; 
32'd191313: dataIn1 = 32'd10552
; 
32'd191314: dataIn1 = 32'd10553
; 
32'd191315: dataIn1 = 32'd204
; 
32'd191316: dataIn1 = 32'd1430
; 
32'd191317: dataIn1 = 32'd1431
; 
32'd191318: dataIn1 = 32'd1441
; 
32'd191319: dataIn1 = 32'd10552
; 
32'd191320: dataIn1 = 32'd10553
; 
32'd191321: dataIn1 = 32'd10554
; 
32'd191322: dataIn1 = 32'd1430
; 
32'd191323: dataIn1 = 32'd1431
; 
32'd191324: dataIn1 = 32'd10553
; 
32'd191325: dataIn1 = 32'd10554
; 
32'd191326: dataIn1 = 32'd10555
; 
32'd191327: dataIn1 = 32'd746
; 
32'd191328: dataIn1 = 32'd1427
; 
32'd191329: dataIn1 = 32'd1430
; 
32'd191330: dataIn1 = 32'd1431
; 
32'd191331: dataIn1 = 32'd10554
; 
32'd191332: dataIn1 = 32'd10555
; 
32'd191333: dataIn1 = 32'd10556
; 
32'd191334: dataIn1 = 32'd746
; 
32'd191335: dataIn1 = 32'd1427
; 
32'd191336: dataIn1 = 32'd10555
; 
32'd191337: dataIn1 = 32'd10556
; 
32'd191338: dataIn1 = 32'd10557
; 
32'd191339: dataIn1 = 32'd746
; 
32'd191340: dataIn1 = 32'd1427
; 
32'd191341: dataIn1 = 32'd1428
; 
32'd191342: dataIn1 = 32'd10556
; 
32'd191343: dataIn1 = 32'd10557
; 
32'd191344: dataIn1 = 32'd10558
; 
32'd191345: dataIn1 = 32'd746
; 
32'd191346: dataIn1 = 32'd749
; 
32'd191347: dataIn1 = 32'd1428
; 
32'd191348: dataIn1 = 32'd1429
; 
32'd191349: dataIn1 = 32'd10557
; 
32'd191350: dataIn1 = 32'd10558
; 
32'd191351: dataIn1 = 32'd10559
; 
32'd191352: dataIn1 = 32'd389
; 
32'd191353: dataIn1 = 32'd746
; 
32'd191354: dataIn1 = 32'd1429
; 
32'd191355: dataIn1 = 32'd10558
; 
32'd191356: dataIn1 = 32'd10559
; 
32'd191357: dataIn1 = 32'd10560
; 
32'd191358: dataIn1 = 32'd389
; 
32'd191359: dataIn1 = 32'd746
; 
32'd191360: dataIn1 = 32'd1424
; 
32'd191361: dataIn1 = 32'd10559
; 
32'd191362: dataIn1 = 32'd10560
; 
32'd191363: dataIn1 = 32'd10561
; 
32'd191364: dataIn1 = 32'd389
; 
32'd191365: dataIn1 = 32'd1424
; 
32'd191366: dataIn1 = 32'd10560
; 
32'd191367: dataIn1 = 32'd10561
; 
32'd191368: dataIn1 = 32'd10707
; 
32'd191369: dataIn1 = 32'd10708
; 
32'd191370: dataIn1 = 32'd957
; 
32'd191371: dataIn1 = 32'd1719
; 
32'd191372: dataIn1 = 32'd10562
; 
32'd191373: dataIn1 = 32'd10762
; 
32'd191374: dataIn1 = 32'd728
; 
32'd191375: dataIn1 = 32'd1395
; 
32'd191376: dataIn1 = 32'd10563
; 
32'd191377: dataIn1 = 32'd11198
; 
32'd191378: dataIn1 = 32'd270
; 
32'd191379: dataIn1 = 32'd1271
; 
32'd191380: dataIn1 = 32'd1488
; 
32'd191381: dataIn1 = 32'd10564
; 
32'd191382: dataIn1 = 32'd11662
; 
32'd191383: dataIn1 = 32'd11663
; 
32'd191384: dataIn1 = 32'd1169
; 
32'd191385: dataIn1 = 32'd1170
; 
32'd191386: dataIn1 = 32'd10565
; 
32'd191387: dataIn1 = 32'd10566
; 
32'd191388: dataIn1 = 32'd11673
; 
32'd191389: dataIn1 = 32'd1158
; 
32'd191390: dataIn1 = 32'd1169
; 
32'd191391: dataIn1 = 32'd10565
; 
32'd191392: dataIn1 = 32'd10566
; 
32'd191393: dataIn1 = 32'd10567
; 
32'd191394: dataIn1 = 32'd1157
; 
32'd191395: dataIn1 = 32'd1158
; 
32'd191396: dataIn1 = 32'd10566
; 
32'd191397: dataIn1 = 32'd10567
; 
32'd191398: dataIn1 = 32'd10568
; 
32'd191399: dataIn1 = 32'd1157
; 
32'd191400: dataIn1 = 32'd10567
; 
32'd191401: dataIn1 = 32'd10568
; 
32'd191402: dataIn1 = 32'd10569
; 
32'd191403: dataIn1 = 32'd1153
; 
32'd191404: dataIn1 = 32'd1157
; 
32'd191405: dataIn1 = 32'd10568
; 
32'd191406: dataIn1 = 32'd10569
; 
32'd191407: dataIn1 = 32'd10570
; 
32'd191408: dataIn1 = 32'd1152
; 
32'd191409: dataIn1 = 32'd1153
; 
32'd191410: dataIn1 = 32'd10569
; 
32'd191411: dataIn1 = 32'd10570
; 
32'd191412: dataIn1 = 32'd10571
; 
32'd191413: dataIn1 = 32'd1152
; 
32'd191414: dataIn1 = 32'd1155
; 
32'd191415: dataIn1 = 32'd10570
; 
32'd191416: dataIn1 = 32'd10571
; 
32'd191417: dataIn1 = 32'd10572
; 
32'd191418: dataIn1 = 32'd1155
; 
32'd191419: dataIn1 = 32'd1159
; 
32'd191420: dataIn1 = 32'd10571
; 
32'd191421: dataIn1 = 32'd10572
; 
32'd191422: dataIn1 = 32'd10573
; 
32'd191423: dataIn1 = 32'd1159
; 
32'd191424: dataIn1 = 32'd1163
; 
32'd191425: dataIn1 = 32'd10572
; 
32'd191426: dataIn1 = 32'd10573
; 
32'd191427: dataIn1 = 32'd10574
; 
32'd191428: dataIn1 = 32'd1163
; 
32'd191429: dataIn1 = 32'd1164
; 
32'd191430: dataIn1 = 32'd10573
; 
32'd191431: dataIn1 = 32'd10574
; 
32'd191432: dataIn1 = 32'd10575
; 
32'd191433: dataIn1 = 32'd1150
; 
32'd191434: dataIn1 = 32'd1164
; 
32'd191435: dataIn1 = 32'd10574
; 
32'd191436: dataIn1 = 32'd10575
; 
32'd191437: dataIn1 = 32'd10576
; 
32'd191438: dataIn1 = 32'd1147
; 
32'd191439: dataIn1 = 32'd1150
; 
32'd191440: dataIn1 = 32'd10575
; 
32'd191441: dataIn1 = 32'd10576
; 
32'd191442: dataIn1 = 32'd10577
; 
32'd191443: dataIn1 = 32'd1144
; 
32'd191444: dataIn1 = 32'd1147
; 
32'd191445: dataIn1 = 32'd10576
; 
32'd191446: dataIn1 = 32'd10577
; 
32'd191447: dataIn1 = 32'd10578
; 
32'd191448: dataIn1 = 32'd1143
; 
32'd191449: dataIn1 = 32'd1144
; 
32'd191450: dataIn1 = 32'd10577
; 
32'd191451: dataIn1 = 32'd10578
; 
32'd191452: dataIn1 = 32'd10579
; 
32'd191453: dataIn1 = 32'd1143
; 
32'd191454: dataIn1 = 32'd1145
; 
32'd191455: dataIn1 = 32'd10578
; 
32'd191456: dataIn1 = 32'd10579
; 
32'd191457: dataIn1 = 32'd10580
; 
32'd191458: dataIn1 = 32'd1145
; 
32'd191459: dataIn1 = 32'd1151
; 
32'd191460: dataIn1 = 32'd10579
; 
32'd191461: dataIn1 = 32'd10580
; 
32'd191462: dataIn1 = 32'd10581
; 
32'd191463: dataIn1 = 32'd1151
; 
32'd191464: dataIn1 = 32'd1188
; 
32'd191465: dataIn1 = 32'd1189
; 
32'd191466: dataIn1 = 32'd10580
; 
32'd191467: dataIn1 = 32'd10581
; 
32'd191468: dataIn1 = 32'd10582
; 
32'd191469: dataIn1 = 32'd1184
; 
32'd191470: dataIn1 = 32'd1188
; 
32'd191471: dataIn1 = 32'd10581
; 
32'd191472: dataIn1 = 32'd10582
; 
32'd191473: dataIn1 = 32'd10583
; 
32'd191474: dataIn1 = 32'd1178
; 
32'd191475: dataIn1 = 32'd1184
; 
32'd191476: dataIn1 = 32'd10582
; 
32'd191477: dataIn1 = 32'd10583
; 
32'd191478: dataIn1 = 32'd10584
; 
32'd191479: dataIn1 = 32'd1176
; 
32'd191480: dataIn1 = 32'd1178
; 
32'd191481: dataIn1 = 32'd10583
; 
32'd191482: dataIn1 = 32'd10584
; 
32'd191483: dataIn1 = 32'd10585
; 
32'd191484: dataIn1 = 32'd1176
; 
32'd191485: dataIn1 = 32'd1177
; 
32'd191486: dataIn1 = 32'd10584
; 
32'd191487: dataIn1 = 32'd10585
; 
32'd191488: dataIn1 = 32'd10586
; 
32'd191489: dataIn1 = 32'd1177
; 
32'd191490: dataIn1 = 32'd1181
; 
32'd191491: dataIn1 = 32'd10585
; 
32'd191492: dataIn1 = 32'd10586
; 
32'd191493: dataIn1 = 32'd10587
; 
32'd191494: dataIn1 = 32'd1181
; 
32'd191495: dataIn1 = 32'd1182
; 
32'd191496: dataIn1 = 32'd10586
; 
32'd191497: dataIn1 = 32'd10587
; 
32'd191498: dataIn1 = 32'd10588
; 
32'd191499: dataIn1 = 32'd1182
; 
32'd191500: dataIn1 = 32'd1194
; 
32'd191501: dataIn1 = 32'd10587
; 
32'd191502: dataIn1 = 32'd10588
; 
32'd191503: dataIn1 = 32'd10589
; 
32'd191504: dataIn1 = 32'd1193
; 
32'd191505: dataIn1 = 32'd1194
; 
32'd191506: dataIn1 = 32'd10588
; 
32'd191507: dataIn1 = 32'd10589
; 
32'd191508: dataIn1 = 32'd10590
; 
32'd191509: dataIn1 = 32'd1193
; 
32'd191510: dataIn1 = 32'd1195
; 
32'd191511: dataIn1 = 32'd10589
; 
32'd191512: dataIn1 = 32'd10590
; 
32'd191513: dataIn1 = 32'd10591
; 
32'd191514: dataIn1 = 32'd1195
; 
32'd191515: dataIn1 = 32'd1205
; 
32'd191516: dataIn1 = 32'd10590
; 
32'd191517: dataIn1 = 32'd10591
; 
32'd191518: dataIn1 = 32'd10592
; 
32'd191519: dataIn1 = 32'd1205
; 
32'd191520: dataIn1 = 32'd10591
; 
32'd191521: dataIn1 = 32'd10592
; 
32'd191522: dataIn1 = 32'd10593
; 
32'd191523: dataIn1 = 32'd1201
; 
32'd191524: dataIn1 = 32'd1205
; 
32'd191525: dataIn1 = 32'd10592
; 
32'd191526: dataIn1 = 32'd10593
; 
32'd191527: dataIn1 = 32'd10594
; 
32'd191528: dataIn1 = 32'd1201
; 
32'd191529: dataIn1 = 32'd10593
; 
32'd191530: dataIn1 = 32'd10594
; 
32'd191531: dataIn1 = 32'd10595
; 
32'd191532: dataIn1 = 32'd1200
; 
32'd191533: dataIn1 = 32'd1201
; 
32'd191534: dataIn1 = 32'd10594
; 
32'd191535: dataIn1 = 32'd10595
; 
32'd191536: dataIn1 = 32'd10596
; 
32'd191537: dataIn1 = 32'd1200
; 
32'd191538: dataIn1 = 32'd10595
; 
32'd191539: dataIn1 = 32'd10596
; 
32'd191540: dataIn1 = 32'd10597
; 
32'd191541: dataIn1 = 32'd1200
; 
32'd191542: dataIn1 = 32'd1202
; 
32'd191543: dataIn1 = 32'd10596
; 
32'd191544: dataIn1 = 32'd10597
; 
32'd191545: dataIn1 = 32'd10598
; 
32'd191546: dataIn1 = 32'd1202
; 
32'd191547: dataIn1 = 32'd10597
; 
32'd191548: dataIn1 = 32'd10598
; 
32'd191549: dataIn1 = 32'd10599
; 
32'd191550: dataIn1 = 32'd1202
; 
32'd191551: dataIn1 = 32'd1207
; 
32'd191552: dataIn1 = 32'd10598
; 
32'd191553: dataIn1 = 32'd10599
; 
32'd191554: dataIn1 = 32'd10600
; 
32'd191555: dataIn1 = 32'd1207
; 
32'd191556: dataIn1 = 32'd10599
; 
32'd191557: dataIn1 = 32'd10600
; 
32'd191558: dataIn1 = 32'd10601
; 
32'd191559: dataIn1 = 32'd1207
; 
32'd191560: dataIn1 = 32'd1235
; 
32'd191561: dataIn1 = 32'd10600
; 
32'd191562: dataIn1 = 32'd10601
; 
32'd191563: dataIn1 = 32'd10602
; 
32'd191564: dataIn1 = 32'd1235
; 
32'd191565: dataIn1 = 32'd10601
; 
32'd191566: dataIn1 = 32'd10602
; 
32'd191567: dataIn1 = 32'd10603
; 
32'd191568: dataIn1 = 32'd1234
; 
32'd191569: dataIn1 = 32'd1235
; 
32'd191570: dataIn1 = 32'd10602
; 
32'd191571: dataIn1 = 32'd10603
; 
32'd191572: dataIn1 = 32'd10604
; 
32'd191573: dataIn1 = 32'd1234
; 
32'd191574: dataIn1 = 32'd10603
; 
32'd191575: dataIn1 = 32'd10604
; 
32'd191576: dataIn1 = 32'd10605
; 
32'd191577: dataIn1 = 32'd1223
; 
32'd191578: dataIn1 = 32'd1234
; 
32'd191579: dataIn1 = 32'd10604
; 
32'd191580: dataIn1 = 32'd10605
; 
32'd191581: dataIn1 = 32'd10606
; 
32'd191582: dataIn1 = 32'd1223
; 
32'd191583: dataIn1 = 32'd10605
; 
32'd191584: dataIn1 = 32'd10606
; 
32'd191585: dataIn1 = 32'd10607
; 
32'd191586: dataIn1 = 32'd1222
; 
32'd191587: dataIn1 = 32'd1223
; 
32'd191588: dataIn1 = 32'd10606
; 
32'd191589: dataIn1 = 32'd10607
; 
32'd191590: dataIn1 = 32'd10608
; 
32'd191591: dataIn1 = 32'd1222
; 
32'd191592: dataIn1 = 32'd10607
; 
32'd191593: dataIn1 = 32'd10608
; 
32'd191594: dataIn1 = 32'd10609
; 
32'd191595: dataIn1 = 32'd1222
; 
32'd191596: dataIn1 = 32'd10608
; 
32'd191597: dataIn1 = 32'd10609
; 
32'd191598: dataIn1 = 32'd10610
; 
32'd191599: dataIn1 = 32'd1218
; 
32'd191600: dataIn1 = 32'd1222
; 
32'd191601: dataIn1 = 32'd10609
; 
32'd191602: dataIn1 = 32'd10610
; 
32'd191603: dataIn1 = 32'd10611
; 
32'd191604: dataIn1 = 32'd1218
; 
32'd191605: dataIn1 = 32'd10610
; 
32'd191606: dataIn1 = 32'd10611
; 
32'd191607: dataIn1 = 32'd10612
; 
32'd191608: dataIn1 = 32'd1217
; 
32'd191609: dataIn1 = 32'd1218
; 
32'd191610: dataIn1 = 32'd10611
; 
32'd191611: dataIn1 = 32'd10612
; 
32'd191612: dataIn1 = 32'd10613
; 
32'd191613: dataIn1 = 32'd1217
; 
32'd191614: dataIn1 = 32'd10612
; 
32'd191615: dataIn1 = 32'd10613
; 
32'd191616: dataIn1 = 32'd10614
; 
32'd191617: dataIn1 = 32'd1217
; 
32'd191618: dataIn1 = 32'd1220
; 
32'd191619: dataIn1 = 32'd10613
; 
32'd191620: dataIn1 = 32'd10614
; 
32'd191621: dataIn1 = 32'd10615
; 
32'd191622: dataIn1 = 32'd1220
; 
32'd191623: dataIn1 = 32'd10614
; 
32'd191624: dataIn1 = 32'd10615
; 
32'd191625: dataIn1 = 32'd10616
; 
32'd191626: dataIn1 = 32'd1220
; 
32'd191627: dataIn1 = 32'd1224
; 
32'd191628: dataIn1 = 32'd10615
; 
32'd191629: dataIn1 = 32'd10616
; 
32'd191630: dataIn1 = 32'd10617
; 
32'd191631: dataIn1 = 32'd1224
; 
32'd191632: dataIn1 = 32'd10616
; 
32'd191633: dataIn1 = 32'd10617
; 
32'd191634: dataIn1 = 32'd10618
; 
32'd191635: dataIn1 = 32'd1224
; 
32'd191636: dataIn1 = 32'd1228
; 
32'd191637: dataIn1 = 32'd10617
; 
32'd191638: dataIn1 = 32'd10618
; 
32'd191639: dataIn1 = 32'd10619
; 
32'd191640: dataIn1 = 32'd1228
; 
32'd191641: dataIn1 = 32'd10618
; 
32'd191642: dataIn1 = 32'd10619
; 
32'd191643: dataIn1 = 32'd10620
; 
32'd191644: dataIn1 = 32'd1228
; 
32'd191645: dataIn1 = 32'd1229
; 
32'd191646: dataIn1 = 32'd10619
; 
32'd191647: dataIn1 = 32'd10620
; 
32'd191648: dataIn1 = 32'd10621
; 
32'd191649: dataIn1 = 32'd1215
; 
32'd191650: dataIn1 = 32'd1229
; 
32'd191651: dataIn1 = 32'd10620
; 
32'd191652: dataIn1 = 32'd10621
; 
32'd191653: dataIn1 = 32'd10622
; 
32'd191654: dataIn1 = 32'd1215
; 
32'd191655: dataIn1 = 32'd10621
; 
32'd191656: dataIn1 = 32'd10622
; 
32'd191657: dataIn1 = 32'd10623
; 
32'd191658: dataIn1 = 32'd1212
; 
32'd191659: dataIn1 = 32'd1215
; 
32'd191660: dataIn1 = 32'd10622
; 
32'd191661: dataIn1 = 32'd10623
; 
32'd191662: dataIn1 = 32'd10624
; 
32'd191663: dataIn1 = 32'd1212
; 
32'd191664: dataIn1 = 32'd10623
; 
32'd191665: dataIn1 = 32'd10624
; 
32'd191666: dataIn1 = 32'd10625
; 
32'd191667: dataIn1 = 32'd1209
; 
32'd191668: dataIn1 = 32'd1212
; 
32'd191669: dataIn1 = 32'd10624
; 
32'd191670: dataIn1 = 32'd10625
; 
32'd191671: dataIn1 = 32'd10626
; 
32'd191672: dataIn1 = 32'd1209
; 
32'd191673: dataIn1 = 32'd10625
; 
32'd191674: dataIn1 = 32'd10626
; 
32'd191675: dataIn1 = 32'd10627
; 
32'd191676: dataIn1 = 32'd1208
; 
32'd191677: dataIn1 = 32'd1209
; 
32'd191678: dataIn1 = 32'd10626
; 
32'd191679: dataIn1 = 32'd10627
; 
32'd191680: dataIn1 = 32'd10628
; 
32'd191681: dataIn1 = 32'd1208
; 
32'd191682: dataIn1 = 32'd10627
; 
32'd191683: dataIn1 = 32'd10628
; 
32'd191684: dataIn1 = 32'd10629
; 
32'd191685: dataIn1 = 32'd1208
; 
32'd191686: dataIn1 = 32'd1210
; 
32'd191687: dataIn1 = 32'd10628
; 
32'd191688: dataIn1 = 32'd10629
; 
32'd191689: dataIn1 = 32'd10630
; 
32'd191690: dataIn1 = 32'd1210
; 
32'd191691: dataIn1 = 32'd10629
; 
32'd191692: dataIn1 = 32'd10630
; 
32'd191693: dataIn1 = 32'd10631
; 
32'd191694: dataIn1 = 32'd1210
; 
32'd191695: dataIn1 = 32'd1216
; 
32'd191696: dataIn1 = 32'd10630
; 
32'd191697: dataIn1 = 32'd10631
; 
32'd191698: dataIn1 = 32'd10632
; 
32'd191699: dataIn1 = 32'd1216
; 
32'd191700: dataIn1 = 32'd10631
; 
32'd191701: dataIn1 = 32'd10632
; 
32'd191702: dataIn1 = 32'd10633
; 
32'd191703: dataIn1 = 32'd1216
; 
32'd191704: dataIn1 = 32'd1255
; 
32'd191705: dataIn1 = 32'd10632
; 
32'd191706: dataIn1 = 32'd10633
; 
32'd191707: dataIn1 = 32'd10634
; 
32'd191708: dataIn1 = 32'd1255
; 
32'd191709: dataIn1 = 32'd10633
; 
32'd191710: dataIn1 = 32'd10634
; 
32'd191711: dataIn1 = 32'd10635
; 
32'd191712: dataIn1 = 32'd1254
; 
32'd191713: dataIn1 = 32'd1255
; 
32'd191714: dataIn1 = 32'd10634
; 
32'd191715: dataIn1 = 32'd10635
; 
32'd191716: dataIn1 = 32'd10636
; 
32'd191717: dataIn1 = 32'd1254
; 
32'd191718: dataIn1 = 32'd10635
; 
32'd191719: dataIn1 = 32'd10636
; 
32'd191720: dataIn1 = 32'd10637
; 
32'd191721: dataIn1 = 32'd1250
; 
32'd191722: dataIn1 = 32'd1254
; 
32'd191723: dataIn1 = 32'd10636
; 
32'd191724: dataIn1 = 32'd10637
; 
32'd191725: dataIn1 = 32'd10638
; 
32'd191726: dataIn1 = 32'd1250
; 
32'd191727: dataIn1 = 32'd10637
; 
32'd191728: dataIn1 = 32'd10638
; 
32'd191729: dataIn1 = 32'd10639
; 
32'd191730: dataIn1 = 32'd1242
; 
32'd191731: dataIn1 = 32'd1250
; 
32'd191732: dataIn1 = 32'd10638
; 
32'd191733: dataIn1 = 32'd10639
; 
32'd191734: dataIn1 = 32'd10640
; 
32'd191735: dataIn1 = 32'd1242
; 
32'd191736: dataIn1 = 32'd10639
; 
32'd191737: dataIn1 = 32'd10640
; 
32'd191738: dataIn1 = 32'd10641
; 
32'd191739: dataIn1 = 32'd1240
; 
32'd191740: dataIn1 = 32'd1242
; 
32'd191741: dataIn1 = 32'd10640
; 
32'd191742: dataIn1 = 32'd10641
; 
32'd191743: dataIn1 = 32'd10642
; 
32'd191744: dataIn1 = 32'd1240
; 
32'd191745: dataIn1 = 32'd10641
; 
32'd191746: dataIn1 = 32'd10642
; 
32'd191747: dataIn1 = 32'd10643
; 
32'd191748: dataIn1 = 32'd1240
; 
32'd191749: dataIn1 = 32'd1241
; 
32'd191750: dataIn1 = 32'd10642
; 
32'd191751: dataIn1 = 32'd10643
; 
32'd191752: dataIn1 = 32'd10644
; 
32'd191753: dataIn1 = 32'd1241
; 
32'd191754: dataIn1 = 32'd10643
; 
32'd191755: dataIn1 = 32'd10644
; 
32'd191756: dataIn1 = 32'd10645
; 
32'd191757: dataIn1 = 32'd1241
; 
32'd191758: dataIn1 = 32'd1245
; 
32'd191759: dataIn1 = 32'd10644
; 
32'd191760: dataIn1 = 32'd10645
; 
32'd191761: dataIn1 = 32'd10646
; 
32'd191762: dataIn1 = 32'd1245
; 
32'd191763: dataIn1 = 32'd10645
; 
32'd191764: dataIn1 = 32'd10646
; 
32'd191765: dataIn1 = 32'd10647
; 
32'd191766: dataIn1 = 32'd1245
; 
32'd191767: dataIn1 = 32'd1246
; 
32'd191768: dataIn1 = 32'd10646
; 
32'd191769: dataIn1 = 32'd10647
; 
32'd191770: dataIn1 = 32'd10648
; 
32'd191771: dataIn1 = 32'd1246
; 
32'd191772: dataIn1 = 32'd10647
; 
32'd191773: dataIn1 = 32'd10648
; 
32'd191774: dataIn1 = 32'd10649
; 
32'd191775: dataIn1 = 32'd1246
; 
32'd191776: dataIn1 = 32'd10648
; 
32'd191777: dataIn1 = 32'd10649
; 
32'd191778: dataIn1 = 32'd10650
; 
32'd191779: dataIn1 = 32'd1246
; 
32'd191780: dataIn1 = 32'd1258
; 
32'd191781: dataIn1 = 32'd10649
; 
32'd191782: dataIn1 = 32'd10650
; 
32'd191783: dataIn1 = 32'd10651
; 
32'd191784: dataIn1 = 32'd1258
; 
32'd191785: dataIn1 = 32'd10650
; 
32'd191786: dataIn1 = 32'd10651
; 
32'd191787: dataIn1 = 32'd10652
; 
32'd191788: dataIn1 = 32'd547
; 
32'd191789: dataIn1 = 32'd1258
; 
32'd191790: dataIn1 = 32'd1259
; 
32'd191791: dataIn1 = 32'd10651
; 
32'd191792: dataIn1 = 32'd10652
; 
32'd191793: dataIn1 = 32'd10653
; 
32'd191794: dataIn1 = 32'd1259
; 
32'd191795: dataIn1 = 32'd10652
; 
32'd191796: dataIn1 = 32'd10653
; 
32'd191797: dataIn1 = 32'd10654
; 
32'd191798: dataIn1 = 32'd267
; 
32'd191799: dataIn1 = 32'd1259
; 
32'd191800: dataIn1 = 32'd10653
; 
32'd191801: dataIn1 = 32'd10654
; 
32'd191802: dataIn1 = 32'd10655
; 
32'd191803: dataIn1 = 32'd267
; 
32'd191804: dataIn1 = 32'd10654
; 
32'd191805: dataIn1 = 32'd10655
; 
32'd191806: dataIn1 = 32'd10656
; 
32'd191807: dataIn1 = 32'd267
; 
32'd191808: dataIn1 = 32'd1266
; 
32'd191809: dataIn1 = 32'd10655
; 
32'd191810: dataIn1 = 32'd10656
; 
32'd191811: dataIn1 = 32'd10657
; 
32'd191812: dataIn1 = 32'd1266
; 
32'd191813: dataIn1 = 32'd10656
; 
32'd191814: dataIn1 = 32'd10657
; 
32'd191815: dataIn1 = 32'd10658
; 
32'd191816: dataIn1 = 32'd550
; 
32'd191817: dataIn1 = 32'd1263
; 
32'd191818: dataIn1 = 32'd1266
; 
32'd191819: dataIn1 = 32'd10657
; 
32'd191820: dataIn1 = 32'd10658
; 
32'd191821: dataIn1 = 32'd10659
; 
32'd191822: dataIn1 = 32'd1263
; 
32'd191823: dataIn1 = 32'd10658
; 
32'd191824: dataIn1 = 32'd10659
; 
32'd191825: dataIn1 = 32'd10660
; 
32'd191826: dataIn1 = 32'd1263
; 
32'd191827: dataIn1 = 32'd1264
; 
32'd191828: dataIn1 = 32'd10659
; 
32'd191829: dataIn1 = 32'd10660
; 
32'd191830: dataIn1 = 32'd10661
; 
32'd191831: dataIn1 = 32'd1264
; 
32'd191832: dataIn1 = 32'd10660
; 
32'd191833: dataIn1 = 32'd10661
; 
32'd191834: dataIn1 = 32'd10662
; 
32'd191835: dataIn1 = 32'd1264
; 
32'd191836: dataIn1 = 32'd1267
; 
32'd191837: dataIn1 = 32'd10661
; 
32'd191838: dataIn1 = 32'd10662
; 
32'd191839: dataIn1 = 32'd10663
; 
32'd191840: dataIn1 = 32'd1267
; 
32'd191841: dataIn1 = 32'd10662
; 
32'd191842: dataIn1 = 32'd10663
; 
32'd191843: dataIn1 = 32'd10664
; 
32'd191844: dataIn1 = 32'd1267
; 
32'd191845: dataIn1 = 32'd10663
; 
32'd191846: dataIn1 = 32'd10664
; 
32'd191847: dataIn1 = 32'd10665
; 
32'd191848: dataIn1 = 32'd1267
; 
32'd191849: dataIn1 = 32'd1467
; 
32'd191850: dataIn1 = 32'd10664
; 
32'd191851: dataIn1 = 32'd10665
; 
32'd191852: dataIn1 = 32'd10666
; 
32'd191853: dataIn1 = 32'd1467
; 
32'd191854: dataIn1 = 32'd10665
; 
32'd191855: dataIn1 = 32'd10666
; 
32'd191856: dataIn1 = 32'd10667
; 
32'd191857: dataIn1 = 32'd1467
; 
32'd191858: dataIn1 = 32'd1468
; 
32'd191859: dataIn1 = 32'd10666
; 
32'd191860: dataIn1 = 32'd10667
; 
32'd191861: dataIn1 = 32'd10668
; 
32'd191862: dataIn1 = 32'd1468
; 
32'd191863: dataIn1 = 32'd10667
; 
32'd191864: dataIn1 = 32'd10668
; 
32'd191865: dataIn1 = 32'd10669
; 
32'd191866: dataIn1 = 32'd1466
; 
32'd191867: dataIn1 = 32'd1468
; 
32'd191868: dataIn1 = 32'd10668
; 
32'd191869: dataIn1 = 32'd10669
; 
32'd191870: dataIn1 = 32'd10670
; 
32'd191871: dataIn1 = 32'd1466
; 
32'd191872: dataIn1 = 32'd10669
; 
32'd191873: dataIn1 = 32'd10670
; 
32'd191874: dataIn1 = 32'd10671
; 
32'd191875: dataIn1 = 32'd397
; 
32'd191876: dataIn1 = 32'd1466
; 
32'd191877: dataIn1 = 32'd1471
; 
32'd191878: dataIn1 = 32'd10670
; 
32'd191879: dataIn1 = 32'd10671
; 
32'd191880: dataIn1 = 32'd10672
; 
32'd191881: dataIn1 = 32'd1471
; 
32'd191882: dataIn1 = 32'd10671
; 
32'd191883: dataIn1 = 32'd10672
; 
32'd191884: dataIn1 = 32'd10673
; 
32'd191885: dataIn1 = 32'd1447
; 
32'd191886: dataIn1 = 32'd1471
; 
32'd191887: dataIn1 = 32'd3461
; 
32'd191888: dataIn1 = 32'd10672
; 
32'd191889: dataIn1 = 32'd10673
; 
32'd191890: dataIn1 = 32'd10674
; 
32'd191891: dataIn1 = 32'd1447
; 
32'd191892: dataIn1 = 32'd10673
; 
32'd191893: dataIn1 = 32'd10674
; 
32'd191894: dataIn1 = 32'd10675
; 
32'd191895: dataIn1 = 32'd757
; 
32'd191896: dataIn1 = 32'd1447
; 
32'd191897: dataIn1 = 32'd10538
; 
32'd191898: dataIn1 = 32'd10539
; 
32'd191899: dataIn1 = 32'd10674
; 
32'd191900: dataIn1 = 32'd10675
; 
32'd191901: dataIn1 = 32'd10536
; 
32'd191902: dataIn1 = 32'd10537
; 
32'd191903: dataIn1 = 32'd10676
; 
32'd191904: dataIn1 = 32'd10677
; 
32'd191905: dataIn1 = 32'd10686
; 
32'd191906: dataIn1 = 32'd10535
; 
32'd191907: dataIn1 = 32'd10536
; 
32'd191908: dataIn1 = 32'd10676
; 
32'd191909: dataIn1 = 32'd10677
; 
32'd191910: dataIn1 = 32'd10678
; 
32'd191911: dataIn1 = 32'd1458
; 
32'd191912: dataIn1 = 32'd10534
; 
32'd191913: dataIn1 = 32'd10535
; 
32'd191914: dataIn1 = 32'd10677
; 
32'd191915: dataIn1 = 32'd10678
; 
32'd191916: dataIn1 = 32'd10679
; 
32'd191917: dataIn1 = 32'd402
; 
32'd191918: dataIn1 = 32'd1458
; 
32'd191919: dataIn1 = 32'd10678
; 
32'd191920: dataIn1 = 32'd10679
; 
32'd191921: dataIn1 = 32'd10680
; 
32'd191922: dataIn1 = 32'd402
; 
32'd191923: dataIn1 = 32'd10679
; 
32'd191924: dataIn1 = 32'd10680
; 
32'd191925: dataIn1 = 32'd10681
; 
32'd191926: dataIn1 = 32'd402
; 
32'd191927: dataIn1 = 32'd1460
; 
32'd191928: dataIn1 = 32'd10680
; 
32'd191929: dataIn1 = 32'd10681
; 
32'd191930: dataIn1 = 32'd10682
; 
32'd191931: dataIn1 = 32'd1460
; 
32'd191932: dataIn1 = 32'd10527
; 
32'd191933: dataIn1 = 32'd10681
; 
32'd191934: dataIn1 = 32'd10682
; 
32'd191935: dataIn1 = 32'd516
; 
32'd191936: dataIn1 = 32'd10683
; 
32'd191937: dataIn1 = 32'd11674
; 
32'd191938: dataIn1 = 32'd766
; 
32'd191939: dataIn1 = 32'd1461
; 
32'd191940: dataIn1 = 32'd10526
; 
32'd191941: dataIn1 = 32'd10527
; 
32'd191942: dataIn1 = 32'd10684
; 
32'd191943: dataIn1 = 32'd10685
; 
32'd191944: dataIn1 = 32'd11672
; 
32'd191945: dataIn1 = 32'd10527
; 
32'd191946: dataIn1 = 32'd10684
; 
32'd191947: dataIn1 = 32'd10685
; 
32'd191948: dataIn1 = 32'd1454
; 
32'd191949: dataIn1 = 32'd1457
; 
32'd191950: dataIn1 = 32'd10537
; 
32'd191951: dataIn1 = 32'd10676
; 
32'd191952: dataIn1 = 32'd10686
; 
32'd191953: dataIn1 = 32'd10687
; 
32'd191954: dataIn1 = 32'd1457
; 
32'd191955: dataIn1 = 32'd10686
; 
32'd191956: dataIn1 = 32'd10687
; 
32'd191957: dataIn1 = 32'd10688
; 
32'd191958: dataIn1 = 32'd1457
; 
32'd191959: dataIn1 = 32'd1465
; 
32'd191960: dataIn1 = 32'd10687
; 
32'd191961: dataIn1 = 32'd10688
; 
32'd191962: dataIn1 = 32'd10689
; 
32'd191963: dataIn1 = 32'd1465
; 
32'd191964: dataIn1 = 32'd10688
; 
32'd191965: dataIn1 = 32'd10689
; 
32'd191966: dataIn1 = 32'd10690
; 
32'd191967: dataIn1 = 32'd1465
; 
32'd191968: dataIn1 = 32'd10689
; 
32'd191969: dataIn1 = 32'd10690
; 
32'd191970: dataIn1 = 32'd10691
; 
32'd191971: dataIn1 = 32'd1465
; 
32'd191972: dataIn1 = 32'd1475
; 
32'd191973: dataIn1 = 32'd10690
; 
32'd191974: dataIn1 = 32'd10691
; 
32'd191975: dataIn1 = 32'd10692
; 
32'd191976: dataIn1 = 32'd1475
; 
32'd191977: dataIn1 = 32'd10691
; 
32'd191978: dataIn1 = 32'd10692
; 
32'd191979: dataIn1 = 32'd10693
; 
32'd191980: dataIn1 = 32'd1475
; 
32'd191981: dataIn1 = 32'd1477
; 
32'd191982: dataIn1 = 32'd10692
; 
32'd191983: dataIn1 = 32'd10693
; 
32'd191984: dataIn1 = 32'd10694
; 
32'd191985: dataIn1 = 32'd1477
; 
32'd191986: dataIn1 = 32'd10693
; 
32'd191987: dataIn1 = 32'd10694
; 
32'd191988: dataIn1 = 32'd10695
; 
32'd191989: dataIn1 = 32'd1473
; 
32'd191990: dataIn1 = 32'd1477
; 
32'd191991: dataIn1 = 32'd10694
; 
32'd191992: dataIn1 = 32'd10695
; 
32'd191993: dataIn1 = 32'd10696
; 
32'd191994: dataIn1 = 32'd1473
; 
32'd191995: dataIn1 = 32'd10695
; 
32'd191996: dataIn1 = 32'd10696
; 
32'd191997: dataIn1 = 32'd10697
; 
32'd191998: dataIn1 = 32'd1472
; 
32'd191999: dataIn1 = 32'd1473
; 
32'd192000: dataIn1 = 32'd10696
; 
32'd192001: dataIn1 = 32'd10697
; 
32'd192002: dataIn1 = 32'd10698
; 
32'd192003: dataIn1 = 32'd1472
; 
32'd192004: dataIn1 = 32'd1480
; 
32'd192005: dataIn1 = 32'd10697
; 
32'd192006: dataIn1 = 32'd10698
; 
32'd192007: dataIn1 = 32'd10699
; 
32'd192008: dataIn1 = 32'd1480
; 
32'd192009: dataIn1 = 32'd10698
; 
32'd192010: dataIn1 = 32'd10699
; 
32'd192011: dataIn1 = 32'd10700
; 
32'd192012: dataIn1 = 32'd1480
; 
32'd192013: dataIn1 = 32'd10699
; 
32'd192014: dataIn1 = 32'd10700
; 
32'd192015: dataIn1 = 32'd10701
; 
32'd192016: dataIn1 = 32'd1479
; 
32'd192017: dataIn1 = 32'd1480
; 
32'd192018: dataIn1 = 32'd10700
; 
32'd192019: dataIn1 = 32'd10701
; 
32'd192020: dataIn1 = 32'd10702
; 
32'd192021: dataIn1 = 32'd1479
; 
32'd192022: dataIn1 = 32'd10701
; 
32'd192023: dataIn1 = 32'd10702
; 
32'd192024: dataIn1 = 32'd10703
; 
32'd192025: dataIn1 = 32'd1448
; 
32'd192026: dataIn1 = 32'd1479
; 
32'd192027: dataIn1 = 32'd10702
; 
32'd192028: dataIn1 = 32'd10703
; 
32'd192029: dataIn1 = 32'd10704
; 
32'd192030: dataIn1 = 32'd1446
; 
32'd192031: dataIn1 = 32'd1448
; 
32'd192032: dataIn1 = 32'd10703
; 
32'd192033: dataIn1 = 32'd10704
; 
32'd192034: dataIn1 = 32'd10705
; 
32'd192035: dataIn1 = 32'd1446
; 
32'd192036: dataIn1 = 32'd10704
; 
32'd192037: dataIn1 = 32'd10705
; 
32'd192038: dataIn1 = 32'd10706
; 
32'd192039: dataIn1 = 32'd1446
; 
32'd192040: dataIn1 = 32'd10538
; 
32'd192041: dataIn1 = 32'd10705
; 
32'd192042: dataIn1 = 32'd10706
; 
32'd192043: dataIn1 = 32'd743
; 
32'd192044: dataIn1 = 32'd1424
; 
32'd192045: dataIn1 = 32'd10561
; 
32'd192046: dataIn1 = 32'd10707
; 
32'd192047: dataIn1 = 32'd10708
; 
32'd192048: dataIn1 = 32'd11738
; 
32'd192049: dataIn1 = 32'd389
; 
32'd192050: dataIn1 = 32'd10561
; 
32'd192051: dataIn1 = 32'd10707
; 
32'd192052: dataIn1 = 32'd10708
; 
32'd192053: dataIn1 = 32'd10709
; 
32'd192054: dataIn1 = 32'd389
; 
32'd192055: dataIn1 = 32'd1425
; 
32'd192056: dataIn1 = 32'd10708
; 
32'd192057: dataIn1 = 32'd10709
; 
32'd192058: dataIn1 = 32'd10710
; 
32'd192059: dataIn1 = 32'd747
; 
32'd192060: dataIn1 = 32'd1425
; 
32'd192061: dataIn1 = 32'd10709
; 
32'd192062: dataIn1 = 32'd10710
; 
32'd192063: dataIn1 = 32'd10711
; 
32'd192064: dataIn1 = 32'd747
; 
32'd192065: dataIn1 = 32'd1426
; 
32'd192066: dataIn1 = 32'd10710
; 
32'd192067: dataIn1 = 32'd10711
; 
32'd192068: dataIn1 = 32'd10712
; 
32'd192069: dataIn1 = 32'd203
; 
32'd192070: dataIn1 = 32'd1426
; 
32'd192071: dataIn1 = 32'd10711
; 
32'd192072: dataIn1 = 32'd10712
; 
32'd192073: dataIn1 = 32'd10713
; 
32'd192074: dataIn1 = 32'd203
; 
32'd192075: dataIn1 = 32'd1416
; 
32'd192076: dataIn1 = 32'd10712
; 
32'd192077: dataIn1 = 32'd10713
; 
32'd192078: dataIn1 = 32'd10714
; 
32'd192079: dataIn1 = 32'd740
; 
32'd192080: dataIn1 = 32'd1416
; 
32'd192081: dataIn1 = 32'd10713
; 
32'd192082: dataIn1 = 32'd10714
; 
32'd192083: dataIn1 = 32'd10715
; 
32'd192084: dataIn1 = 32'd740
; 
32'd192085: dataIn1 = 32'd1415
; 
32'd192086: dataIn1 = 32'd10714
; 
32'd192087: dataIn1 = 32'd10715
; 
32'd192088: dataIn1 = 32'd10716
; 
32'd192089: dataIn1 = 32'd387
; 
32'd192090: dataIn1 = 32'd1415
; 
32'd192091: dataIn1 = 32'd10715
; 
32'd192092: dataIn1 = 32'd10716
; 
32'd192093: dataIn1 = 32'd10717
; 
32'd192094: dataIn1 = 32'd387
; 
32'd192095: dataIn1 = 32'd1414
; 
32'd192096: dataIn1 = 32'd10716
; 
32'd192097: dataIn1 = 32'd10717
; 
32'd192098: dataIn1 = 32'd10718
; 
32'd192099: dataIn1 = 32'd739
; 
32'd192100: dataIn1 = 32'd1414
; 
32'd192101: dataIn1 = 32'd10717
; 
32'd192102: dataIn1 = 32'd10718
; 
32'd192103: dataIn1 = 32'd10719
; 
32'd192104: dataIn1 = 32'd739
; 
32'd192105: dataIn1 = 32'd1413
; 
32'd192106: dataIn1 = 32'd10718
; 
32'd192107: dataIn1 = 32'd10719
; 
32'd192108: dataIn1 = 32'd10720
; 
32'd192109: dataIn1 = 32'd201
; 
32'd192110: dataIn1 = 32'd1413
; 
32'd192111: dataIn1 = 32'd10719
; 
32'd192112: dataIn1 = 32'd10720
; 
32'd192113: dataIn1 = 32'd10721
; 
32'd192114: dataIn1 = 32'd201
; 
32'd192115: dataIn1 = 32'd1417
; 
32'd192116: dataIn1 = 32'd10720
; 
32'd192117: dataIn1 = 32'd10721
; 
32'd192118: dataIn1 = 32'd10722
; 
32'd192119: dataIn1 = 32'd741
; 
32'd192120: dataIn1 = 32'd1417
; 
32'd192121: dataIn1 = 32'd10721
; 
32'd192122: dataIn1 = 32'd10722
; 
32'd192123: dataIn1 = 32'd10723
; 
32'd192124: dataIn1 = 32'd741
; 
32'd192125: dataIn1 = 32'd1418
; 
32'd192126: dataIn1 = 32'd10722
; 
32'd192127: dataIn1 = 32'd10723
; 
32'd192128: dataIn1 = 32'd10724
; 
32'd192129: dataIn1 = 32'd388
; 
32'd192130: dataIn1 = 32'd1418
; 
32'd192131: dataIn1 = 32'd10723
; 
32'd192132: dataIn1 = 32'd10724
; 
32'd192133: dataIn1 = 32'd10725
; 
32'd192134: dataIn1 = 32'd388
; 
32'd192135: dataIn1 = 32'd1420
; 
32'd192136: dataIn1 = 32'd10724
; 
32'd192137: dataIn1 = 32'd10725
; 
32'd192138: dataIn1 = 32'd10726
; 
32'd192139: dataIn1 = 32'd742
; 
32'd192140: dataIn1 = 32'd1420
; 
32'd192141: dataIn1 = 32'd10725
; 
32'd192142: dataIn1 = 32'd10726
; 
32'd192143: dataIn1 = 32'd10727
; 
32'd192144: dataIn1 = 32'd742
; 
32'd192145: dataIn1 = 32'd1419
; 
32'd192146: dataIn1 = 32'd10726
; 
32'd192147: dataIn1 = 32'd10727
; 
32'd192148: dataIn1 = 32'd10728
; 
32'd192149: dataIn1 = 32'd200
; 
32'd192150: dataIn1 = 32'd1419
; 
32'd192151: dataIn1 = 32'd10727
; 
32'd192152: dataIn1 = 32'd10728
; 
32'd192153: dataIn1 = 32'd10729
; 
32'd192154: dataIn1 = 32'd200
; 
32'd192155: dataIn1 = 32'd1412
; 
32'd192156: dataIn1 = 32'd10728
; 
32'd192157: dataIn1 = 32'd10729
; 
32'd192158: dataIn1 = 32'd10730
; 
32'd192159: dataIn1 = 32'd738
; 
32'd192160: dataIn1 = 32'd1412
; 
32'd192161: dataIn1 = 32'd10729
; 
32'd192162: dataIn1 = 32'd10730
; 
32'd192163: dataIn1 = 32'd10731
; 
32'd192164: dataIn1 = 32'd738
; 
32'd192165: dataIn1 = 32'd1411
; 
32'd192166: dataIn1 = 32'd10730
; 
32'd192167: dataIn1 = 32'd10731
; 
32'd192168: dataIn1 = 32'd10732
; 
32'd192169: dataIn1 = 32'd386
; 
32'd192170: dataIn1 = 32'd1411
; 
32'd192171: dataIn1 = 32'd10731
; 
32'd192172: dataIn1 = 32'd10732
; 
32'd192173: dataIn1 = 32'd10733
; 
32'd192174: dataIn1 = 32'd386
; 
32'd192175: dataIn1 = 32'd1409
; 
32'd192176: dataIn1 = 32'd10732
; 
32'd192177: dataIn1 = 32'd10733
; 
32'd192178: dataIn1 = 32'd10734
; 
32'd192179: dataIn1 = 32'd737
; 
32'd192180: dataIn1 = 32'd1409
; 
32'd192181: dataIn1 = 32'd10733
; 
32'd192182: dataIn1 = 32'd10734
; 
32'd192183: dataIn1 = 32'd10735
; 
32'd192184: dataIn1 = 32'd737
; 
32'd192185: dataIn1 = 32'd1410
; 
32'd192186: dataIn1 = 32'd10734
; 
32'd192187: dataIn1 = 32'd10735
; 
32'd192188: dataIn1 = 32'd10736
; 
32'd192189: dataIn1 = 32'd198
; 
32'd192190: dataIn1 = 32'd1410
; 
32'd192191: dataIn1 = 32'd10735
; 
32'd192192: dataIn1 = 32'd10736
; 
32'd192193: dataIn1 = 32'd10737
; 
32'd192194: dataIn1 = 32'd198
; 
32'd192195: dataIn1 = 32'd1406
; 
32'd192196: dataIn1 = 32'd10736
; 
32'd192197: dataIn1 = 32'd10737
; 
32'd192198: dataIn1 = 32'd10738
; 
32'd192199: dataIn1 = 32'd735
; 
32'd192200: dataIn1 = 32'd1406
; 
32'd192201: dataIn1 = 32'd10737
; 
32'd192202: dataIn1 = 32'd10738
; 
32'd192203: dataIn1 = 32'd10739
; 
32'd192204: dataIn1 = 32'd735
; 
32'd192205: dataIn1 = 32'd1405
; 
32'd192206: dataIn1 = 32'd10738
; 
32'd192207: dataIn1 = 32'd10739
; 
32'd192208: dataIn1 = 32'd10740
; 
32'd192209: dataIn1 = 32'd385
; 
32'd192210: dataIn1 = 32'd1405
; 
32'd192211: dataIn1 = 32'd10739
; 
32'd192212: dataIn1 = 32'd10740
; 
32'd192213: dataIn1 = 32'd10741
; 
32'd192214: dataIn1 = 32'd385
; 
32'd192215: dataIn1 = 32'd1407
; 
32'd192216: dataIn1 = 32'd10740
; 
32'd192217: dataIn1 = 32'd10741
; 
32'd192218: dataIn1 = 32'd10742
; 
32'd192219: dataIn1 = 32'd736
; 
32'd192220: dataIn1 = 32'd1407
; 
32'd192221: dataIn1 = 32'd10741
; 
32'd192222: dataIn1 = 32'd10742
; 
32'd192223: dataIn1 = 32'd10743
; 
32'd192224: dataIn1 = 32'd736
; 
32'd192225: dataIn1 = 32'd1408
; 
32'd192226: dataIn1 = 32'd10742
; 
32'd192227: dataIn1 = 32'd10743
; 
32'd192228: dataIn1 = 32'd10744
; 
32'd192229: dataIn1 = 32'd196
; 
32'd192230: dataIn1 = 32'd1408
; 
32'd192231: dataIn1 = 32'd10743
; 
32'd192232: dataIn1 = 32'd10744
; 
32'd192233: dataIn1 = 32'd10745
; 
32'd192234: dataIn1 = 32'd196
; 
32'd192235: dataIn1 = 32'd1400
; 
32'd192236: dataIn1 = 32'd10744
; 
32'd192237: dataIn1 = 32'd10745
; 
32'd192238: dataIn1 = 32'd10746
; 
32'd192239: dataIn1 = 32'd732
; 
32'd192240: dataIn1 = 32'd1400
; 
32'd192241: dataIn1 = 32'd10745
; 
32'd192242: dataIn1 = 32'd10746
; 
32'd192243: dataIn1 = 32'd10747
; 
32'd192244: dataIn1 = 32'd732
; 
32'd192245: dataIn1 = 32'd1399
; 
32'd192246: dataIn1 = 32'd10746
; 
32'd192247: dataIn1 = 32'd10747
; 
32'd192248: dataIn1 = 32'd10748
; 
32'd192249: dataIn1 = 32'd383
; 
32'd192250: dataIn1 = 32'd1399
; 
32'd192251: dataIn1 = 32'd10747
; 
32'd192252: dataIn1 = 32'd10748
; 
32'd192253: dataIn1 = 32'd10749
; 
32'd192254: dataIn1 = 32'd383
; 
32'd192255: dataIn1 = 32'd1398
; 
32'd192256: dataIn1 = 32'd10748
; 
32'd192257: dataIn1 = 32'd10749
; 
32'd192258: dataIn1 = 32'd10750
; 
32'd192259: dataIn1 = 32'd731
; 
32'd192260: dataIn1 = 32'd1398
; 
32'd192261: dataIn1 = 32'd10749
; 
32'd192262: dataIn1 = 32'd10750
; 
32'd192263: dataIn1 = 32'd10751
; 
32'd192264: dataIn1 = 32'd731
; 
32'd192265: dataIn1 = 32'd1397
; 
32'd192266: dataIn1 = 32'd10750
; 
32'd192267: dataIn1 = 32'd10751
; 
32'd192268: dataIn1 = 32'd10752
; 
32'd192269: dataIn1 = 32'd1397
; 
32'd192270: dataIn1 = 32'd10751
; 
32'd192271: dataIn1 = 32'd10752
; 
32'd192272: dataIn1 = 32'd10753
; 
32'd192273: dataIn1 = 32'd194
; 
32'd192274: dataIn1 = 32'd1397
; 
32'd192275: dataIn1 = 32'd10752
; 
32'd192276: dataIn1 = 32'd10753
; 
32'd192277: dataIn1 = 32'd10754
; 
32'd192278: dataIn1 = 32'd194
; 
32'd192279: dataIn1 = 32'd733
; 
32'd192280: dataIn1 = 32'd1401
; 
32'd192281: dataIn1 = 32'd10753
; 
32'd192282: dataIn1 = 32'd10754
; 
32'd192283: dataIn1 = 32'd10755
; 
32'd192284: dataIn1 = 32'd733
; 
32'd192285: dataIn1 = 32'd1402
; 
32'd192286: dataIn1 = 32'd10754
; 
32'd192287: dataIn1 = 32'd10755
; 
32'd192288: dataIn1 = 32'd10756
; 
32'd192289: dataIn1 = 32'd1402
; 
32'd192290: dataIn1 = 32'd10755
; 
32'd192291: dataIn1 = 32'd10756
; 
32'd192292: dataIn1 = 32'd10757
; 
32'd192293: dataIn1 = 32'd384
; 
32'd192294: dataIn1 = 32'd1402
; 
32'd192295: dataIn1 = 32'd10756
; 
32'd192296: dataIn1 = 32'd10757
; 
32'd192297: dataIn1 = 32'd10758
; 
32'd192298: dataIn1 = 32'd384
; 
32'd192299: dataIn1 = 32'd1404
; 
32'd192300: dataIn1 = 32'd10757
; 
32'd192301: dataIn1 = 32'd10758
; 
32'd192302: dataIn1 = 32'd10759
; 
32'd192303: dataIn1 = 32'd734
; 
32'd192304: dataIn1 = 32'd1404
; 
32'd192305: dataIn1 = 32'd10758
; 
32'd192306: dataIn1 = 32'd10759
; 
32'd192307: dataIn1 = 32'd10760
; 
32'd192308: dataIn1 = 32'd197
; 
32'd192309: dataIn1 = 32'd734
; 
32'd192310: dataIn1 = 32'd1403
; 
32'd192311: dataIn1 = 32'd10759
; 
32'd192312: dataIn1 = 32'd10760
; 
32'd192313: dataIn1 = 32'd10761
; 
32'd192314: dataIn1 = 32'd197
; 
32'd192315: dataIn1 = 32'd10760
; 
32'd192316: dataIn1 = 32'd10761
; 
32'd192317: dataIn1 = 32'd953
; 
32'd192318: dataIn1 = 32'd1719
; 
32'd192319: dataIn1 = 32'd10562
; 
32'd192320: dataIn1 = 32'd10762
; 
32'd192321: dataIn1 = 32'd10763
; 
32'd192322: dataIn1 = 32'd953
; 
32'd192323: dataIn1 = 32'd10762
; 
32'd192324: dataIn1 = 32'd10763
; 
32'd192325: dataIn1 = 32'd10764
; 
32'd192326: dataIn1 = 32'd953
; 
32'd192327: dataIn1 = 32'd1712
; 
32'd192328: dataIn1 = 32'd10763
; 
32'd192329: dataIn1 = 32'd10764
; 
32'd192330: dataIn1 = 32'd10765
; 
32'd192331: dataIn1 = 32'd951
; 
32'd192332: dataIn1 = 32'd1712
; 
32'd192333: dataIn1 = 32'd10764
; 
32'd192334: dataIn1 = 32'd10765
; 
32'd192335: dataIn1 = 32'd10766
; 
32'd192336: dataIn1 = 32'd951
; 
32'd192337: dataIn1 = 32'd1711
; 
32'd192338: dataIn1 = 32'd10765
; 
32'd192339: dataIn1 = 32'd10766
; 
32'd192340: dataIn1 = 32'd10767
; 
32'd192341: dataIn1 = 32'd952
; 
32'd192342: dataIn1 = 32'd1711
; 
32'd192343: dataIn1 = 32'd10766
; 
32'd192344: dataIn1 = 32'd10767
; 
32'd192345: dataIn1 = 32'd10768
; 
32'd192346: dataIn1 = 32'd952
; 
32'd192347: dataIn1 = 32'd1715
; 
32'd192348: dataIn1 = 32'd10767
; 
32'd192349: dataIn1 = 32'd10768
; 
32'd192350: dataIn1 = 32'd10769
; 
32'd192351: dataIn1 = 32'd955
; 
32'd192352: dataIn1 = 32'd1715
; 
32'd192353: dataIn1 = 32'd10768
; 
32'd192354: dataIn1 = 32'd10769
; 
32'd192355: dataIn1 = 32'd10770
; 
32'd192356: dataIn1 = 32'd955
; 
32'd192357: dataIn1 = 32'd1718
; 
32'd192358: dataIn1 = 32'd10769
; 
32'd192359: dataIn1 = 32'd10770
; 
32'd192360: dataIn1 = 32'd10771
; 
32'd192361: dataIn1 = 32'd944
; 
32'd192362: dataIn1 = 32'd1718
; 
32'd192363: dataIn1 = 32'd10770
; 
32'd192364: dataIn1 = 32'd10771
; 
32'd192365: dataIn1 = 32'd10772
; 
32'd192366: dataIn1 = 32'd944
; 
32'd192367: dataIn1 = 32'd1699
; 
32'd192368: dataIn1 = 32'd10771
; 
32'd192369: dataIn1 = 32'd10772
; 
32'd192370: dataIn1 = 32'd10773
; 
32'd192371: dataIn1 = 32'd940
; 
32'd192372: dataIn1 = 32'd1699
; 
32'd192373: dataIn1 = 32'd10772
; 
32'd192374: dataIn1 = 32'd10773
; 
32'd192375: dataIn1 = 32'd10774
; 
32'd192376: dataIn1 = 32'd940
; 
32'd192377: dataIn1 = 32'd1695
; 
32'd192378: dataIn1 = 32'd10773
; 
32'd192379: dataIn1 = 32'd10774
; 
32'd192380: dataIn1 = 32'd10775
; 
32'd192381: dataIn1 = 32'd939
; 
32'd192382: dataIn1 = 32'd1695
; 
32'd192383: dataIn1 = 32'd10774
; 
32'd192384: dataIn1 = 32'd10775
; 
32'd192385: dataIn1 = 32'd10776
; 
32'd192386: dataIn1 = 32'd939
; 
32'd192387: dataIn1 = 32'd1696
; 
32'd192388: dataIn1 = 32'd10775
; 
32'd192389: dataIn1 = 32'd10776
; 
32'd192390: dataIn1 = 32'd10777
; 
32'd192391: dataIn1 = 32'd941
; 
32'd192392: dataIn1 = 32'd1696
; 
32'd192393: dataIn1 = 32'd10776
; 
32'd192394: dataIn1 = 32'd10777
; 
32'd192395: dataIn1 = 32'd10778
; 
32'd192396: dataIn1 = 32'd941
; 
32'd192397: dataIn1 = 32'd1710
; 
32'd192398: dataIn1 = 32'd10777
; 
32'd192399: dataIn1 = 32'd10778
; 
32'd192400: dataIn1 = 32'd10779
; 
32'd192401: dataIn1 = 32'd948
; 
32'd192402: dataIn1 = 32'd1710
; 
32'd192403: dataIn1 = 32'd10778
; 
32'd192404: dataIn1 = 32'd10779
; 
32'd192405: dataIn1 = 32'd10780
; 
32'd192406: dataIn1 = 32'd948
; 
32'd192407: dataIn1 = 32'd1703
; 
32'd192408: dataIn1 = 32'd10779
; 
32'd192409: dataIn1 = 32'd10780
; 
32'd192410: dataIn1 = 32'd10781
; 
32'd192411: dataIn1 = 32'd945
; 
32'd192412: dataIn1 = 32'd1703
; 
32'd192413: dataIn1 = 32'd10780
; 
32'd192414: dataIn1 = 32'd10781
; 
32'd192415: dataIn1 = 32'd10782
; 
32'd192416: dataIn1 = 32'd945
; 
32'd192417: dataIn1 = 32'd1702
; 
32'd192418: dataIn1 = 32'd10781
; 
32'd192419: dataIn1 = 32'd10782
; 
32'd192420: dataIn1 = 32'd10783
; 
32'd192421: dataIn1 = 32'd946
; 
32'd192422: dataIn1 = 32'd1702
; 
32'd192423: dataIn1 = 32'd10782
; 
32'd192424: dataIn1 = 32'd10783
; 
32'd192425: dataIn1 = 32'd10784
; 
32'd192426: dataIn1 = 32'd946
; 
32'd192427: dataIn1 = 32'd1706
; 
32'd192428: dataIn1 = 32'd10783
; 
32'd192429: dataIn1 = 32'd10784
; 
32'd192430: dataIn1 = 32'd10785
; 
32'd192431: dataIn1 = 32'd950
; 
32'd192432: dataIn1 = 32'd1706
; 
32'd192433: dataIn1 = 32'd10784
; 
32'd192434: dataIn1 = 32'd10785
; 
32'd192435: dataIn1 = 32'd10786
; 
32'd192436: dataIn1 = 32'd950
; 
32'd192437: dataIn1 = 32'd1709
; 
32'd192438: dataIn1 = 32'd10785
; 
32'd192439: dataIn1 = 32'd10786
; 
32'd192440: dataIn1 = 32'd10787
; 
32'd192441: dataIn1 = 32'd937
; 
32'd192442: dataIn1 = 32'd1709
; 
32'd192443: dataIn1 = 32'd10786
; 
32'd192444: dataIn1 = 32'd10787
; 
32'd192445: dataIn1 = 32'd10788
; 
32'd192446: dataIn1 = 32'd937
; 
32'd192447: dataIn1 = 32'd1692
; 
32'd192448: dataIn1 = 32'd10787
; 
32'd192449: dataIn1 = 32'd10788
; 
32'd192450: dataIn1 = 32'd10789
; 
32'd192451: dataIn1 = 32'd935
; 
32'd192452: dataIn1 = 32'd1692
; 
32'd192453: dataIn1 = 32'd10788
; 
32'd192454: dataIn1 = 32'd10789
; 
32'd192455: dataIn1 = 32'd10790
; 
32'd192456: dataIn1 = 32'd935
; 
32'd192457: dataIn1 = 32'd1688
; 
32'd192458: dataIn1 = 32'd10789
; 
32'd192459: dataIn1 = 32'd10790
; 
32'd192460: dataIn1 = 32'd10791
; 
32'd192461: dataIn1 = 32'd934
; 
32'd192462: dataIn1 = 32'd1688
; 
32'd192463: dataIn1 = 32'd10790
; 
32'd192464: dataIn1 = 32'd10791
; 
32'd192465: dataIn1 = 32'd10792
; 
32'd192466: dataIn1 = 32'd934
; 
32'd192467: dataIn1 = 32'd1689
; 
32'd192468: dataIn1 = 32'd10791
; 
32'd192469: dataIn1 = 32'd10792
; 
32'd192470: dataIn1 = 32'd10793
; 
32'd192471: dataIn1 = 32'd933
; 
32'd192472: dataIn1 = 32'd1689
; 
32'd192473: dataIn1 = 32'd10792
; 
32'd192474: dataIn1 = 32'd10793
; 
32'd192475: dataIn1 = 32'd10794
; 
32'd192476: dataIn1 = 32'd933
; 
32'd192477: dataIn1 = 32'd1687
; 
32'd192478: dataIn1 = 32'd10793
; 
32'd192479: dataIn1 = 32'd10794
; 
32'd192480: dataIn1 = 32'd10795
; 
32'd192481: dataIn1 = 32'd929
; 
32'd192482: dataIn1 = 32'd1687
; 
32'd192483: dataIn1 = 32'd10794
; 
32'd192484: dataIn1 = 32'd10795
; 
32'd192485: dataIn1 = 32'd10796
; 
32'd192486: dataIn1 = 32'd929
; 
32'd192487: dataIn1 = 32'd1680
; 
32'd192488: dataIn1 = 32'd10795
; 
32'd192489: dataIn1 = 32'd10796
; 
32'd192490: dataIn1 = 32'd10797
; 
32'd192491: dataIn1 = 32'd927
; 
32'd192492: dataIn1 = 32'd1680
; 
32'd192493: dataIn1 = 32'd10796
; 
32'd192494: dataIn1 = 32'd10797
; 
32'd192495: dataIn1 = 32'd10798
; 
32'd192496: dataIn1 = 32'd927
; 
32'd192497: dataIn1 = 32'd1679
; 
32'd192498: dataIn1 = 32'd10797
; 
32'd192499: dataIn1 = 32'd10798
; 
32'd192500: dataIn1 = 32'd10799
; 
32'd192501: dataIn1 = 32'd928
; 
32'd192502: dataIn1 = 32'd1679
; 
32'd192503: dataIn1 = 32'd10798
; 
32'd192504: dataIn1 = 32'd10799
; 
32'd192505: dataIn1 = 32'd10800
; 
32'd192506: dataIn1 = 32'd928
; 
32'd192507: dataIn1 = 32'd1683
; 
32'd192508: dataIn1 = 32'd10799
; 
32'd192509: dataIn1 = 32'd10800
; 
32'd192510: dataIn1 = 32'd10801
; 
32'd192511: dataIn1 = 32'd931
; 
32'd192512: dataIn1 = 32'd1683
; 
32'd192513: dataIn1 = 32'd10800
; 
32'd192514: dataIn1 = 32'd10801
; 
32'd192515: dataIn1 = 32'd10802
; 
32'd192516: dataIn1 = 32'd931
; 
32'd192517: dataIn1 = 32'd1686
; 
32'd192518: dataIn1 = 32'd10801
; 
32'd192519: dataIn1 = 32'd10802
; 
32'd192520: dataIn1 = 32'd10803
; 
32'd192521: dataIn1 = 32'd920
; 
32'd192522: dataIn1 = 32'd1686
; 
32'd192523: dataIn1 = 32'd10802
; 
32'd192524: dataIn1 = 32'd10803
; 
32'd192525: dataIn1 = 32'd10804
; 
32'd192526: dataIn1 = 32'd920
; 
32'd192527: dataIn1 = 32'd1667
; 
32'd192528: dataIn1 = 32'd10803
; 
32'd192529: dataIn1 = 32'd10804
; 
32'd192530: dataIn1 = 32'd10805
; 
32'd192531: dataIn1 = 32'd916
; 
32'd192532: dataIn1 = 32'd1667
; 
32'd192533: dataIn1 = 32'd10804
; 
32'd192534: dataIn1 = 32'd10805
; 
32'd192535: dataIn1 = 32'd10806
; 
32'd192536: dataIn1 = 32'd916
; 
32'd192537: dataIn1 = 32'd1663
; 
32'd192538: dataIn1 = 32'd10805
; 
32'd192539: dataIn1 = 32'd10806
; 
32'd192540: dataIn1 = 32'd10807
; 
32'd192541: dataIn1 = 32'd915
; 
32'd192542: dataIn1 = 32'd1663
; 
32'd192543: dataIn1 = 32'd10806
; 
32'd192544: dataIn1 = 32'd10807
; 
32'd192545: dataIn1 = 32'd10808
; 
32'd192546: dataIn1 = 32'd915
; 
32'd192547: dataIn1 = 32'd1664
; 
32'd192548: dataIn1 = 32'd10807
; 
32'd192549: dataIn1 = 32'd10808
; 
32'd192550: dataIn1 = 32'd10809
; 
32'd192551: dataIn1 = 32'd917
; 
32'd192552: dataIn1 = 32'd1664
; 
32'd192553: dataIn1 = 32'd10808
; 
32'd192554: dataIn1 = 32'd10809
; 
32'd192555: dataIn1 = 32'd10810
; 
32'd192556: dataIn1 = 32'd917
; 
32'd192557: dataIn1 = 32'd1678
; 
32'd192558: dataIn1 = 32'd10809
; 
32'd192559: dataIn1 = 32'd10810
; 
32'd192560: dataIn1 = 32'd10811
; 
32'd192561: dataIn1 = 32'd924
; 
32'd192562: dataIn1 = 32'd1678
; 
32'd192563: dataIn1 = 32'd10810
; 
32'd192564: dataIn1 = 32'd10811
; 
32'd192565: dataIn1 = 32'd10812
; 
32'd192566: dataIn1 = 32'd924
; 
32'd192567: dataIn1 = 32'd1671
; 
32'd192568: dataIn1 = 32'd10811
; 
32'd192569: dataIn1 = 32'd10812
; 
32'd192570: dataIn1 = 32'd10813
; 
32'd192571: dataIn1 = 32'd921
; 
32'd192572: dataIn1 = 32'd1671
; 
32'd192573: dataIn1 = 32'd10812
; 
32'd192574: dataIn1 = 32'd10813
; 
32'd192575: dataIn1 = 32'd10814
; 
32'd192576: dataIn1 = 32'd921
; 
32'd192577: dataIn1 = 32'd1670
; 
32'd192578: dataIn1 = 32'd10813
; 
32'd192579: dataIn1 = 32'd10814
; 
32'd192580: dataIn1 = 32'd10815
; 
32'd192581: dataIn1 = 32'd922
; 
32'd192582: dataIn1 = 32'd1670
; 
32'd192583: dataIn1 = 32'd10814
; 
32'd192584: dataIn1 = 32'd10815
; 
32'd192585: dataIn1 = 32'd10816
; 
32'd192586: dataIn1 = 32'd922
; 
32'd192587: dataIn1 = 32'd1674
; 
32'd192588: dataIn1 = 32'd10815
; 
32'd192589: dataIn1 = 32'd10816
; 
32'd192590: dataIn1 = 32'd10817
; 
32'd192591: dataIn1 = 32'd926
; 
32'd192592: dataIn1 = 32'd1674
; 
32'd192593: dataIn1 = 32'd10816
; 
32'd192594: dataIn1 = 32'd10817
; 
32'd192595: dataIn1 = 32'd10818
; 
32'd192596: dataIn1 = 32'd926
; 
32'd192597: dataIn1 = 32'd1677
; 
32'd192598: dataIn1 = 32'd10817
; 
32'd192599: dataIn1 = 32'd10818
; 
32'd192600: dataIn1 = 32'd10819
; 
32'd192601: dataIn1 = 32'd913
; 
32'd192602: dataIn1 = 32'd1677
; 
32'd192603: dataIn1 = 32'd10818
; 
32'd192604: dataIn1 = 32'd10819
; 
32'd192605: dataIn1 = 32'd10820
; 
32'd192606: dataIn1 = 32'd913
; 
32'd192607: dataIn1 = 32'd1660
; 
32'd192608: dataIn1 = 32'd10819
; 
32'd192609: dataIn1 = 32'd10820
; 
32'd192610: dataIn1 = 32'd10821
; 
32'd192611: dataIn1 = 32'd911
; 
32'd192612: dataIn1 = 32'd1660
; 
32'd192613: dataIn1 = 32'd10820
; 
32'd192614: dataIn1 = 32'd10821
; 
32'd192615: dataIn1 = 32'd10822
; 
32'd192616: dataIn1 = 32'd911
; 
32'd192617: dataIn1 = 32'd1656
; 
32'd192618: dataIn1 = 32'd10821
; 
32'd192619: dataIn1 = 32'd10822
; 
32'd192620: dataIn1 = 32'd10823
; 
32'd192621: dataIn1 = 32'd910
; 
32'd192622: dataIn1 = 32'd1656
; 
32'd192623: dataIn1 = 32'd10822
; 
32'd192624: dataIn1 = 32'd10823
; 
32'd192625: dataIn1 = 32'd10824
; 
32'd192626: dataIn1 = 32'd910
; 
32'd192627: dataIn1 = 32'd1657
; 
32'd192628: dataIn1 = 32'd10823
; 
32'd192629: dataIn1 = 32'd10824
; 
32'd192630: dataIn1 = 32'd10825
; 
32'd192631: dataIn1 = 32'd909
; 
32'd192632: dataIn1 = 32'd1657
; 
32'd192633: dataIn1 = 32'd10824
; 
32'd192634: dataIn1 = 32'd10825
; 
32'd192635: dataIn1 = 32'd10826
; 
32'd192636: dataIn1 = 32'd909
; 
32'd192637: dataIn1 = 32'd1655
; 
32'd192638: dataIn1 = 32'd10825
; 
32'd192639: dataIn1 = 32'd10826
; 
32'd192640: dataIn1 = 32'd10827
; 
32'd192641: dataIn1 = 32'd905
; 
32'd192642: dataIn1 = 32'd1655
; 
32'd192643: dataIn1 = 32'd10826
; 
32'd192644: dataIn1 = 32'd10827
; 
32'd192645: dataIn1 = 32'd10828
; 
32'd192646: dataIn1 = 32'd905
; 
32'd192647: dataIn1 = 32'd1648
; 
32'd192648: dataIn1 = 32'd10827
; 
32'd192649: dataIn1 = 32'd10828
; 
32'd192650: dataIn1 = 32'd10829
; 
32'd192651: dataIn1 = 32'd903
; 
32'd192652: dataIn1 = 32'd1648
; 
32'd192653: dataIn1 = 32'd10828
; 
32'd192654: dataIn1 = 32'd10829
; 
32'd192655: dataIn1 = 32'd10830
; 
32'd192656: dataIn1 = 32'd903
; 
32'd192657: dataIn1 = 32'd1647
; 
32'd192658: dataIn1 = 32'd10829
; 
32'd192659: dataIn1 = 32'd10830
; 
32'd192660: dataIn1 = 32'd10831
; 
32'd192661: dataIn1 = 32'd904
; 
32'd192662: dataIn1 = 32'd1647
; 
32'd192663: dataIn1 = 32'd10830
; 
32'd192664: dataIn1 = 32'd10831
; 
32'd192665: dataIn1 = 32'd10832
; 
32'd192666: dataIn1 = 32'd904
; 
32'd192667: dataIn1 = 32'd1651
; 
32'd192668: dataIn1 = 32'd10831
; 
32'd192669: dataIn1 = 32'd10832
; 
32'd192670: dataIn1 = 32'd10833
; 
32'd192671: dataIn1 = 32'd907
; 
32'd192672: dataIn1 = 32'd1651
; 
32'd192673: dataIn1 = 32'd10832
; 
32'd192674: dataIn1 = 32'd10833
; 
32'd192675: dataIn1 = 32'd10834
; 
32'd192676: dataIn1 = 32'd907
; 
32'd192677: dataIn1 = 32'd1654
; 
32'd192678: dataIn1 = 32'd10833
; 
32'd192679: dataIn1 = 32'd10834
; 
32'd192680: dataIn1 = 32'd10835
; 
32'd192681: dataIn1 = 32'd896
; 
32'd192682: dataIn1 = 32'd1654
; 
32'd192683: dataIn1 = 32'd10834
; 
32'd192684: dataIn1 = 32'd10835
; 
32'd192685: dataIn1 = 32'd10836
; 
32'd192686: dataIn1 = 32'd896
; 
32'd192687: dataIn1 = 32'd1635
; 
32'd192688: dataIn1 = 32'd10835
; 
32'd192689: dataIn1 = 32'd10836
; 
32'd192690: dataIn1 = 32'd10837
; 
32'd192691: dataIn1 = 32'd892
; 
32'd192692: dataIn1 = 32'd1635
; 
32'd192693: dataIn1 = 32'd10836
; 
32'd192694: dataIn1 = 32'd10837
; 
32'd192695: dataIn1 = 32'd10838
; 
32'd192696: dataIn1 = 32'd892
; 
32'd192697: dataIn1 = 32'd1631
; 
32'd192698: dataIn1 = 32'd10837
; 
32'd192699: dataIn1 = 32'd10838
; 
32'd192700: dataIn1 = 32'd10839
; 
32'd192701: dataIn1 = 32'd891
; 
32'd192702: dataIn1 = 32'd1631
; 
32'd192703: dataIn1 = 32'd10838
; 
32'd192704: dataIn1 = 32'd10839
; 
32'd192705: dataIn1 = 32'd10840
; 
32'd192706: dataIn1 = 32'd891
; 
32'd192707: dataIn1 = 32'd1632
; 
32'd192708: dataIn1 = 32'd10839
; 
32'd192709: dataIn1 = 32'd10840
; 
32'd192710: dataIn1 = 32'd10841
; 
32'd192711: dataIn1 = 32'd893
; 
32'd192712: dataIn1 = 32'd1632
; 
32'd192713: dataIn1 = 32'd10840
; 
32'd192714: dataIn1 = 32'd10841
; 
32'd192715: dataIn1 = 32'd10842
; 
32'd192716: dataIn1 = 32'd893
; 
32'd192717: dataIn1 = 32'd1646
; 
32'd192718: dataIn1 = 32'd10841
; 
32'd192719: dataIn1 = 32'd10842
; 
32'd192720: dataIn1 = 32'd10843
; 
32'd192721: dataIn1 = 32'd900
; 
32'd192722: dataIn1 = 32'd1646
; 
32'd192723: dataIn1 = 32'd10842
; 
32'd192724: dataIn1 = 32'd10843
; 
32'd192725: dataIn1 = 32'd10844
; 
32'd192726: dataIn1 = 32'd900
; 
32'd192727: dataIn1 = 32'd1639
; 
32'd192728: dataIn1 = 32'd10843
; 
32'd192729: dataIn1 = 32'd10844
; 
32'd192730: dataIn1 = 32'd10845
; 
32'd192731: dataIn1 = 32'd897
; 
32'd192732: dataIn1 = 32'd1639
; 
32'd192733: dataIn1 = 32'd10844
; 
32'd192734: dataIn1 = 32'd10845
; 
32'd192735: dataIn1 = 32'd10846
; 
32'd192736: dataIn1 = 32'd897
; 
32'd192737: dataIn1 = 32'd1638
; 
32'd192738: dataIn1 = 32'd10845
; 
32'd192739: dataIn1 = 32'd10846
; 
32'd192740: dataIn1 = 32'd10847
; 
32'd192741: dataIn1 = 32'd898
; 
32'd192742: dataIn1 = 32'd1638
; 
32'd192743: dataIn1 = 32'd10846
; 
32'd192744: dataIn1 = 32'd10847
; 
32'd192745: dataIn1 = 32'd10848
; 
32'd192746: dataIn1 = 32'd898
; 
32'd192747: dataIn1 = 32'd1642
; 
32'd192748: dataIn1 = 32'd10847
; 
32'd192749: dataIn1 = 32'd10848
; 
32'd192750: dataIn1 = 32'd10849
; 
32'd192751: dataIn1 = 32'd902
; 
32'd192752: dataIn1 = 32'd1642
; 
32'd192753: dataIn1 = 32'd10848
; 
32'd192754: dataIn1 = 32'd10849
; 
32'd192755: dataIn1 = 32'd10850
; 
32'd192756: dataIn1 = 32'd902
; 
32'd192757: dataIn1 = 32'd1645
; 
32'd192758: dataIn1 = 32'd10849
; 
32'd192759: dataIn1 = 32'd10850
; 
32'd192760: dataIn1 = 32'd10851
; 
32'd192761: dataIn1 = 32'd889
; 
32'd192762: dataIn1 = 32'd1645
; 
32'd192763: dataIn1 = 32'd10850
; 
32'd192764: dataIn1 = 32'd10851
; 
32'd192765: dataIn1 = 32'd10852
; 
32'd192766: dataIn1 = 32'd889
; 
32'd192767: dataIn1 = 32'd1628
; 
32'd192768: dataIn1 = 32'd10851
; 
32'd192769: dataIn1 = 32'd10852
; 
32'd192770: dataIn1 = 32'd10853
; 
32'd192771: dataIn1 = 32'd887
; 
32'd192772: dataIn1 = 32'd1628
; 
32'd192773: dataIn1 = 32'd10852
; 
32'd192774: dataIn1 = 32'd10853
; 
32'd192775: dataIn1 = 32'd10854
; 
32'd192776: dataIn1 = 32'd887
; 
32'd192777: dataIn1 = 32'd1624
; 
32'd192778: dataIn1 = 32'd10853
; 
32'd192779: dataIn1 = 32'd10854
; 
32'd192780: dataIn1 = 32'd10855
; 
32'd192781: dataIn1 = 32'd886
; 
32'd192782: dataIn1 = 32'd1624
; 
32'd192783: dataIn1 = 32'd10854
; 
32'd192784: dataIn1 = 32'd10855
; 
32'd192785: dataIn1 = 32'd10856
; 
32'd192786: dataIn1 = 32'd886
; 
32'd192787: dataIn1 = 32'd1625
; 
32'd192788: dataIn1 = 32'd10855
; 
32'd192789: dataIn1 = 32'd10856
; 
32'd192790: dataIn1 = 32'd10857
; 
32'd192791: dataIn1 = 32'd885
; 
32'd192792: dataIn1 = 32'd1625
; 
32'd192793: dataIn1 = 32'd10856
; 
32'd192794: dataIn1 = 32'd10857
; 
32'd192795: dataIn1 = 32'd10858
; 
32'd192796: dataIn1 = 32'd885
; 
32'd192797: dataIn1 = 32'd1623
; 
32'd192798: dataIn1 = 32'd10857
; 
32'd192799: dataIn1 = 32'd10858
; 
32'd192800: dataIn1 = 32'd10859
; 
32'd192801: dataIn1 = 32'd881
; 
32'd192802: dataIn1 = 32'd1623
; 
32'd192803: dataIn1 = 32'd10858
; 
32'd192804: dataIn1 = 32'd10859
; 
32'd192805: dataIn1 = 32'd10860
; 
32'd192806: dataIn1 = 32'd881
; 
32'd192807: dataIn1 = 32'd1616
; 
32'd192808: dataIn1 = 32'd10859
; 
32'd192809: dataIn1 = 32'd10860
; 
32'd192810: dataIn1 = 32'd10861
; 
32'd192811: dataIn1 = 32'd879
; 
32'd192812: dataIn1 = 32'd1616
; 
32'd192813: dataIn1 = 32'd10860
; 
32'd192814: dataIn1 = 32'd10861
; 
32'd192815: dataIn1 = 32'd10862
; 
32'd192816: dataIn1 = 32'd879
; 
32'd192817: dataIn1 = 32'd1615
; 
32'd192818: dataIn1 = 32'd10861
; 
32'd192819: dataIn1 = 32'd10862
; 
32'd192820: dataIn1 = 32'd10863
; 
32'd192821: dataIn1 = 32'd880
; 
32'd192822: dataIn1 = 32'd1615
; 
32'd192823: dataIn1 = 32'd10862
; 
32'd192824: dataIn1 = 32'd10863
; 
32'd192825: dataIn1 = 32'd10864
; 
32'd192826: dataIn1 = 32'd880
; 
32'd192827: dataIn1 = 32'd1619
; 
32'd192828: dataIn1 = 32'd10863
; 
32'd192829: dataIn1 = 32'd10864
; 
32'd192830: dataIn1 = 32'd10865
; 
32'd192831: dataIn1 = 32'd883
; 
32'd192832: dataIn1 = 32'd1619
; 
32'd192833: dataIn1 = 32'd10864
; 
32'd192834: dataIn1 = 32'd10865
; 
32'd192835: dataIn1 = 32'd10866
; 
32'd192836: dataIn1 = 32'd883
; 
32'd192837: dataIn1 = 32'd1622
; 
32'd192838: dataIn1 = 32'd10865
; 
32'd192839: dataIn1 = 32'd10866
; 
32'd192840: dataIn1 = 32'd10867
; 
32'd192841: dataIn1 = 32'd872
; 
32'd192842: dataIn1 = 32'd1622
; 
32'd192843: dataIn1 = 32'd10866
; 
32'd192844: dataIn1 = 32'd10867
; 
32'd192845: dataIn1 = 32'd10868
; 
32'd192846: dataIn1 = 32'd872
; 
32'd192847: dataIn1 = 32'd1603
; 
32'd192848: dataIn1 = 32'd10867
; 
32'd192849: dataIn1 = 32'd10868
; 
32'd192850: dataIn1 = 32'd10869
; 
32'd192851: dataIn1 = 32'd868
; 
32'd192852: dataIn1 = 32'd1603
; 
32'd192853: dataIn1 = 32'd10868
; 
32'd192854: dataIn1 = 32'd10869
; 
32'd192855: dataIn1 = 32'd10870
; 
32'd192856: dataIn1 = 32'd868
; 
32'd192857: dataIn1 = 32'd1599
; 
32'd192858: dataIn1 = 32'd10869
; 
32'd192859: dataIn1 = 32'd10870
; 
32'd192860: dataIn1 = 32'd10871
; 
32'd192861: dataIn1 = 32'd867
; 
32'd192862: dataIn1 = 32'd1599
; 
32'd192863: dataIn1 = 32'd10870
; 
32'd192864: dataIn1 = 32'd10871
; 
32'd192865: dataIn1 = 32'd10872
; 
32'd192866: dataIn1 = 32'd867
; 
32'd192867: dataIn1 = 32'd1600
; 
32'd192868: dataIn1 = 32'd10871
; 
32'd192869: dataIn1 = 32'd10872
; 
32'd192870: dataIn1 = 32'd10873
; 
32'd192871: dataIn1 = 32'd869
; 
32'd192872: dataIn1 = 32'd1600
; 
32'd192873: dataIn1 = 32'd10872
; 
32'd192874: dataIn1 = 32'd10873
; 
32'd192875: dataIn1 = 32'd10874
; 
32'd192876: dataIn1 = 32'd869
; 
32'd192877: dataIn1 = 32'd1614
; 
32'd192878: dataIn1 = 32'd10873
; 
32'd192879: dataIn1 = 32'd10874
; 
32'd192880: dataIn1 = 32'd10875
; 
32'd192881: dataIn1 = 32'd876
; 
32'd192882: dataIn1 = 32'd1614
; 
32'd192883: dataIn1 = 32'd10874
; 
32'd192884: dataIn1 = 32'd10875
; 
32'd192885: dataIn1 = 32'd10876
; 
32'd192886: dataIn1 = 32'd876
; 
32'd192887: dataIn1 = 32'd1607
; 
32'd192888: dataIn1 = 32'd10875
; 
32'd192889: dataIn1 = 32'd10876
; 
32'd192890: dataIn1 = 32'd10877
; 
32'd192891: dataIn1 = 32'd873
; 
32'd192892: dataIn1 = 32'd1607
; 
32'd192893: dataIn1 = 32'd10876
; 
32'd192894: dataIn1 = 32'd10877
; 
32'd192895: dataIn1 = 32'd10878
; 
32'd192896: dataIn1 = 32'd873
; 
32'd192897: dataIn1 = 32'd1606
; 
32'd192898: dataIn1 = 32'd10877
; 
32'd192899: dataIn1 = 32'd10878
; 
32'd192900: dataIn1 = 32'd10879
; 
32'd192901: dataIn1 = 32'd874
; 
32'd192902: dataIn1 = 32'd1606
; 
32'd192903: dataIn1 = 32'd10878
; 
32'd192904: dataIn1 = 32'd10879
; 
32'd192905: dataIn1 = 32'd10880
; 
32'd192906: dataIn1 = 32'd874
; 
32'd192907: dataIn1 = 32'd1610
; 
32'd192908: dataIn1 = 32'd10879
; 
32'd192909: dataIn1 = 32'd10880
; 
32'd192910: dataIn1 = 32'd10881
; 
32'd192911: dataIn1 = 32'd878
; 
32'd192912: dataIn1 = 32'd1610
; 
32'd192913: dataIn1 = 32'd10880
; 
32'd192914: dataIn1 = 32'd10881
; 
32'd192915: dataIn1 = 32'd10882
; 
32'd192916: dataIn1 = 32'd878
; 
32'd192917: dataIn1 = 32'd1613
; 
32'd192918: dataIn1 = 32'd10881
; 
32'd192919: dataIn1 = 32'd10882
; 
32'd192920: dataIn1 = 32'd10883
; 
32'd192921: dataIn1 = 32'd865
; 
32'd192922: dataIn1 = 32'd1613
; 
32'd192923: dataIn1 = 32'd10882
; 
32'd192924: dataIn1 = 32'd10883
; 
32'd192925: dataIn1 = 32'd10884
; 
32'd192926: dataIn1 = 32'd865
; 
32'd192927: dataIn1 = 32'd1596
; 
32'd192928: dataIn1 = 32'd10883
; 
32'd192929: dataIn1 = 32'd10884
; 
32'd192930: dataIn1 = 32'd10885
; 
32'd192931: dataIn1 = 32'd863
; 
32'd192932: dataIn1 = 32'd1596
; 
32'd192933: dataIn1 = 32'd10884
; 
32'd192934: dataIn1 = 32'd10885
; 
32'd192935: dataIn1 = 32'd10886
; 
32'd192936: dataIn1 = 32'd863
; 
32'd192937: dataIn1 = 32'd1592
; 
32'd192938: dataIn1 = 32'd10885
; 
32'd192939: dataIn1 = 32'd10886
; 
32'd192940: dataIn1 = 32'd10887
; 
32'd192941: dataIn1 = 32'd862
; 
32'd192942: dataIn1 = 32'd1592
; 
32'd192943: dataIn1 = 32'd10886
; 
32'd192944: dataIn1 = 32'd10887
; 
32'd192945: dataIn1 = 32'd10888
; 
32'd192946: dataIn1 = 32'd862
; 
32'd192947: dataIn1 = 32'd1593
; 
32'd192948: dataIn1 = 32'd10887
; 
32'd192949: dataIn1 = 32'd10888
; 
32'd192950: dataIn1 = 32'd10889
; 
32'd192951: dataIn1 = 32'd861
; 
32'd192952: dataIn1 = 32'd1593
; 
32'd192953: dataIn1 = 32'd10888
; 
32'd192954: dataIn1 = 32'd10889
; 
32'd192955: dataIn1 = 32'd10890
; 
32'd192956: dataIn1 = 32'd861
; 
32'd192957: dataIn1 = 32'd1591
; 
32'd192958: dataIn1 = 32'd10889
; 
32'd192959: dataIn1 = 32'd10890
; 
32'd192960: dataIn1 = 32'd10891
; 
32'd192961: dataIn1 = 32'd857
; 
32'd192962: dataIn1 = 32'd1591
; 
32'd192963: dataIn1 = 32'd10890
; 
32'd192964: dataIn1 = 32'd10891
; 
32'd192965: dataIn1 = 32'd10892
; 
32'd192966: dataIn1 = 32'd857
; 
32'd192967: dataIn1 = 32'd1584
; 
32'd192968: dataIn1 = 32'd10891
; 
32'd192969: dataIn1 = 32'd10892
; 
32'd192970: dataIn1 = 32'd10893
; 
32'd192971: dataIn1 = 32'd855
; 
32'd192972: dataIn1 = 32'd1584
; 
32'd192973: dataIn1 = 32'd10892
; 
32'd192974: dataIn1 = 32'd10893
; 
32'd192975: dataIn1 = 32'd10894
; 
32'd192976: dataIn1 = 32'd855
; 
32'd192977: dataIn1 = 32'd1583
; 
32'd192978: dataIn1 = 32'd10893
; 
32'd192979: dataIn1 = 32'd10894
; 
32'd192980: dataIn1 = 32'd10895
; 
32'd192981: dataIn1 = 32'd856
; 
32'd192982: dataIn1 = 32'd1583
; 
32'd192983: dataIn1 = 32'd10894
; 
32'd192984: dataIn1 = 32'd10895
; 
32'd192985: dataIn1 = 32'd10896
; 
32'd192986: dataIn1 = 32'd856
; 
32'd192987: dataIn1 = 32'd1587
; 
32'd192988: dataIn1 = 32'd10895
; 
32'd192989: dataIn1 = 32'd10896
; 
32'd192990: dataIn1 = 32'd10897
; 
32'd192991: dataIn1 = 32'd859
; 
32'd192992: dataIn1 = 32'd1587
; 
32'd192993: dataIn1 = 32'd10896
; 
32'd192994: dataIn1 = 32'd10897
; 
32'd192995: dataIn1 = 32'd10898
; 
32'd192996: dataIn1 = 32'd859
; 
32'd192997: dataIn1 = 32'd1590
; 
32'd192998: dataIn1 = 32'd10897
; 
32'd192999: dataIn1 = 32'd10898
; 
32'd193000: dataIn1 = 32'd10899
; 
32'd193001: dataIn1 = 32'd848
; 
32'd193002: dataIn1 = 32'd1590
; 
32'd193003: dataIn1 = 32'd10898
; 
32'd193004: dataIn1 = 32'd10899
; 
32'd193005: dataIn1 = 32'd10900
; 
32'd193006: dataIn1 = 32'd848
; 
32'd193007: dataIn1 = 32'd1571
; 
32'd193008: dataIn1 = 32'd10899
; 
32'd193009: dataIn1 = 32'd10900
; 
32'd193010: dataIn1 = 32'd10901
; 
32'd193011: dataIn1 = 32'd844
; 
32'd193012: dataIn1 = 32'd1571
; 
32'd193013: dataIn1 = 32'd10900
; 
32'd193014: dataIn1 = 32'd10901
; 
32'd193015: dataIn1 = 32'd10902
; 
32'd193016: dataIn1 = 32'd844
; 
32'd193017: dataIn1 = 32'd1567
; 
32'd193018: dataIn1 = 32'd10901
; 
32'd193019: dataIn1 = 32'd10902
; 
32'd193020: dataIn1 = 32'd10903
; 
32'd193021: dataIn1 = 32'd843
; 
32'd193022: dataIn1 = 32'd1567
; 
32'd193023: dataIn1 = 32'd10902
; 
32'd193024: dataIn1 = 32'd10903
; 
32'd193025: dataIn1 = 32'd10904
; 
32'd193026: dataIn1 = 32'd843
; 
32'd193027: dataIn1 = 32'd1568
; 
32'd193028: dataIn1 = 32'd10903
; 
32'd193029: dataIn1 = 32'd10904
; 
32'd193030: dataIn1 = 32'd10905
; 
32'd193031: dataIn1 = 32'd845
; 
32'd193032: dataIn1 = 32'd1568
; 
32'd193033: dataIn1 = 32'd10904
; 
32'd193034: dataIn1 = 32'd10905
; 
32'd193035: dataIn1 = 32'd10906
; 
32'd193036: dataIn1 = 32'd845
; 
32'd193037: dataIn1 = 32'd1582
; 
32'd193038: dataIn1 = 32'd10905
; 
32'd193039: dataIn1 = 32'd10906
; 
32'd193040: dataIn1 = 32'd10907
; 
32'd193041: dataIn1 = 32'd852
; 
32'd193042: dataIn1 = 32'd1582
; 
32'd193043: dataIn1 = 32'd10906
; 
32'd193044: dataIn1 = 32'd10907
; 
32'd193045: dataIn1 = 32'd10908
; 
32'd193046: dataIn1 = 32'd852
; 
32'd193047: dataIn1 = 32'd1575
; 
32'd193048: dataIn1 = 32'd10907
; 
32'd193049: dataIn1 = 32'd10908
; 
32'd193050: dataIn1 = 32'd10909
; 
32'd193051: dataIn1 = 32'd849
; 
32'd193052: dataIn1 = 32'd1575
; 
32'd193053: dataIn1 = 32'd10908
; 
32'd193054: dataIn1 = 32'd10909
; 
32'd193055: dataIn1 = 32'd10910
; 
32'd193056: dataIn1 = 32'd849
; 
32'd193057: dataIn1 = 32'd1574
; 
32'd193058: dataIn1 = 32'd10909
; 
32'd193059: dataIn1 = 32'd10910
; 
32'd193060: dataIn1 = 32'd10911
; 
32'd193061: dataIn1 = 32'd850
; 
32'd193062: dataIn1 = 32'd1574
; 
32'd193063: dataIn1 = 32'd10910
; 
32'd193064: dataIn1 = 32'd10911
; 
32'd193065: dataIn1 = 32'd10912
; 
32'd193066: dataIn1 = 32'd850
; 
32'd193067: dataIn1 = 32'd1578
; 
32'd193068: dataIn1 = 32'd10911
; 
32'd193069: dataIn1 = 32'd10912
; 
32'd193070: dataIn1 = 32'd10913
; 
32'd193071: dataIn1 = 32'd854
; 
32'd193072: dataIn1 = 32'd1578
; 
32'd193073: dataIn1 = 32'd10912
; 
32'd193074: dataIn1 = 32'd10913
; 
32'd193075: dataIn1 = 32'd10914
; 
32'd193076: dataIn1 = 32'd854
; 
32'd193077: dataIn1 = 32'd1581
; 
32'd193078: dataIn1 = 32'd10913
; 
32'd193079: dataIn1 = 32'd10914
; 
32'd193080: dataIn1 = 32'd10915
; 
32'd193081: dataIn1 = 32'd841
; 
32'd193082: dataIn1 = 32'd1581
; 
32'd193083: dataIn1 = 32'd10914
; 
32'd193084: dataIn1 = 32'd10915
; 
32'd193085: dataIn1 = 32'd10916
; 
32'd193086: dataIn1 = 32'd841
; 
32'd193087: dataIn1 = 32'd1564
; 
32'd193088: dataIn1 = 32'd10915
; 
32'd193089: dataIn1 = 32'd10916
; 
32'd193090: dataIn1 = 32'd10917
; 
32'd193091: dataIn1 = 32'd839
; 
32'd193092: dataIn1 = 32'd1564
; 
32'd193093: dataIn1 = 32'd10916
; 
32'd193094: dataIn1 = 32'd10917
; 
32'd193095: dataIn1 = 32'd10918
; 
32'd193096: dataIn1 = 32'd839
; 
32'd193097: dataIn1 = 32'd1560
; 
32'd193098: dataIn1 = 32'd10917
; 
32'd193099: dataIn1 = 32'd10918
; 
32'd193100: dataIn1 = 32'd10919
; 
32'd193101: dataIn1 = 32'd838
; 
32'd193102: dataIn1 = 32'd1560
; 
32'd193103: dataIn1 = 32'd10918
; 
32'd193104: dataIn1 = 32'd10919
; 
32'd193105: dataIn1 = 32'd10920
; 
32'd193106: dataIn1 = 32'd838
; 
32'd193107: dataIn1 = 32'd1561
; 
32'd193108: dataIn1 = 32'd10919
; 
32'd193109: dataIn1 = 32'd10920
; 
32'd193110: dataIn1 = 32'd10921
; 
32'd193111: dataIn1 = 32'd837
; 
32'd193112: dataIn1 = 32'd1561
; 
32'd193113: dataIn1 = 32'd10920
; 
32'd193114: dataIn1 = 32'd10921
; 
32'd193115: dataIn1 = 32'd10922
; 
32'd193116: dataIn1 = 32'd837
; 
32'd193117: dataIn1 = 32'd1559
; 
32'd193118: dataIn1 = 32'd10921
; 
32'd193119: dataIn1 = 32'd10922
; 
32'd193120: dataIn1 = 32'd10923
; 
32'd193121: dataIn1 = 32'd833
; 
32'd193122: dataIn1 = 32'd1559
; 
32'd193123: dataIn1 = 32'd10922
; 
32'd193124: dataIn1 = 32'd10923
; 
32'd193125: dataIn1 = 32'd10924
; 
32'd193126: dataIn1 = 32'd833
; 
32'd193127: dataIn1 = 32'd1552
; 
32'd193128: dataIn1 = 32'd10923
; 
32'd193129: dataIn1 = 32'd10924
; 
32'd193130: dataIn1 = 32'd10925
; 
32'd193131: dataIn1 = 32'd831
; 
32'd193132: dataIn1 = 32'd1552
; 
32'd193133: dataIn1 = 32'd10924
; 
32'd193134: dataIn1 = 32'd10925
; 
32'd193135: dataIn1 = 32'd10926
; 
32'd193136: dataIn1 = 32'd831
; 
32'd193137: dataIn1 = 32'd1551
; 
32'd193138: dataIn1 = 32'd10925
; 
32'd193139: dataIn1 = 32'd10926
; 
32'd193140: dataIn1 = 32'd10927
; 
32'd193141: dataIn1 = 32'd832
; 
32'd193142: dataIn1 = 32'd1551
; 
32'd193143: dataIn1 = 32'd10926
; 
32'd193144: dataIn1 = 32'd10927
; 
32'd193145: dataIn1 = 32'd10928
; 
32'd193146: dataIn1 = 32'd832
; 
32'd193147: dataIn1 = 32'd1555
; 
32'd193148: dataIn1 = 32'd10927
; 
32'd193149: dataIn1 = 32'd10928
; 
32'd193150: dataIn1 = 32'd10929
; 
32'd193151: dataIn1 = 32'd835
; 
32'd193152: dataIn1 = 32'd1555
; 
32'd193153: dataIn1 = 32'd10928
; 
32'd193154: dataIn1 = 32'd10929
; 
32'd193155: dataIn1 = 32'd10930
; 
32'd193156: dataIn1 = 32'd835
; 
32'd193157: dataIn1 = 32'd1558
; 
32'd193158: dataIn1 = 32'd10929
; 
32'd193159: dataIn1 = 32'd10930
; 
32'd193160: dataIn1 = 32'd10931
; 
32'd193161: dataIn1 = 32'd824
; 
32'd193162: dataIn1 = 32'd1558
; 
32'd193163: dataIn1 = 32'd10930
; 
32'd193164: dataIn1 = 32'd10931
; 
32'd193165: dataIn1 = 32'd10932
; 
32'd193166: dataIn1 = 32'd824
; 
32'd193167: dataIn1 = 32'd1539
; 
32'd193168: dataIn1 = 32'd10931
; 
32'd193169: dataIn1 = 32'd10932
; 
32'd193170: dataIn1 = 32'd10933
; 
32'd193171: dataIn1 = 32'd820
; 
32'd193172: dataIn1 = 32'd1539
; 
32'd193173: dataIn1 = 32'd10932
; 
32'd193174: dataIn1 = 32'd10933
; 
32'd193175: dataIn1 = 32'd10934
; 
32'd193176: dataIn1 = 32'd820
; 
32'd193177: dataIn1 = 32'd1535
; 
32'd193178: dataIn1 = 32'd10933
; 
32'd193179: dataIn1 = 32'd10934
; 
32'd193180: dataIn1 = 32'd10935
; 
32'd193181: dataIn1 = 32'd819
; 
32'd193182: dataIn1 = 32'd1535
; 
32'd193183: dataIn1 = 32'd10934
; 
32'd193184: dataIn1 = 32'd10935
; 
32'd193185: dataIn1 = 32'd10936
; 
32'd193186: dataIn1 = 32'd819
; 
32'd193187: dataIn1 = 32'd1536
; 
32'd193188: dataIn1 = 32'd10935
; 
32'd193189: dataIn1 = 32'd10936
; 
32'd193190: dataIn1 = 32'd10937
; 
32'd193191: dataIn1 = 32'd821
; 
32'd193192: dataIn1 = 32'd1536
; 
32'd193193: dataIn1 = 32'd10936
; 
32'd193194: dataIn1 = 32'd10937
; 
32'd193195: dataIn1 = 32'd10938
; 
32'd193196: dataIn1 = 32'd821
; 
32'd193197: dataIn1 = 32'd1550
; 
32'd193198: dataIn1 = 32'd10937
; 
32'd193199: dataIn1 = 32'd10938
; 
32'd193200: dataIn1 = 32'd10939
; 
32'd193201: dataIn1 = 32'd828
; 
32'd193202: dataIn1 = 32'd1550
; 
32'd193203: dataIn1 = 32'd10938
; 
32'd193204: dataIn1 = 32'd10939
; 
32'd193205: dataIn1 = 32'd10940
; 
32'd193206: dataIn1 = 32'd828
; 
32'd193207: dataIn1 = 32'd1543
; 
32'd193208: dataIn1 = 32'd10939
; 
32'd193209: dataIn1 = 32'd10940
; 
32'd193210: dataIn1 = 32'd10941
; 
32'd193211: dataIn1 = 32'd825
; 
32'd193212: dataIn1 = 32'd1543
; 
32'd193213: dataIn1 = 32'd10940
; 
32'd193214: dataIn1 = 32'd10941
; 
32'd193215: dataIn1 = 32'd10942
; 
32'd193216: dataIn1 = 32'd825
; 
32'd193217: dataIn1 = 32'd1542
; 
32'd193218: dataIn1 = 32'd10941
; 
32'd193219: dataIn1 = 32'd10942
; 
32'd193220: dataIn1 = 32'd10943
; 
32'd193221: dataIn1 = 32'd826
; 
32'd193222: dataIn1 = 32'd1542
; 
32'd193223: dataIn1 = 32'd10942
; 
32'd193224: dataIn1 = 32'd10943
; 
32'd193225: dataIn1 = 32'd10944
; 
32'd193226: dataIn1 = 32'd826
; 
32'd193227: dataIn1 = 32'd1546
; 
32'd193228: dataIn1 = 32'd10943
; 
32'd193229: dataIn1 = 32'd10944
; 
32'd193230: dataIn1 = 32'd10945
; 
32'd193231: dataIn1 = 32'd830
; 
32'd193232: dataIn1 = 32'd1546
; 
32'd193233: dataIn1 = 32'd10944
; 
32'd193234: dataIn1 = 32'd10945
; 
32'd193235: dataIn1 = 32'd10946
; 
32'd193236: dataIn1 = 32'd830
; 
32'd193237: dataIn1 = 32'd1549
; 
32'd193238: dataIn1 = 32'd10945
; 
32'd193239: dataIn1 = 32'd10946
; 
32'd193240: dataIn1 = 32'd10947
; 
32'd193241: dataIn1 = 32'd817
; 
32'd193242: dataIn1 = 32'd1549
; 
32'd193243: dataIn1 = 32'd10946
; 
32'd193244: dataIn1 = 32'd10947
; 
32'd193245: dataIn1 = 32'd10948
; 
32'd193246: dataIn1 = 32'd817
; 
32'd193247: dataIn1 = 32'd1532
; 
32'd193248: dataIn1 = 32'd10947
; 
32'd193249: dataIn1 = 32'd10948
; 
32'd193250: dataIn1 = 32'd10949
; 
32'd193251: dataIn1 = 32'd815
; 
32'd193252: dataIn1 = 32'd1532
; 
32'd193253: dataIn1 = 32'd10948
; 
32'd193254: dataIn1 = 32'd10949
; 
32'd193255: dataIn1 = 32'd10950
; 
32'd193256: dataIn1 = 32'd815
; 
32'd193257: dataIn1 = 32'd1528
; 
32'd193258: dataIn1 = 32'd10949
; 
32'd193259: dataIn1 = 32'd10950
; 
32'd193260: dataIn1 = 32'd10951
; 
32'd193261: dataIn1 = 32'd814
; 
32'd193262: dataIn1 = 32'd1528
; 
32'd193263: dataIn1 = 32'd10950
; 
32'd193264: dataIn1 = 32'd10951
; 
32'd193265: dataIn1 = 32'd10952
; 
32'd193266: dataIn1 = 32'd814
; 
32'd193267: dataIn1 = 32'd1529
; 
32'd193268: dataIn1 = 32'd10951
; 
32'd193269: dataIn1 = 32'd10952
; 
32'd193270: dataIn1 = 32'd10953
; 
32'd193271: dataIn1 = 32'd813
; 
32'd193272: dataIn1 = 32'd1529
; 
32'd193273: dataIn1 = 32'd10952
; 
32'd193274: dataIn1 = 32'd10953
; 
32'd193275: dataIn1 = 32'd10954
; 
32'd193276: dataIn1 = 32'd813
; 
32'd193277: dataIn1 = 32'd1527
; 
32'd193278: dataIn1 = 32'd10953
; 
32'd193279: dataIn1 = 32'd10954
; 
32'd193280: dataIn1 = 32'd10955
; 
32'd193281: dataIn1 = 32'd809
; 
32'd193282: dataIn1 = 32'd1527
; 
32'd193283: dataIn1 = 32'd10954
; 
32'd193284: dataIn1 = 32'd10955
; 
32'd193285: dataIn1 = 32'd10956
; 
32'd193286: dataIn1 = 32'd809
; 
32'd193287: dataIn1 = 32'd1520
; 
32'd193288: dataIn1 = 32'd10955
; 
32'd193289: dataIn1 = 32'd10956
; 
32'd193290: dataIn1 = 32'd10957
; 
32'd193291: dataIn1 = 32'd807
; 
32'd193292: dataIn1 = 32'd1520
; 
32'd193293: dataIn1 = 32'd10956
; 
32'd193294: dataIn1 = 32'd10957
; 
32'd193295: dataIn1 = 32'd10958
; 
32'd193296: dataIn1 = 32'd807
; 
32'd193297: dataIn1 = 32'd1519
; 
32'd193298: dataIn1 = 32'd10957
; 
32'd193299: dataIn1 = 32'd10958
; 
32'd193300: dataIn1 = 32'd10959
; 
32'd193301: dataIn1 = 32'd808
; 
32'd193302: dataIn1 = 32'd1519
; 
32'd193303: dataIn1 = 32'd10958
; 
32'd193304: dataIn1 = 32'd10959
; 
32'd193305: dataIn1 = 32'd10960
; 
32'd193306: dataIn1 = 32'd808
; 
32'd193307: dataIn1 = 32'd1523
; 
32'd193308: dataIn1 = 32'd10959
; 
32'd193309: dataIn1 = 32'd10960
; 
32'd193310: dataIn1 = 32'd10961
; 
32'd193311: dataIn1 = 32'd811
; 
32'd193312: dataIn1 = 32'd1523
; 
32'd193313: dataIn1 = 32'd10960
; 
32'd193314: dataIn1 = 32'd10961
; 
32'd193315: dataIn1 = 32'd10962
; 
32'd193316: dataIn1 = 32'd811
; 
32'd193317: dataIn1 = 32'd1526
; 
32'd193318: dataIn1 = 32'd10961
; 
32'd193319: dataIn1 = 32'd10962
; 
32'd193320: dataIn1 = 32'd10963
; 
32'd193321: dataIn1 = 32'd797
; 
32'd193322: dataIn1 = 32'd1526
; 
32'd193323: dataIn1 = 32'd10962
; 
32'd193324: dataIn1 = 32'd10963
; 
32'd193325: dataIn1 = 32'd10964
; 
32'd193326: dataIn1 = 32'd797
; 
32'd193327: dataIn1 = 32'd1503
; 
32'd193328: dataIn1 = 32'd10963
; 
32'd193329: dataIn1 = 32'd10964
; 
32'd193330: dataIn1 = 32'd10965
; 
32'd193331: dataIn1 = 32'd793
; 
32'd193332: dataIn1 = 32'd1503
; 
32'd193333: dataIn1 = 32'd10964
; 
32'd193334: dataIn1 = 32'd10965
; 
32'd193335: dataIn1 = 32'd10966
; 
32'd193336: dataIn1 = 32'd793
; 
32'd193337: dataIn1 = 32'd1499
; 
32'd193338: dataIn1 = 32'd10965
; 
32'd193339: dataIn1 = 32'd10966
; 
32'd193340: dataIn1 = 32'd10967
; 
32'd193341: dataIn1 = 32'd792
; 
32'd193342: dataIn1 = 32'd1499
; 
32'd193343: dataIn1 = 32'd10966
; 
32'd193344: dataIn1 = 32'd10967
; 
32'd193345: dataIn1 = 32'd10968
; 
32'd193346: dataIn1 = 32'd792
; 
32'd193347: dataIn1 = 32'd1500
; 
32'd193348: dataIn1 = 32'd10967
; 
32'd193349: dataIn1 = 32'd10968
; 
32'd193350: dataIn1 = 32'd10969
; 
32'd193351: dataIn1 = 32'd794
; 
32'd193352: dataIn1 = 32'd1500
; 
32'd193353: dataIn1 = 32'd10968
; 
32'd193354: dataIn1 = 32'd10969
; 
32'd193355: dataIn1 = 32'd10970
; 
32'd193356: dataIn1 = 32'd794
; 
32'd193357: dataIn1 = 32'd1515
; 
32'd193358: dataIn1 = 32'd1516
; 
32'd193359: dataIn1 = 32'd10969
; 
32'd193360: dataIn1 = 32'd10970
; 
32'd193361: dataIn1 = 32'd10971
; 
32'd193362: dataIn1 = 32'd1516
; 
32'd193363: dataIn1 = 32'd10970
; 
32'd193364: dataIn1 = 32'd10971
; 
32'd193365: dataIn1 = 32'd10972
; 
32'd193366: dataIn1 = 32'd1516
; 
32'd193367: dataIn1 = 32'd10971
; 
32'd193368: dataIn1 = 32'd10972
; 
32'd193369: dataIn1 = 32'd10973
; 
32'd193370: dataIn1 = 32'd414
; 
32'd193371: dataIn1 = 32'd1516
; 
32'd193372: dataIn1 = 32'd1517
; 
32'd193373: dataIn1 = 32'd10972
; 
32'd193374: dataIn1 = 32'd10973
; 
32'd193375: dataIn1 = 32'd10974
; 
32'd193376: dataIn1 = 32'd414
; 
32'd193377: dataIn1 = 32'd1514
; 
32'd193378: dataIn1 = 32'd10973
; 
32'd193379: dataIn1 = 32'd10974
; 
32'd193380: dataIn1 = 32'd10975
; 
32'd193381: dataIn1 = 32'd1514
; 
32'd193382: dataIn1 = 32'd10974
; 
32'd193383: dataIn1 = 32'd10975
; 
32'd193384: dataIn1 = 32'd10976
; 
32'd193385: dataIn1 = 32'd1514
; 
32'd193386: dataIn1 = 32'd1518
; 
32'd193387: dataIn1 = 32'd2760
; 
32'd193388: dataIn1 = 32'd10975
; 
32'd193389: dataIn1 = 32'd10976
; 
32'd193390: dataIn1 = 32'd10977
; 
32'd193391: dataIn1 = 32'd1518
; 
32'd193392: dataIn1 = 32'd10976
; 
32'd193393: dataIn1 = 32'd10977
; 
32'd193394: dataIn1 = 32'd10978
; 
32'd193395: dataIn1 = 32'd585
; 
32'd193396: dataIn1 = 32'd1518
; 
32'd193397: dataIn1 = 32'd10977
; 
32'd193398: dataIn1 = 32'd10978
; 
32'd193399: dataIn1 = 32'd10979
; 
32'd193400: dataIn1 = 32'd585
; 
32'd193401: dataIn1 = 32'd1300
; 
32'd193402: dataIn1 = 32'd10978
; 
32'd193403: dataIn1 = 32'd10979
; 
32'd193404: dataIn1 = 32'd10980
; 
32'd193405: dataIn1 = 32'd1300
; 
32'd193406: dataIn1 = 32'd10979
; 
32'd193407: dataIn1 = 32'd10980
; 
32'd193408: dataIn1 = 32'd10981
; 
32'd193409: dataIn1 = 32'd584
; 
32'd193410: dataIn1 = 32'd1300
; 
32'd193411: dataIn1 = 32'd10980
; 
32'd193412: dataIn1 = 32'd10981
; 
32'd193413: dataIn1 = 32'd10982
; 
32'd193414: dataIn1 = 32'd584
; 
32'd193415: dataIn1 = 32'd10981
; 
32'd193416: dataIn1 = 32'd10982
; 
32'd193417: dataIn1 = 32'd10983
; 
32'd193418: dataIn1 = 32'd584
; 
32'd193419: dataIn1 = 32'd2484
; 
32'd193420: dataIn1 = 32'd10982
; 
32'd193421: dataIn1 = 32'd10983
; 
32'd193422: dataIn1 = 32'd10984
; 
32'd193423: dataIn1 = 32'd2484
; 
32'd193424: dataIn1 = 32'd10983
; 
32'd193425: dataIn1 = 32'd10984
; 
32'd193426: dataIn1 = 32'd10985
; 
32'd193427: dataIn1 = 32'd583
; 
32'd193428: dataIn1 = 32'd2484
; 
32'd193429: dataIn1 = 32'd2757
; 
32'd193430: dataIn1 = 32'd10984
; 
32'd193431: dataIn1 = 32'd10985
; 
32'd193432: dataIn1 = 32'd10986
; 
32'd193433: dataIn1 = 32'd583
; 
32'd193434: dataIn1 = 32'd10985
; 
32'd193435: dataIn1 = 32'd10986
; 
32'd193436: dataIn1 = 32'd10987
; 
32'd193437: dataIn1 = 32'd583
; 
32'd193438: dataIn1 = 32'd1299
; 
32'd193439: dataIn1 = 32'd10986
; 
32'd193440: dataIn1 = 32'd10987
; 
32'd193441: dataIn1 = 32'd10988
; 
32'd193442: dataIn1 = 32'd1299
; 
32'd193443: dataIn1 = 32'd10987
; 
32'd193444: dataIn1 = 32'd10988
; 
32'd193445: dataIn1 = 32'd10989
; 
32'd193446: dataIn1 = 32'd1299
; 
32'd193447: dataIn1 = 32'd3053
; 
32'd193448: dataIn1 = 32'd3054
; 
32'd193449: dataIn1 = 32'd10988
; 
32'd193450: dataIn1 = 32'd10989
; 
32'd193451: dataIn1 = 32'd10990
; 
32'd193452: dataIn1 = 32'd2763
; 
32'd193453: dataIn1 = 32'd3053
; 
32'd193454: dataIn1 = 32'd10989
; 
32'd193455: dataIn1 = 32'd10990
; 
32'd193456: dataIn1 = 32'd10991
; 
32'd193457: dataIn1 = 32'd2762
; 
32'd193458: dataIn1 = 32'd2763
; 
32'd193459: dataIn1 = 32'd10990
; 
32'd193460: dataIn1 = 32'd10991
; 
32'd193461: dataIn1 = 32'd10992
; 
32'd193462: dataIn1 = 32'd2762
; 
32'd193463: dataIn1 = 32'd3045
; 
32'd193464: dataIn1 = 32'd10991
; 
32'd193465: dataIn1 = 32'd10992
; 
32'd193466: dataIn1 = 32'd10993
; 
32'd193467: dataIn1 = 32'd3045
; 
32'd193468: dataIn1 = 32'd3046
; 
32'd193469: dataIn1 = 32'd10992
; 
32'd193470: dataIn1 = 32'd10993
; 
32'd193471: dataIn1 = 32'd10994
; 
32'd193472: dataIn1 = 32'd2778
; 
32'd193473: dataIn1 = 32'd3046
; 
32'd193474: dataIn1 = 32'd10993
; 
32'd193475: dataIn1 = 32'd10994
; 
32'd193476: dataIn1 = 32'd10995
; 
32'd193477: dataIn1 = 32'd2777
; 
32'd193478: dataIn1 = 32'd2778
; 
32'd193479: dataIn1 = 32'd10994
; 
32'd193480: dataIn1 = 32'd10995
; 
32'd193481: dataIn1 = 32'd10996
; 
32'd193482: dataIn1 = 32'd2777
; 
32'd193483: dataIn1 = 32'd3059
; 
32'd193484: dataIn1 = 32'd10995
; 
32'd193485: dataIn1 = 32'd10996
; 
32'd193486: dataIn1 = 32'd10997
; 
32'd193487: dataIn1 = 32'd3058
; 
32'd193488: dataIn1 = 32'd3059
; 
32'd193489: dataIn1 = 32'd10996
; 
32'd193490: dataIn1 = 32'd10997
; 
32'd193491: dataIn1 = 32'd10998
; 
32'd193492: dataIn1 = 32'd2772
; 
32'd193493: dataIn1 = 32'd3058
; 
32'd193494: dataIn1 = 32'd10997
; 
32'd193495: dataIn1 = 32'd10998
; 
32'd193496: dataIn1 = 32'd10999
; 
32'd193497: dataIn1 = 32'd2772
; 
32'd193498: dataIn1 = 32'd2774
; 
32'd193499: dataIn1 = 32'd10998
; 
32'd193500: dataIn1 = 32'd10999
; 
32'd193501: dataIn1 = 32'd11000
; 
32'd193502: dataIn1 = 32'd2774
; 
32'd193503: dataIn1 = 32'd3068
; 
32'd193504: dataIn1 = 32'd10999
; 
32'd193505: dataIn1 = 32'd11000
; 
32'd193506: dataIn1 = 32'd11001
; 
32'd193507: dataIn1 = 32'd3067
; 
32'd193508: dataIn1 = 32'd3068
; 
32'd193509: dataIn1 = 32'd11000
; 
32'd193510: dataIn1 = 32'd11001
; 
32'd193511: dataIn1 = 32'd11002
; 
32'd193512: dataIn1 = 32'd2784
; 
32'd193513: dataIn1 = 32'd3067
; 
32'd193514: dataIn1 = 32'd11001
; 
32'd193515: dataIn1 = 32'd11002
; 
32'd193516: dataIn1 = 32'd11003
; 
32'd193517: dataIn1 = 32'd2783
; 
32'd193518: dataIn1 = 32'd2784
; 
32'd193519: dataIn1 = 32'd11002
; 
32'd193520: dataIn1 = 32'd11003
; 
32'd193521: dataIn1 = 32'd11004
; 
32'd193522: dataIn1 = 32'd2783
; 
32'd193523: dataIn1 = 32'd3074
; 
32'd193524: dataIn1 = 32'd11003
; 
32'd193525: dataIn1 = 32'd11004
; 
32'd193526: dataIn1 = 32'd11005
; 
32'd193527: dataIn1 = 32'd3074
; 
32'd193528: dataIn1 = 32'd3075
; 
32'd193529: dataIn1 = 32'd11004
; 
32'd193530: dataIn1 = 32'd11005
; 
32'd193531: dataIn1 = 32'd11006
; 
32'd193532: dataIn1 = 32'd2789
; 
32'd193533: dataIn1 = 32'd3075
; 
32'd193534: dataIn1 = 32'd11005
; 
32'd193535: dataIn1 = 32'd11006
; 
32'd193536: dataIn1 = 32'd11007
; 
32'd193537: dataIn1 = 32'd2787
; 
32'd193538: dataIn1 = 32'd2789
; 
32'd193539: dataIn1 = 32'd11006
; 
32'd193540: dataIn1 = 32'd11007
; 
32'd193541: dataIn1 = 32'd11008
; 
32'd193542: dataIn1 = 32'd2787
; 
32'd193543: dataIn1 = 32'd3079
; 
32'd193544: dataIn1 = 32'd11007
; 
32'd193545: dataIn1 = 32'd11008
; 
32'd193546: dataIn1 = 32'd11009
; 
32'd193547: dataIn1 = 32'd3079
; 
32'd193548: dataIn1 = 32'd3080
; 
32'd193549: dataIn1 = 32'd11008
; 
32'd193550: dataIn1 = 32'd11009
; 
32'd193551: dataIn1 = 32'd11010
; 
32'd193552: dataIn1 = 32'd2809
; 
32'd193553: dataIn1 = 32'd3080
; 
32'd193554: dataIn1 = 32'd11009
; 
32'd193555: dataIn1 = 32'd11010
; 
32'd193556: dataIn1 = 32'd11011
; 
32'd193557: dataIn1 = 32'd2808
; 
32'd193558: dataIn1 = 32'd2809
; 
32'd193559: dataIn1 = 32'd11010
; 
32'd193560: dataIn1 = 32'd11011
; 
32'd193561: dataIn1 = 32'd11012
; 
32'd193562: dataIn1 = 32'd2808
; 
32'd193563: dataIn1 = 32'd3108
; 
32'd193564: dataIn1 = 32'd11011
; 
32'd193565: dataIn1 = 32'd11012
; 
32'd193566: dataIn1 = 32'd11013
; 
32'd193567: dataIn1 = 32'd3108
; 
32'd193568: dataIn1 = 32'd3109
; 
32'd193569: dataIn1 = 32'd11012
; 
32'd193570: dataIn1 = 32'd11013
; 
32'd193571: dataIn1 = 32'd11014
; 
32'd193572: dataIn1 = 32'd2798
; 
32'd193573: dataIn1 = 32'd3109
; 
32'd193574: dataIn1 = 32'd11013
; 
32'd193575: dataIn1 = 32'd11014
; 
32'd193576: dataIn1 = 32'd11015
; 
32'd193577: dataIn1 = 32'd2797
; 
32'd193578: dataIn1 = 32'd2798
; 
32'd193579: dataIn1 = 32'd11014
; 
32'd193580: dataIn1 = 32'd11015
; 
32'd193581: dataIn1 = 32'd11016
; 
32'd193582: dataIn1 = 32'd2797
; 
32'd193583: dataIn1 = 32'd3101
; 
32'd193584: dataIn1 = 32'd11015
; 
32'd193585: dataIn1 = 32'd11016
; 
32'd193586: dataIn1 = 32'd11017
; 
32'd193587: dataIn1 = 32'd3100
; 
32'd193588: dataIn1 = 32'd3101
; 
32'd193589: dataIn1 = 32'd11016
; 
32'd193590: dataIn1 = 32'd11017
; 
32'd193591: dataIn1 = 32'd11018
; 
32'd193592: dataIn1 = 32'd2802
; 
32'd193593: dataIn1 = 32'd3100
; 
32'd193594: dataIn1 = 32'd11017
; 
32'd193595: dataIn1 = 32'd11018
; 
32'd193596: dataIn1 = 32'd11019
; 
32'd193597: dataIn1 = 32'd2802
; 
32'd193598: dataIn1 = 32'd2804
; 
32'd193599: dataIn1 = 32'd11018
; 
32'd193600: dataIn1 = 32'd11019
; 
32'd193601: dataIn1 = 32'd11020
; 
32'd193602: dataIn1 = 32'd2804
; 
32'd193603: dataIn1 = 32'd3096
; 
32'd193604: dataIn1 = 32'd11019
; 
32'd193605: dataIn1 = 32'd11020
; 
32'd193606: dataIn1 = 32'd11021
; 
32'd193607: dataIn1 = 32'd3095
; 
32'd193608: dataIn1 = 32'd3096
; 
32'd193609: dataIn1 = 32'd11020
; 
32'd193610: dataIn1 = 32'd11021
; 
32'd193611: dataIn1 = 32'd11022
; 
32'd193612: dataIn1 = 32'd2794
; 
32'd193613: dataIn1 = 32'd3095
; 
32'd193614: dataIn1 = 32'd11021
; 
32'd193615: dataIn1 = 32'd11022
; 
32'd193616: dataIn1 = 32'd11023
; 
32'd193617: dataIn1 = 32'd2793
; 
32'd193618: dataIn1 = 32'd2794
; 
32'd193619: dataIn1 = 32'd11022
; 
32'd193620: dataIn1 = 32'd11023
; 
32'd193621: dataIn1 = 32'd11024
; 
32'd193622: dataIn1 = 32'd2793
; 
32'd193623: dataIn1 = 32'd3087
; 
32'd193624: dataIn1 = 32'd11023
; 
32'd193625: dataIn1 = 32'd11024
; 
32'd193626: dataIn1 = 32'd11025
; 
32'd193627: dataIn1 = 32'd3087
; 
32'd193628: dataIn1 = 32'd3088
; 
32'd193629: dataIn1 = 32'd11024
; 
32'd193630: dataIn1 = 32'd11025
; 
32'd193631: dataIn1 = 32'd11026
; 
32'd193632: dataIn1 = 32'd2818
; 
32'd193633: dataIn1 = 32'd3088
; 
32'd193634: dataIn1 = 32'd11025
; 
32'd193635: dataIn1 = 32'd11026
; 
32'd193636: dataIn1 = 32'd11027
; 
32'd193637: dataIn1 = 32'd2817
; 
32'd193638: dataIn1 = 32'd2818
; 
32'd193639: dataIn1 = 32'd11026
; 
32'd193640: dataIn1 = 32'd11027
; 
32'd193641: dataIn1 = 32'd11028
; 
32'd193642: dataIn1 = 32'd2817
; 
32'd193643: dataIn1 = 32'd3115
; 
32'd193644: dataIn1 = 32'd11027
; 
32'd193645: dataIn1 = 32'd11028
; 
32'd193646: dataIn1 = 32'd11029
; 
32'd193647: dataIn1 = 32'd3114
; 
32'd193648: dataIn1 = 32'd3115
; 
32'd193649: dataIn1 = 32'd11028
; 
32'd193650: dataIn1 = 32'd11029
; 
32'd193651: dataIn1 = 32'd11030
; 
32'd193652: dataIn1 = 32'd2812
; 
32'd193653: dataIn1 = 32'd3114
; 
32'd193654: dataIn1 = 32'd11029
; 
32'd193655: dataIn1 = 32'd11030
; 
32'd193656: dataIn1 = 32'd11031
; 
32'd193657: dataIn1 = 32'd2812
; 
32'd193658: dataIn1 = 32'd2814
; 
32'd193659: dataIn1 = 32'd11030
; 
32'd193660: dataIn1 = 32'd11031
; 
32'd193661: dataIn1 = 32'd11032
; 
32'd193662: dataIn1 = 32'd2814
; 
32'd193663: dataIn1 = 32'd3124
; 
32'd193664: dataIn1 = 32'd11031
; 
32'd193665: dataIn1 = 32'd11032
; 
32'd193666: dataIn1 = 32'd11033
; 
32'd193667: dataIn1 = 32'd3123
; 
32'd193668: dataIn1 = 32'd3124
; 
32'd193669: dataIn1 = 32'd11032
; 
32'd193670: dataIn1 = 32'd11033
; 
32'd193671: dataIn1 = 32'd11034
; 
32'd193672: dataIn1 = 32'd2824
; 
32'd193673: dataIn1 = 32'd3123
; 
32'd193674: dataIn1 = 32'd11033
; 
32'd193675: dataIn1 = 32'd11034
; 
32'd193676: dataIn1 = 32'd11035
; 
32'd193677: dataIn1 = 32'd2823
; 
32'd193678: dataIn1 = 32'd2824
; 
32'd193679: dataIn1 = 32'd11034
; 
32'd193680: dataIn1 = 32'd11035
; 
32'd193681: dataIn1 = 32'd11036
; 
32'd193682: dataIn1 = 32'd2823
; 
32'd193683: dataIn1 = 32'd3130
; 
32'd193684: dataIn1 = 32'd11035
; 
32'd193685: dataIn1 = 32'd11036
; 
32'd193686: dataIn1 = 32'd11037
; 
32'd193687: dataIn1 = 32'd3130
; 
32'd193688: dataIn1 = 32'd3131
; 
32'd193689: dataIn1 = 32'd11036
; 
32'd193690: dataIn1 = 32'd11037
; 
32'd193691: dataIn1 = 32'd11038
; 
32'd193692: dataIn1 = 32'd2829
; 
32'd193693: dataIn1 = 32'd3131
; 
32'd193694: dataIn1 = 32'd11037
; 
32'd193695: dataIn1 = 32'd11038
; 
32'd193696: dataIn1 = 32'd11039
; 
32'd193697: dataIn1 = 32'd2827
; 
32'd193698: dataIn1 = 32'd2829
; 
32'd193699: dataIn1 = 32'd11038
; 
32'd193700: dataIn1 = 32'd11039
; 
32'd193701: dataIn1 = 32'd11040
; 
32'd193702: dataIn1 = 32'd2827
; 
32'd193703: dataIn1 = 32'd3135
; 
32'd193704: dataIn1 = 32'd11039
; 
32'd193705: dataIn1 = 32'd11040
; 
32'd193706: dataIn1 = 32'd11041
; 
32'd193707: dataIn1 = 32'd3135
; 
32'd193708: dataIn1 = 32'd3136
; 
32'd193709: dataIn1 = 32'd11040
; 
32'd193710: dataIn1 = 32'd11041
; 
32'd193711: dataIn1 = 32'd11042
; 
32'd193712: dataIn1 = 32'd2849
; 
32'd193713: dataIn1 = 32'd3136
; 
32'd193714: dataIn1 = 32'd11041
; 
32'd193715: dataIn1 = 32'd11042
; 
32'd193716: dataIn1 = 32'd11043
; 
32'd193717: dataIn1 = 32'd2848
; 
32'd193718: dataIn1 = 32'd2849
; 
32'd193719: dataIn1 = 32'd11042
; 
32'd193720: dataIn1 = 32'd11043
; 
32'd193721: dataIn1 = 32'd11044
; 
32'd193722: dataIn1 = 32'd2848
; 
32'd193723: dataIn1 = 32'd3164
; 
32'd193724: dataIn1 = 32'd11043
; 
32'd193725: dataIn1 = 32'd11044
; 
32'd193726: dataIn1 = 32'd11045
; 
32'd193727: dataIn1 = 32'd3164
; 
32'd193728: dataIn1 = 32'd3165
; 
32'd193729: dataIn1 = 32'd11044
; 
32'd193730: dataIn1 = 32'd11045
; 
32'd193731: dataIn1 = 32'd11046
; 
32'd193732: dataIn1 = 32'd2838
; 
32'd193733: dataIn1 = 32'd3165
; 
32'd193734: dataIn1 = 32'd11045
; 
32'd193735: dataIn1 = 32'd11046
; 
32'd193736: dataIn1 = 32'd11047
; 
32'd193737: dataIn1 = 32'd2837
; 
32'd193738: dataIn1 = 32'd2838
; 
32'd193739: dataIn1 = 32'd11046
; 
32'd193740: dataIn1 = 32'd11047
; 
32'd193741: dataIn1 = 32'd11048
; 
32'd193742: dataIn1 = 32'd2837
; 
32'd193743: dataIn1 = 32'd3157
; 
32'd193744: dataIn1 = 32'd11047
; 
32'd193745: dataIn1 = 32'd11048
; 
32'd193746: dataIn1 = 32'd11049
; 
32'd193747: dataIn1 = 32'd3156
; 
32'd193748: dataIn1 = 32'd3157
; 
32'd193749: dataIn1 = 32'd11048
; 
32'd193750: dataIn1 = 32'd11049
; 
32'd193751: dataIn1 = 32'd11050
; 
32'd193752: dataIn1 = 32'd2842
; 
32'd193753: dataIn1 = 32'd3156
; 
32'd193754: dataIn1 = 32'd11049
; 
32'd193755: dataIn1 = 32'd11050
; 
32'd193756: dataIn1 = 32'd11051
; 
32'd193757: dataIn1 = 32'd2842
; 
32'd193758: dataIn1 = 32'd2844
; 
32'd193759: dataIn1 = 32'd11050
; 
32'd193760: dataIn1 = 32'd11051
; 
32'd193761: dataIn1 = 32'd11052
; 
32'd193762: dataIn1 = 32'd2844
; 
32'd193763: dataIn1 = 32'd3152
; 
32'd193764: dataIn1 = 32'd11051
; 
32'd193765: dataIn1 = 32'd11052
; 
32'd193766: dataIn1 = 32'd11053
; 
32'd193767: dataIn1 = 32'd3151
; 
32'd193768: dataIn1 = 32'd3152
; 
32'd193769: dataIn1 = 32'd11052
; 
32'd193770: dataIn1 = 32'd11053
; 
32'd193771: dataIn1 = 32'd11054
; 
32'd193772: dataIn1 = 32'd2834
; 
32'd193773: dataIn1 = 32'd3151
; 
32'd193774: dataIn1 = 32'd11053
; 
32'd193775: dataIn1 = 32'd11054
; 
32'd193776: dataIn1 = 32'd11055
; 
32'd193777: dataIn1 = 32'd2833
; 
32'd193778: dataIn1 = 32'd2834
; 
32'd193779: dataIn1 = 32'd11054
; 
32'd193780: dataIn1 = 32'd11055
; 
32'd193781: dataIn1 = 32'd11056
; 
32'd193782: dataIn1 = 32'd2833
; 
32'd193783: dataIn1 = 32'd3143
; 
32'd193784: dataIn1 = 32'd11055
; 
32'd193785: dataIn1 = 32'd11056
; 
32'd193786: dataIn1 = 32'd11057
; 
32'd193787: dataIn1 = 32'd3143
; 
32'd193788: dataIn1 = 32'd3144
; 
32'd193789: dataIn1 = 32'd11056
; 
32'd193790: dataIn1 = 32'd11057
; 
32'd193791: dataIn1 = 32'd11058
; 
32'd193792: dataIn1 = 32'd2858
; 
32'd193793: dataIn1 = 32'd3144
; 
32'd193794: dataIn1 = 32'd11057
; 
32'd193795: dataIn1 = 32'd11058
; 
32'd193796: dataIn1 = 32'd11059
; 
32'd193797: dataIn1 = 32'd2857
; 
32'd193798: dataIn1 = 32'd2858
; 
32'd193799: dataIn1 = 32'd11058
; 
32'd193800: dataIn1 = 32'd11059
; 
32'd193801: dataIn1 = 32'd11060
; 
32'd193802: dataIn1 = 32'd2857
; 
32'd193803: dataIn1 = 32'd3171
; 
32'd193804: dataIn1 = 32'd11059
; 
32'd193805: dataIn1 = 32'd11060
; 
32'd193806: dataIn1 = 32'd11061
; 
32'd193807: dataIn1 = 32'd3170
; 
32'd193808: dataIn1 = 32'd3171
; 
32'd193809: dataIn1 = 32'd11060
; 
32'd193810: dataIn1 = 32'd11061
; 
32'd193811: dataIn1 = 32'd11062
; 
32'd193812: dataIn1 = 32'd2852
; 
32'd193813: dataIn1 = 32'd3170
; 
32'd193814: dataIn1 = 32'd11061
; 
32'd193815: dataIn1 = 32'd11062
; 
32'd193816: dataIn1 = 32'd11063
; 
32'd193817: dataIn1 = 32'd2852
; 
32'd193818: dataIn1 = 32'd2854
; 
32'd193819: dataIn1 = 32'd11062
; 
32'd193820: dataIn1 = 32'd11063
; 
32'd193821: dataIn1 = 32'd11064
; 
32'd193822: dataIn1 = 32'd2854
; 
32'd193823: dataIn1 = 32'd3180
; 
32'd193824: dataIn1 = 32'd11063
; 
32'd193825: dataIn1 = 32'd11064
; 
32'd193826: dataIn1 = 32'd11065
; 
32'd193827: dataIn1 = 32'd3179
; 
32'd193828: dataIn1 = 32'd3180
; 
32'd193829: dataIn1 = 32'd11064
; 
32'd193830: dataIn1 = 32'd11065
; 
32'd193831: dataIn1 = 32'd11066
; 
32'd193832: dataIn1 = 32'd2864
; 
32'd193833: dataIn1 = 32'd3179
; 
32'd193834: dataIn1 = 32'd11065
; 
32'd193835: dataIn1 = 32'd11066
; 
32'd193836: dataIn1 = 32'd11067
; 
32'd193837: dataIn1 = 32'd2863
; 
32'd193838: dataIn1 = 32'd2864
; 
32'd193839: dataIn1 = 32'd11066
; 
32'd193840: dataIn1 = 32'd11067
; 
32'd193841: dataIn1 = 32'd11068
; 
32'd193842: dataIn1 = 32'd2863
; 
32'd193843: dataIn1 = 32'd3186
; 
32'd193844: dataIn1 = 32'd11067
; 
32'd193845: dataIn1 = 32'd11068
; 
32'd193846: dataIn1 = 32'd11069
; 
32'd193847: dataIn1 = 32'd3186
; 
32'd193848: dataIn1 = 32'd3187
; 
32'd193849: dataIn1 = 32'd11068
; 
32'd193850: dataIn1 = 32'd11069
; 
32'd193851: dataIn1 = 32'd11070
; 
32'd193852: dataIn1 = 32'd2869
; 
32'd193853: dataIn1 = 32'd3187
; 
32'd193854: dataIn1 = 32'd11069
; 
32'd193855: dataIn1 = 32'd11070
; 
32'd193856: dataIn1 = 32'd11071
; 
32'd193857: dataIn1 = 32'd2867
; 
32'd193858: dataIn1 = 32'd2869
; 
32'd193859: dataIn1 = 32'd11070
; 
32'd193860: dataIn1 = 32'd11071
; 
32'd193861: dataIn1 = 32'd11072
; 
32'd193862: dataIn1 = 32'd2867
; 
32'd193863: dataIn1 = 32'd3191
; 
32'd193864: dataIn1 = 32'd11071
; 
32'd193865: dataIn1 = 32'd11072
; 
32'd193866: dataIn1 = 32'd11073
; 
32'd193867: dataIn1 = 32'd3191
; 
32'd193868: dataIn1 = 32'd3192
; 
32'd193869: dataIn1 = 32'd11072
; 
32'd193870: dataIn1 = 32'd11073
; 
32'd193871: dataIn1 = 32'd11074
; 
32'd193872: dataIn1 = 32'd2889
; 
32'd193873: dataIn1 = 32'd3192
; 
32'd193874: dataIn1 = 32'd11073
; 
32'd193875: dataIn1 = 32'd11074
; 
32'd193876: dataIn1 = 32'd11075
; 
32'd193877: dataIn1 = 32'd2888
; 
32'd193878: dataIn1 = 32'd2889
; 
32'd193879: dataIn1 = 32'd11074
; 
32'd193880: dataIn1 = 32'd11075
; 
32'd193881: dataIn1 = 32'd11076
; 
32'd193882: dataIn1 = 32'd2888
; 
32'd193883: dataIn1 = 32'd3220
; 
32'd193884: dataIn1 = 32'd11075
; 
32'd193885: dataIn1 = 32'd11076
; 
32'd193886: dataIn1 = 32'd11077
; 
32'd193887: dataIn1 = 32'd3220
; 
32'd193888: dataIn1 = 32'd3221
; 
32'd193889: dataIn1 = 32'd11076
; 
32'd193890: dataIn1 = 32'd11077
; 
32'd193891: dataIn1 = 32'd11078
; 
32'd193892: dataIn1 = 32'd2878
; 
32'd193893: dataIn1 = 32'd3221
; 
32'd193894: dataIn1 = 32'd11077
; 
32'd193895: dataIn1 = 32'd11078
; 
32'd193896: dataIn1 = 32'd11079
; 
32'd193897: dataIn1 = 32'd2877
; 
32'd193898: dataIn1 = 32'd2878
; 
32'd193899: dataIn1 = 32'd11078
; 
32'd193900: dataIn1 = 32'd11079
; 
32'd193901: dataIn1 = 32'd11080
; 
32'd193902: dataIn1 = 32'd2877
; 
32'd193903: dataIn1 = 32'd3213
; 
32'd193904: dataIn1 = 32'd11079
; 
32'd193905: dataIn1 = 32'd11080
; 
32'd193906: dataIn1 = 32'd11081
; 
32'd193907: dataIn1 = 32'd3212
; 
32'd193908: dataIn1 = 32'd3213
; 
32'd193909: dataIn1 = 32'd11080
; 
32'd193910: dataIn1 = 32'd11081
; 
32'd193911: dataIn1 = 32'd11082
; 
32'd193912: dataIn1 = 32'd2882
; 
32'd193913: dataIn1 = 32'd3212
; 
32'd193914: dataIn1 = 32'd11081
; 
32'd193915: dataIn1 = 32'd11082
; 
32'd193916: dataIn1 = 32'd11083
; 
32'd193917: dataIn1 = 32'd2882
; 
32'd193918: dataIn1 = 32'd2884
; 
32'd193919: dataIn1 = 32'd11082
; 
32'd193920: dataIn1 = 32'd11083
; 
32'd193921: dataIn1 = 32'd11084
; 
32'd193922: dataIn1 = 32'd2884
; 
32'd193923: dataIn1 = 32'd3208
; 
32'd193924: dataIn1 = 32'd11083
; 
32'd193925: dataIn1 = 32'd11084
; 
32'd193926: dataIn1 = 32'd11085
; 
32'd193927: dataIn1 = 32'd3207
; 
32'd193928: dataIn1 = 32'd3208
; 
32'd193929: dataIn1 = 32'd11084
; 
32'd193930: dataIn1 = 32'd11085
; 
32'd193931: dataIn1 = 32'd11086
; 
32'd193932: dataIn1 = 32'd2874
; 
32'd193933: dataIn1 = 32'd3207
; 
32'd193934: dataIn1 = 32'd11085
; 
32'd193935: dataIn1 = 32'd11086
; 
32'd193936: dataIn1 = 32'd11087
; 
32'd193937: dataIn1 = 32'd2873
; 
32'd193938: dataIn1 = 32'd2874
; 
32'd193939: dataIn1 = 32'd11086
; 
32'd193940: dataIn1 = 32'd11087
; 
32'd193941: dataIn1 = 32'd11088
; 
32'd193942: dataIn1 = 32'd2873
; 
32'd193943: dataIn1 = 32'd3199
; 
32'd193944: dataIn1 = 32'd11087
; 
32'd193945: dataIn1 = 32'd11088
; 
32'd193946: dataIn1 = 32'd11089
; 
32'd193947: dataIn1 = 32'd3199
; 
32'd193948: dataIn1 = 32'd3200
; 
32'd193949: dataIn1 = 32'd11088
; 
32'd193950: dataIn1 = 32'd11089
; 
32'd193951: dataIn1 = 32'd11090
; 
32'd193952: dataIn1 = 32'd2898
; 
32'd193953: dataIn1 = 32'd3200
; 
32'd193954: dataIn1 = 32'd11089
; 
32'd193955: dataIn1 = 32'd11090
; 
32'd193956: dataIn1 = 32'd11091
; 
32'd193957: dataIn1 = 32'd2897
; 
32'd193958: dataIn1 = 32'd2898
; 
32'd193959: dataIn1 = 32'd11090
; 
32'd193960: dataIn1 = 32'd11091
; 
32'd193961: dataIn1 = 32'd11092
; 
32'd193962: dataIn1 = 32'd2897
; 
32'd193963: dataIn1 = 32'd3227
; 
32'd193964: dataIn1 = 32'd11091
; 
32'd193965: dataIn1 = 32'd11092
; 
32'd193966: dataIn1 = 32'd11093
; 
32'd193967: dataIn1 = 32'd3226
; 
32'd193968: dataIn1 = 32'd3227
; 
32'd193969: dataIn1 = 32'd11092
; 
32'd193970: dataIn1 = 32'd11093
; 
32'd193971: dataIn1 = 32'd11094
; 
32'd193972: dataIn1 = 32'd2892
; 
32'd193973: dataIn1 = 32'd3226
; 
32'd193974: dataIn1 = 32'd11093
; 
32'd193975: dataIn1 = 32'd11094
; 
32'd193976: dataIn1 = 32'd11095
; 
32'd193977: dataIn1 = 32'd2892
; 
32'd193978: dataIn1 = 32'd2894
; 
32'd193979: dataIn1 = 32'd11094
; 
32'd193980: dataIn1 = 32'd11095
; 
32'd193981: dataIn1 = 32'd11096
; 
32'd193982: dataIn1 = 32'd2894
; 
32'd193983: dataIn1 = 32'd3236
; 
32'd193984: dataIn1 = 32'd11095
; 
32'd193985: dataIn1 = 32'd11096
; 
32'd193986: dataIn1 = 32'd11097
; 
32'd193987: dataIn1 = 32'd3235
; 
32'd193988: dataIn1 = 32'd3236
; 
32'd193989: dataIn1 = 32'd11096
; 
32'd193990: dataIn1 = 32'd11097
; 
32'd193991: dataIn1 = 32'd11098
; 
32'd193992: dataIn1 = 32'd2904
; 
32'd193993: dataIn1 = 32'd3235
; 
32'd193994: dataIn1 = 32'd11097
; 
32'd193995: dataIn1 = 32'd11098
; 
32'd193996: dataIn1 = 32'd11099
; 
32'd193997: dataIn1 = 32'd2903
; 
32'd193998: dataIn1 = 32'd2904
; 
32'd193999: dataIn1 = 32'd11098
; 
32'd194000: dataIn1 = 32'd11099
; 
32'd194001: dataIn1 = 32'd11100
; 
32'd194002: dataIn1 = 32'd2903
; 
32'd194003: dataIn1 = 32'd3242
; 
32'd194004: dataIn1 = 32'd11099
; 
32'd194005: dataIn1 = 32'd11100
; 
32'd194006: dataIn1 = 32'd11101
; 
32'd194007: dataIn1 = 32'd3242
; 
32'd194008: dataIn1 = 32'd3243
; 
32'd194009: dataIn1 = 32'd11100
; 
32'd194010: dataIn1 = 32'd11101
; 
32'd194011: dataIn1 = 32'd11102
; 
32'd194012: dataIn1 = 32'd2909
; 
32'd194013: dataIn1 = 32'd3243
; 
32'd194014: dataIn1 = 32'd11101
; 
32'd194015: dataIn1 = 32'd11102
; 
32'd194016: dataIn1 = 32'd11103
; 
32'd194017: dataIn1 = 32'd2907
; 
32'd194018: dataIn1 = 32'd2909
; 
32'd194019: dataIn1 = 32'd11102
; 
32'd194020: dataIn1 = 32'd11103
; 
32'd194021: dataIn1 = 32'd11104
; 
32'd194022: dataIn1 = 32'd2907
; 
32'd194023: dataIn1 = 32'd3247
; 
32'd194024: dataIn1 = 32'd11103
; 
32'd194025: dataIn1 = 32'd11104
; 
32'd194026: dataIn1 = 32'd11105
; 
32'd194027: dataIn1 = 32'd3247
; 
32'd194028: dataIn1 = 32'd3248
; 
32'd194029: dataIn1 = 32'd11104
; 
32'd194030: dataIn1 = 32'd11105
; 
32'd194031: dataIn1 = 32'd11106
; 
32'd194032: dataIn1 = 32'd2929
; 
32'd194033: dataIn1 = 32'd3248
; 
32'd194034: dataIn1 = 32'd11105
; 
32'd194035: dataIn1 = 32'd11106
; 
32'd194036: dataIn1 = 32'd11107
; 
32'd194037: dataIn1 = 32'd2928
; 
32'd194038: dataIn1 = 32'd2929
; 
32'd194039: dataIn1 = 32'd11106
; 
32'd194040: dataIn1 = 32'd11107
; 
32'd194041: dataIn1 = 32'd11108
; 
32'd194042: dataIn1 = 32'd2928
; 
32'd194043: dataIn1 = 32'd3276
; 
32'd194044: dataIn1 = 32'd11107
; 
32'd194045: dataIn1 = 32'd11108
; 
32'd194046: dataIn1 = 32'd11109
; 
32'd194047: dataIn1 = 32'd3276
; 
32'd194048: dataIn1 = 32'd3277
; 
32'd194049: dataIn1 = 32'd11108
; 
32'd194050: dataIn1 = 32'd11109
; 
32'd194051: dataIn1 = 32'd11110
; 
32'd194052: dataIn1 = 32'd2918
; 
32'd194053: dataIn1 = 32'd3277
; 
32'd194054: dataIn1 = 32'd11109
; 
32'd194055: dataIn1 = 32'd11110
; 
32'd194056: dataIn1 = 32'd11111
; 
32'd194057: dataIn1 = 32'd2917
; 
32'd194058: dataIn1 = 32'd2918
; 
32'd194059: dataIn1 = 32'd11110
; 
32'd194060: dataIn1 = 32'd11111
; 
32'd194061: dataIn1 = 32'd11112
; 
32'd194062: dataIn1 = 32'd2917
; 
32'd194063: dataIn1 = 32'd3269
; 
32'd194064: dataIn1 = 32'd11111
; 
32'd194065: dataIn1 = 32'd11112
; 
32'd194066: dataIn1 = 32'd11113
; 
32'd194067: dataIn1 = 32'd3268
; 
32'd194068: dataIn1 = 32'd3269
; 
32'd194069: dataIn1 = 32'd11112
; 
32'd194070: dataIn1 = 32'd11113
; 
32'd194071: dataIn1 = 32'd11114
; 
32'd194072: dataIn1 = 32'd2922
; 
32'd194073: dataIn1 = 32'd3268
; 
32'd194074: dataIn1 = 32'd11113
; 
32'd194075: dataIn1 = 32'd11114
; 
32'd194076: dataIn1 = 32'd11115
; 
32'd194077: dataIn1 = 32'd2922
; 
32'd194078: dataIn1 = 32'd2924
; 
32'd194079: dataIn1 = 32'd11114
; 
32'd194080: dataIn1 = 32'd11115
; 
32'd194081: dataIn1 = 32'd11116
; 
32'd194082: dataIn1 = 32'd2924
; 
32'd194083: dataIn1 = 32'd3264
; 
32'd194084: dataIn1 = 32'd11115
; 
32'd194085: dataIn1 = 32'd11116
; 
32'd194086: dataIn1 = 32'd11117
; 
32'd194087: dataIn1 = 32'd3263
; 
32'd194088: dataIn1 = 32'd3264
; 
32'd194089: dataIn1 = 32'd11116
; 
32'd194090: dataIn1 = 32'd11117
; 
32'd194091: dataIn1 = 32'd11118
; 
32'd194092: dataIn1 = 32'd2914
; 
32'd194093: dataIn1 = 32'd3263
; 
32'd194094: dataIn1 = 32'd11117
; 
32'd194095: dataIn1 = 32'd11118
; 
32'd194096: dataIn1 = 32'd11119
; 
32'd194097: dataIn1 = 32'd2913
; 
32'd194098: dataIn1 = 32'd2914
; 
32'd194099: dataIn1 = 32'd11118
; 
32'd194100: dataIn1 = 32'd11119
; 
32'd194101: dataIn1 = 32'd11120
; 
32'd194102: dataIn1 = 32'd2913
; 
32'd194103: dataIn1 = 32'd3255
; 
32'd194104: dataIn1 = 32'd11119
; 
32'd194105: dataIn1 = 32'd11120
; 
32'd194106: dataIn1 = 32'd11121
; 
32'd194107: dataIn1 = 32'd3255
; 
32'd194108: dataIn1 = 32'd3256
; 
32'd194109: dataIn1 = 32'd11120
; 
32'd194110: dataIn1 = 32'd11121
; 
32'd194111: dataIn1 = 32'd11122
; 
32'd194112: dataIn1 = 32'd2938
; 
32'd194113: dataIn1 = 32'd3256
; 
32'd194114: dataIn1 = 32'd11121
; 
32'd194115: dataIn1 = 32'd11122
; 
32'd194116: dataIn1 = 32'd11123
; 
32'd194117: dataIn1 = 32'd2937
; 
32'd194118: dataIn1 = 32'd2938
; 
32'd194119: dataIn1 = 32'd11122
; 
32'd194120: dataIn1 = 32'd11123
; 
32'd194121: dataIn1 = 32'd11124
; 
32'd194122: dataIn1 = 32'd2937
; 
32'd194123: dataIn1 = 32'd3283
; 
32'd194124: dataIn1 = 32'd11123
; 
32'd194125: dataIn1 = 32'd11124
; 
32'd194126: dataIn1 = 32'd11125
; 
32'd194127: dataIn1 = 32'd3282
; 
32'd194128: dataIn1 = 32'd3283
; 
32'd194129: dataIn1 = 32'd11124
; 
32'd194130: dataIn1 = 32'd11125
; 
32'd194131: dataIn1 = 32'd11126
; 
32'd194132: dataIn1 = 32'd2932
; 
32'd194133: dataIn1 = 32'd3282
; 
32'd194134: dataIn1 = 32'd11125
; 
32'd194135: dataIn1 = 32'd11126
; 
32'd194136: dataIn1 = 32'd11127
; 
32'd194137: dataIn1 = 32'd2932
; 
32'd194138: dataIn1 = 32'd2934
; 
32'd194139: dataIn1 = 32'd11126
; 
32'd194140: dataIn1 = 32'd11127
; 
32'd194141: dataIn1 = 32'd11128
; 
32'd194142: dataIn1 = 32'd2934
; 
32'd194143: dataIn1 = 32'd3292
; 
32'd194144: dataIn1 = 32'd11127
; 
32'd194145: dataIn1 = 32'd11128
; 
32'd194146: dataIn1 = 32'd11129
; 
32'd194147: dataIn1 = 32'd3291
; 
32'd194148: dataIn1 = 32'd3292
; 
32'd194149: dataIn1 = 32'd11128
; 
32'd194150: dataIn1 = 32'd11129
; 
32'd194151: dataIn1 = 32'd11130
; 
32'd194152: dataIn1 = 32'd2944
; 
32'd194153: dataIn1 = 32'd3291
; 
32'd194154: dataIn1 = 32'd11129
; 
32'd194155: dataIn1 = 32'd11130
; 
32'd194156: dataIn1 = 32'd11131
; 
32'd194157: dataIn1 = 32'd2943
; 
32'd194158: dataIn1 = 32'd2944
; 
32'd194159: dataIn1 = 32'd11130
; 
32'd194160: dataIn1 = 32'd11131
; 
32'd194161: dataIn1 = 32'd11132
; 
32'd194162: dataIn1 = 32'd2943
; 
32'd194163: dataIn1 = 32'd3298
; 
32'd194164: dataIn1 = 32'd11131
; 
32'd194165: dataIn1 = 32'd11132
; 
32'd194166: dataIn1 = 32'd11133
; 
32'd194167: dataIn1 = 32'd3298
; 
32'd194168: dataIn1 = 32'd3299
; 
32'd194169: dataIn1 = 32'd11132
; 
32'd194170: dataIn1 = 32'd11133
; 
32'd194171: dataIn1 = 32'd11134
; 
32'd194172: dataIn1 = 32'd2949
; 
32'd194173: dataIn1 = 32'd3299
; 
32'd194174: dataIn1 = 32'd11133
; 
32'd194175: dataIn1 = 32'd11134
; 
32'd194176: dataIn1 = 32'd11135
; 
32'd194177: dataIn1 = 32'd2947
; 
32'd194178: dataIn1 = 32'd2949
; 
32'd194179: dataIn1 = 32'd11134
; 
32'd194180: dataIn1 = 32'd11135
; 
32'd194181: dataIn1 = 32'd11136
; 
32'd194182: dataIn1 = 32'd2947
; 
32'd194183: dataIn1 = 32'd3303
; 
32'd194184: dataIn1 = 32'd11135
; 
32'd194185: dataIn1 = 32'd11136
; 
32'd194186: dataIn1 = 32'd11137
; 
32'd194187: dataIn1 = 32'd3303
; 
32'd194188: dataIn1 = 32'd3304
; 
32'd194189: dataIn1 = 32'd11136
; 
32'd194190: dataIn1 = 32'd11137
; 
32'd194191: dataIn1 = 32'd11138
; 
32'd194192: dataIn1 = 32'd2969
; 
32'd194193: dataIn1 = 32'd3304
; 
32'd194194: dataIn1 = 32'd11137
; 
32'd194195: dataIn1 = 32'd11138
; 
32'd194196: dataIn1 = 32'd11139
; 
32'd194197: dataIn1 = 32'd2968
; 
32'd194198: dataIn1 = 32'd2969
; 
32'd194199: dataIn1 = 32'd11138
; 
32'd194200: dataIn1 = 32'd11139
; 
32'd194201: dataIn1 = 32'd11140
; 
32'd194202: dataIn1 = 32'd2968
; 
32'd194203: dataIn1 = 32'd3332
; 
32'd194204: dataIn1 = 32'd11139
; 
32'd194205: dataIn1 = 32'd11140
; 
32'd194206: dataIn1 = 32'd11141
; 
32'd194207: dataIn1 = 32'd3332
; 
32'd194208: dataIn1 = 32'd3333
; 
32'd194209: dataIn1 = 32'd11140
; 
32'd194210: dataIn1 = 32'd11141
; 
32'd194211: dataIn1 = 32'd11142
; 
32'd194212: dataIn1 = 32'd2958
; 
32'd194213: dataIn1 = 32'd3333
; 
32'd194214: dataIn1 = 32'd11141
; 
32'd194215: dataIn1 = 32'd11142
; 
32'd194216: dataIn1 = 32'd11143
; 
32'd194217: dataIn1 = 32'd2957
; 
32'd194218: dataIn1 = 32'd2958
; 
32'd194219: dataIn1 = 32'd11142
; 
32'd194220: dataIn1 = 32'd11143
; 
32'd194221: dataIn1 = 32'd11144
; 
32'd194222: dataIn1 = 32'd2957
; 
32'd194223: dataIn1 = 32'd3325
; 
32'd194224: dataIn1 = 32'd11143
; 
32'd194225: dataIn1 = 32'd11144
; 
32'd194226: dataIn1 = 32'd11145
; 
32'd194227: dataIn1 = 32'd3324
; 
32'd194228: dataIn1 = 32'd3325
; 
32'd194229: dataIn1 = 32'd11144
; 
32'd194230: dataIn1 = 32'd11145
; 
32'd194231: dataIn1 = 32'd11146
; 
32'd194232: dataIn1 = 32'd2962
; 
32'd194233: dataIn1 = 32'd3324
; 
32'd194234: dataIn1 = 32'd11145
; 
32'd194235: dataIn1 = 32'd11146
; 
32'd194236: dataIn1 = 32'd11147
; 
32'd194237: dataIn1 = 32'd2962
; 
32'd194238: dataIn1 = 32'd2964
; 
32'd194239: dataIn1 = 32'd11146
; 
32'd194240: dataIn1 = 32'd11147
; 
32'd194241: dataIn1 = 32'd11148
; 
32'd194242: dataIn1 = 32'd2964
; 
32'd194243: dataIn1 = 32'd3320
; 
32'd194244: dataIn1 = 32'd11147
; 
32'd194245: dataIn1 = 32'd11148
; 
32'd194246: dataIn1 = 32'd11149
; 
32'd194247: dataIn1 = 32'd3319
; 
32'd194248: dataIn1 = 32'd3320
; 
32'd194249: dataIn1 = 32'd11148
; 
32'd194250: dataIn1 = 32'd11149
; 
32'd194251: dataIn1 = 32'd11150
; 
32'd194252: dataIn1 = 32'd2954
; 
32'd194253: dataIn1 = 32'd3319
; 
32'd194254: dataIn1 = 32'd11149
; 
32'd194255: dataIn1 = 32'd11150
; 
32'd194256: dataIn1 = 32'd11151
; 
32'd194257: dataIn1 = 32'd2953
; 
32'd194258: dataIn1 = 32'd2954
; 
32'd194259: dataIn1 = 32'd11150
; 
32'd194260: dataIn1 = 32'd11151
; 
32'd194261: dataIn1 = 32'd11152
; 
32'd194262: dataIn1 = 32'd2953
; 
32'd194263: dataIn1 = 32'd3311
; 
32'd194264: dataIn1 = 32'd11151
; 
32'd194265: dataIn1 = 32'd11152
; 
32'd194266: dataIn1 = 32'd11153
; 
32'd194267: dataIn1 = 32'd3311
; 
32'd194268: dataIn1 = 32'd3312
; 
32'd194269: dataIn1 = 32'd11152
; 
32'd194270: dataIn1 = 32'd11153
; 
32'd194271: dataIn1 = 32'd11154
; 
32'd194272: dataIn1 = 32'd2978
; 
32'd194273: dataIn1 = 32'd3312
; 
32'd194274: dataIn1 = 32'd11153
; 
32'd194275: dataIn1 = 32'd11154
; 
32'd194276: dataIn1 = 32'd11155
; 
32'd194277: dataIn1 = 32'd2977
; 
32'd194278: dataIn1 = 32'd2978
; 
32'd194279: dataIn1 = 32'd11154
; 
32'd194280: dataIn1 = 32'd11155
; 
32'd194281: dataIn1 = 32'd11156
; 
32'd194282: dataIn1 = 32'd2977
; 
32'd194283: dataIn1 = 32'd3339
; 
32'd194284: dataIn1 = 32'd11155
; 
32'd194285: dataIn1 = 32'd11156
; 
32'd194286: dataIn1 = 32'd11157
; 
32'd194287: dataIn1 = 32'd3338
; 
32'd194288: dataIn1 = 32'd3339
; 
32'd194289: dataIn1 = 32'd11156
; 
32'd194290: dataIn1 = 32'd11157
; 
32'd194291: dataIn1 = 32'd11158
; 
32'd194292: dataIn1 = 32'd2972
; 
32'd194293: dataIn1 = 32'd3338
; 
32'd194294: dataIn1 = 32'd11157
; 
32'd194295: dataIn1 = 32'd11158
; 
32'd194296: dataIn1 = 32'd11159
; 
32'd194297: dataIn1 = 32'd2972
; 
32'd194298: dataIn1 = 32'd2974
; 
32'd194299: dataIn1 = 32'd11158
; 
32'd194300: dataIn1 = 32'd11159
; 
32'd194301: dataIn1 = 32'd11160
; 
32'd194302: dataIn1 = 32'd2974
; 
32'd194303: dataIn1 = 32'd3348
; 
32'd194304: dataIn1 = 32'd11159
; 
32'd194305: dataIn1 = 32'd11160
; 
32'd194306: dataIn1 = 32'd11161
; 
32'd194307: dataIn1 = 32'd3347
; 
32'd194308: dataIn1 = 32'd3348
; 
32'd194309: dataIn1 = 32'd11160
; 
32'd194310: dataIn1 = 32'd11161
; 
32'd194311: dataIn1 = 32'd11162
; 
32'd194312: dataIn1 = 32'd2984
; 
32'd194313: dataIn1 = 32'd3347
; 
32'd194314: dataIn1 = 32'd11161
; 
32'd194315: dataIn1 = 32'd11162
; 
32'd194316: dataIn1 = 32'd11163
; 
32'd194317: dataIn1 = 32'd2983
; 
32'd194318: dataIn1 = 32'd2984
; 
32'd194319: dataIn1 = 32'd11162
; 
32'd194320: dataIn1 = 32'd11163
; 
32'd194321: dataIn1 = 32'd11164
; 
32'd194322: dataIn1 = 32'd2983
; 
32'd194323: dataIn1 = 32'd3354
; 
32'd194324: dataIn1 = 32'd11163
; 
32'd194325: dataIn1 = 32'd11164
; 
32'd194326: dataIn1 = 32'd11165
; 
32'd194327: dataIn1 = 32'd3354
; 
32'd194328: dataIn1 = 32'd3355
; 
32'd194329: dataIn1 = 32'd11164
; 
32'd194330: dataIn1 = 32'd11165
; 
32'd194331: dataIn1 = 32'd11166
; 
32'd194332: dataIn1 = 32'd2989
; 
32'd194333: dataIn1 = 32'd3355
; 
32'd194334: dataIn1 = 32'd11165
; 
32'd194335: dataIn1 = 32'd11166
; 
32'd194336: dataIn1 = 32'd11167
; 
32'd194337: dataIn1 = 32'd2987
; 
32'd194338: dataIn1 = 32'd2989
; 
32'd194339: dataIn1 = 32'd11166
; 
32'd194340: dataIn1 = 32'd11167
; 
32'd194341: dataIn1 = 32'd11168
; 
32'd194342: dataIn1 = 32'd2987
; 
32'd194343: dataIn1 = 32'd3359
; 
32'd194344: dataIn1 = 32'd11167
; 
32'd194345: dataIn1 = 32'd11168
; 
32'd194346: dataIn1 = 32'd11169
; 
32'd194347: dataIn1 = 32'd3359
; 
32'd194348: dataIn1 = 32'd3360
; 
32'd194349: dataIn1 = 32'd11168
; 
32'd194350: dataIn1 = 32'd11169
; 
32'd194351: dataIn1 = 32'd11170
; 
32'd194352: dataIn1 = 32'd3360
; 
32'd194353: dataIn1 = 32'd11169
; 
32'd194354: dataIn1 = 32'd11170
; 
32'd194355: dataIn1 = 32'd11171
; 
32'd194356: dataIn1 = 32'd3009
; 
32'd194357: dataIn1 = 32'd3360
; 
32'd194358: dataIn1 = 32'd11170
; 
32'd194359: dataIn1 = 32'd11171
; 
32'd194360: dataIn1 = 32'd11172
; 
32'd194361: dataIn1 = 32'd3008
; 
32'd194362: dataIn1 = 32'd3009
; 
32'd194363: dataIn1 = 32'd3388
; 
32'd194364: dataIn1 = 32'd11171
; 
32'd194365: dataIn1 = 32'd11172
; 
32'd194366: dataIn1 = 32'd11173
; 
32'd194367: dataIn1 = 32'd3388
; 
32'd194368: dataIn1 = 32'd3389
; 
32'd194369: dataIn1 = 32'd11172
; 
32'd194370: dataIn1 = 32'd11173
; 
32'd194371: dataIn1 = 32'd11174
; 
32'd194372: dataIn1 = 32'd2998
; 
32'd194373: dataIn1 = 32'd3389
; 
32'd194374: dataIn1 = 32'd11173
; 
32'd194375: dataIn1 = 32'd11174
; 
32'd194376: dataIn1 = 32'd11175
; 
32'd194377: dataIn1 = 32'd2997
; 
32'd194378: dataIn1 = 32'd2998
; 
32'd194379: dataIn1 = 32'd11174
; 
32'd194380: dataIn1 = 32'd11175
; 
32'd194381: dataIn1 = 32'd11176
; 
32'd194382: dataIn1 = 32'd2997
; 
32'd194383: dataIn1 = 32'd3381
; 
32'd194384: dataIn1 = 32'd11175
; 
32'd194385: dataIn1 = 32'd11176
; 
32'd194386: dataIn1 = 32'd11177
; 
32'd194387: dataIn1 = 32'd3380
; 
32'd194388: dataIn1 = 32'd3381
; 
32'd194389: dataIn1 = 32'd11176
; 
32'd194390: dataIn1 = 32'd11177
; 
32'd194391: dataIn1 = 32'd11178
; 
32'd194392: dataIn1 = 32'd3002
; 
32'd194393: dataIn1 = 32'd3380
; 
32'd194394: dataIn1 = 32'd11177
; 
32'd194395: dataIn1 = 32'd11178
; 
32'd194396: dataIn1 = 32'd11179
; 
32'd194397: dataIn1 = 32'd3002
; 
32'd194398: dataIn1 = 32'd11178
; 
32'd194399: dataIn1 = 32'd11179
; 
32'd194400: dataIn1 = 32'd11180
; 
32'd194401: dataIn1 = 32'd3002
; 
32'd194402: dataIn1 = 32'd3004
; 
32'd194403: dataIn1 = 32'd11179
; 
32'd194404: dataIn1 = 32'd11180
; 
32'd194405: dataIn1 = 32'd11181
; 
32'd194406: dataIn1 = 32'd3004
; 
32'd194407: dataIn1 = 32'd3376
; 
32'd194408: dataIn1 = 32'd11180
; 
32'd194409: dataIn1 = 32'd11181
; 
32'd194410: dataIn1 = 32'd11182
; 
32'd194411: dataIn1 = 32'd3375
; 
32'd194412: dataIn1 = 32'd3376
; 
32'd194413: dataIn1 = 32'd11181
; 
32'd194414: dataIn1 = 32'd11182
; 
32'd194415: dataIn1 = 32'd11183
; 
32'd194416: dataIn1 = 32'd2994
; 
32'd194417: dataIn1 = 32'd3375
; 
32'd194418: dataIn1 = 32'd11182
; 
32'd194419: dataIn1 = 32'd11183
; 
32'd194420: dataIn1 = 32'd11184
; 
32'd194421: dataIn1 = 32'd2993
; 
32'd194422: dataIn1 = 32'd2994
; 
32'd194423: dataIn1 = 32'd11183
; 
32'd194424: dataIn1 = 32'd11184
; 
32'd194425: dataIn1 = 32'd11185
; 
32'd194426: dataIn1 = 32'd2993
; 
32'd194427: dataIn1 = 32'd3367
; 
32'd194428: dataIn1 = 32'd11184
; 
32'd194429: dataIn1 = 32'd11185
; 
32'd194430: dataIn1 = 32'd11186
; 
32'd194431: dataIn1 = 32'd3367
; 
32'd194432: dataIn1 = 32'd3368
; 
32'd194433: dataIn1 = 32'd11185
; 
32'd194434: dataIn1 = 32'd11186
; 
32'd194435: dataIn1 = 32'd11187
; 
32'd194436: dataIn1 = 32'd3018
; 
32'd194437: dataIn1 = 32'd3368
; 
32'd194438: dataIn1 = 32'd11186
; 
32'd194439: dataIn1 = 32'd11187
; 
32'd194440: dataIn1 = 32'd11188
; 
32'd194441: dataIn1 = 32'd3017
; 
32'd194442: dataIn1 = 32'd3018
; 
32'd194443: dataIn1 = 32'd11187
; 
32'd194444: dataIn1 = 32'd11188
; 
32'd194445: dataIn1 = 32'd11189
; 
32'd194446: dataIn1 = 32'd3017
; 
32'd194447: dataIn1 = 32'd3395
; 
32'd194448: dataIn1 = 32'd11188
; 
32'd194449: dataIn1 = 32'd11189
; 
32'd194450: dataIn1 = 32'd11190
; 
32'd194451: dataIn1 = 32'd3394
; 
32'd194452: dataIn1 = 32'd3395
; 
32'd194453: dataIn1 = 32'd11189
; 
32'd194454: dataIn1 = 32'd11190
; 
32'd194455: dataIn1 = 32'd11191
; 
32'd194456: dataIn1 = 32'd3012
; 
32'd194457: dataIn1 = 32'd3394
; 
32'd194458: dataIn1 = 32'd11190
; 
32'd194459: dataIn1 = 32'd11191
; 
32'd194460: dataIn1 = 32'd11192
; 
32'd194461: dataIn1 = 32'd3012
; 
32'd194462: dataIn1 = 32'd3014
; 
32'd194463: dataIn1 = 32'd11191
; 
32'd194464: dataIn1 = 32'd11192
; 
32'd194465: dataIn1 = 32'd11193
; 
32'd194466: dataIn1 = 32'd3014
; 
32'd194467: dataIn1 = 32'd3404
; 
32'd194468: dataIn1 = 32'd11192
; 
32'd194469: dataIn1 = 32'd11193
; 
32'd194470: dataIn1 = 32'd11194
; 
32'd194471: dataIn1 = 32'd3403
; 
32'd194472: dataIn1 = 32'd3404
; 
32'd194473: dataIn1 = 32'd11193
; 
32'd194474: dataIn1 = 32'd11194
; 
32'd194475: dataIn1 = 32'd11195
; 
32'd194476: dataIn1 = 32'd3023
; 
32'd194477: dataIn1 = 32'd3024
; 
32'd194478: dataIn1 = 32'd3403
; 
32'd194479: dataIn1 = 32'd11194
; 
32'd194480: dataIn1 = 32'd11195
; 
32'd194481: dataIn1 = 32'd11196
; 
32'd194482: dataIn1 = 32'd3023
; 
32'd194483: dataIn1 = 32'd11195
; 
32'd194484: dataIn1 = 32'd11196
; 
32'd194485: dataIn1 = 32'd11197
; 
32'd194486: dataIn1 = 32'd3023
; 
32'd194487: dataIn1 = 32'd3441
; 
32'd194488: dataIn1 = 32'd11196
; 
32'd194489: dataIn1 = 32'd11197
; 
32'd194490: dataIn1 = 32'd727
; 
32'd194491: dataIn1 = 32'd1395
; 
32'd194492: dataIn1 = 32'd10563
; 
32'd194493: dataIn1 = 32'd11198
; 
32'd194494: dataIn1 = 32'd11199
; 
32'd194495: dataIn1 = 32'd727
; 
32'd194496: dataIn1 = 32'd1394
; 
32'd194497: dataIn1 = 32'd11198
; 
32'd194498: dataIn1 = 32'd11199
; 
32'd194499: dataIn1 = 32'd11200
; 
32'd194500: dataIn1 = 32'd1394
; 
32'd194501: dataIn1 = 32'd11199
; 
32'd194502: dataIn1 = 32'd11200
; 
32'd194503: dataIn1 = 32'd11201
; 
32'd194504: dataIn1 = 32'd725
; 
32'd194505: dataIn1 = 32'd1394
; 
32'd194506: dataIn1 = 32'd11200
; 
32'd194507: dataIn1 = 32'd11201
; 
32'd194508: dataIn1 = 32'd11202
; 
32'd194509: dataIn1 = 32'd725
; 
32'd194510: dataIn1 = 32'd1392
; 
32'd194511: dataIn1 = 32'd11201
; 
32'd194512: dataIn1 = 32'd11202
; 
32'd194513: dataIn1 = 32'd11203
; 
32'd194514: dataIn1 = 32'd724
; 
32'd194515: dataIn1 = 32'd1392
; 
32'd194516: dataIn1 = 32'd11202
; 
32'd194517: dataIn1 = 32'd11203
; 
32'd194518: dataIn1 = 32'd11204
; 
32'd194519: dataIn1 = 32'd724
; 
32'd194520: dataIn1 = 32'd1393
; 
32'd194521: dataIn1 = 32'd11203
; 
32'd194522: dataIn1 = 32'd11204
; 
32'd194523: dataIn1 = 32'd11205
; 
32'd194524: dataIn1 = 32'd726
; 
32'd194525: dataIn1 = 32'd1393
; 
32'd194526: dataIn1 = 32'd11204
; 
32'd194527: dataIn1 = 32'd11205
; 
32'd194528: dataIn1 = 32'd11206
; 
32'd194529: dataIn1 = 32'd722
; 
32'd194530: dataIn1 = 32'd726
; 
32'd194531: dataIn1 = 32'd1396
; 
32'd194532: dataIn1 = 32'd11205
; 
32'd194533: dataIn1 = 32'd11206
; 
32'd194534: dataIn1 = 32'd11207
; 
32'd194535: dataIn1 = 32'd722
; 
32'd194536: dataIn1 = 32'd11206
; 
32'd194537: dataIn1 = 32'd11207
; 
32'd194538: dataIn1 = 32'd11208
; 
32'd194539: dataIn1 = 32'd722
; 
32'd194540: dataIn1 = 32'd1390
; 
32'd194541: dataIn1 = 32'd11207
; 
32'd194542: dataIn1 = 32'd11208
; 
32'd194543: dataIn1 = 32'd11209
; 
32'd194544: dataIn1 = 32'd1390
; 
32'd194545: dataIn1 = 32'd11208
; 
32'd194546: dataIn1 = 32'd11209
; 
32'd194547: dataIn1 = 32'd11210
; 
32'd194548: dataIn1 = 32'd720
; 
32'd194549: dataIn1 = 32'd1390
; 
32'd194550: dataIn1 = 32'd11209
; 
32'd194551: dataIn1 = 32'd11210
; 
32'd194552: dataIn1 = 32'd11211
; 
32'd194553: dataIn1 = 32'd720
; 
32'd194554: dataIn1 = 32'd11210
; 
32'd194555: dataIn1 = 32'd11211
; 
32'd194556: dataIn1 = 32'd11212
; 
32'd194557: dataIn1 = 32'd720
; 
32'd194558: dataIn1 = 32'd1389
; 
32'd194559: dataIn1 = 32'd11211
; 
32'd194560: dataIn1 = 32'd11212
; 
32'd194561: dataIn1 = 32'd11213
; 
32'd194562: dataIn1 = 32'd721
; 
32'd194563: dataIn1 = 32'd1389
; 
32'd194564: dataIn1 = 32'd11212
; 
32'd194565: dataIn1 = 32'd11213
; 
32'd194566: dataIn1 = 32'd11214
; 
32'd194567: dataIn1 = 32'd721
; 
32'd194568: dataIn1 = 32'd11213
; 
32'd194569: dataIn1 = 32'd11214
; 
32'd194570: dataIn1 = 32'd11215
; 
32'd194571: dataIn1 = 32'd721
; 
32'd194572: dataIn1 = 32'd11214
; 
32'd194573: dataIn1 = 32'd11215
; 
32'd194574: dataIn1 = 32'd11216
; 
32'd194575: dataIn1 = 32'd721
; 
32'd194576: dataIn1 = 32'd1391
; 
32'd194577: dataIn1 = 32'd11215
; 
32'd194578: dataIn1 = 32'd11216
; 
32'd194579: dataIn1 = 32'd11217
; 
32'd194580: dataIn1 = 32'd712
; 
32'd194581: dataIn1 = 32'd1391
; 
32'd194582: dataIn1 = 32'd11216
; 
32'd194583: dataIn1 = 32'd11217
; 
32'd194584: dataIn1 = 32'd11218
; 
32'd194585: dataIn1 = 32'd712
; 
32'd194586: dataIn1 = 32'd11217
; 
32'd194587: dataIn1 = 32'd11218
; 
32'd194588: dataIn1 = 32'd11219
; 
32'd194589: dataIn1 = 32'd712
; 
32'd194590: dataIn1 = 32'd11218
; 
32'd194591: dataIn1 = 32'd11219
; 
32'd194592: dataIn1 = 32'd11220
; 
32'd194593: dataIn1 = 32'd712
; 
32'd194594: dataIn1 = 32'd1384
; 
32'd194595: dataIn1 = 32'd11219
; 
32'd194596: dataIn1 = 32'd11220
; 
32'd194597: dataIn1 = 32'd11221
; 
32'd194598: dataIn1 = 32'd1384
; 
32'd194599: dataIn1 = 32'd11220
; 
32'd194600: dataIn1 = 32'd11221
; 
32'd194601: dataIn1 = 32'd11222
; 
32'd194602: dataIn1 = 32'd711
; 
32'd194603: dataIn1 = 32'd1384
; 
32'd194604: dataIn1 = 32'd11221
; 
32'd194605: dataIn1 = 32'd11222
; 
32'd194606: dataIn1 = 32'd11223
; 
32'd194607: dataIn1 = 32'd711
; 
32'd194608: dataIn1 = 32'd1383
; 
32'd194609: dataIn1 = 32'd11222
; 
32'd194610: dataIn1 = 32'd11223
; 
32'd194611: dataIn1 = 32'd11224
; 
32'd194612: dataIn1 = 32'd1383
; 
32'd194613: dataIn1 = 32'd11223
; 
32'd194614: dataIn1 = 32'd11224
; 
32'd194615: dataIn1 = 32'd11225
; 
32'd194616: dataIn1 = 32'd709
; 
32'd194617: dataIn1 = 32'd1383
; 
32'd194618: dataIn1 = 32'd11224
; 
32'd194619: dataIn1 = 32'd11225
; 
32'd194620: dataIn1 = 32'd11226
; 
32'd194621: dataIn1 = 32'd709
; 
32'd194622: dataIn1 = 32'd11225
; 
32'd194623: dataIn1 = 32'd11226
; 
32'd194624: dataIn1 = 32'd11227
; 
32'd194625: dataIn1 = 32'd709
; 
32'd194626: dataIn1 = 32'd1381
; 
32'd194627: dataIn1 = 32'd11226
; 
32'd194628: dataIn1 = 32'd11227
; 
32'd194629: dataIn1 = 32'd11228
; 
32'd194630: dataIn1 = 32'd1381
; 
32'd194631: dataIn1 = 32'd11227
; 
32'd194632: dataIn1 = 32'd11228
; 
32'd194633: dataIn1 = 32'd11229
; 
32'd194634: dataIn1 = 32'd707
; 
32'd194635: dataIn1 = 32'd1381
; 
32'd194636: dataIn1 = 32'd11228
; 
32'd194637: dataIn1 = 32'd11229
; 
32'd194638: dataIn1 = 32'd11230
; 
32'd194639: dataIn1 = 32'd707
; 
32'd194640: dataIn1 = 32'd11229
; 
32'd194641: dataIn1 = 32'd11230
; 
32'd194642: dataIn1 = 32'd11231
; 
32'd194643: dataIn1 = 32'd707
; 
32'd194644: dataIn1 = 32'd1382
; 
32'd194645: dataIn1 = 32'd11230
; 
32'd194646: dataIn1 = 32'd11231
; 
32'd194647: dataIn1 = 32'd11232
; 
32'd194648: dataIn1 = 32'd1382
; 
32'd194649: dataIn1 = 32'd11231
; 
32'd194650: dataIn1 = 32'd11232
; 
32'd194651: dataIn1 = 32'd11233
; 
32'd194652: dataIn1 = 32'd1382
; 
32'd194653: dataIn1 = 32'd11232
; 
32'd194654: dataIn1 = 32'd11233
; 
32'd194655: dataIn1 = 32'd11234
; 
32'd194656: dataIn1 = 32'd710
; 
32'd194657: dataIn1 = 32'd1382
; 
32'd194658: dataIn1 = 32'd11233
; 
32'd194659: dataIn1 = 32'd11234
; 
32'd194660: dataIn1 = 32'd11235
; 
32'd194661: dataIn1 = 32'd710
; 
32'd194662: dataIn1 = 32'd11234
; 
32'd194663: dataIn1 = 32'd11235
; 
32'd194664: dataIn1 = 32'd11236
; 
32'd194665: dataIn1 = 32'd710
; 
32'd194666: dataIn1 = 32'd1385
; 
32'd194667: dataIn1 = 32'd11235
; 
32'd194668: dataIn1 = 32'd11236
; 
32'd194669: dataIn1 = 32'd11237
; 
32'd194670: dataIn1 = 32'd715
; 
32'd194671: dataIn1 = 32'd1385
; 
32'd194672: dataIn1 = 32'd11236
; 
32'd194673: dataIn1 = 32'd11237
; 
32'd194674: dataIn1 = 32'd11238
; 
32'd194675: dataIn1 = 32'd715
; 
32'd194676: dataIn1 = 32'd11237
; 
32'd194677: dataIn1 = 32'd11238
; 
32'd194678: dataIn1 = 32'd11239
; 
32'd194679: dataIn1 = 32'd715
; 
32'd194680: dataIn1 = 32'd1387
; 
32'd194681: dataIn1 = 32'd11238
; 
32'd194682: dataIn1 = 32'd11239
; 
32'd194683: dataIn1 = 32'd11240
; 
32'd194684: dataIn1 = 32'd1387
; 
32'd194685: dataIn1 = 32'd11239
; 
32'd194686: dataIn1 = 32'd11240
; 
32'd194687: dataIn1 = 32'd11241
; 
32'd194688: dataIn1 = 32'd716
; 
32'd194689: dataIn1 = 32'd1387
; 
32'd194690: dataIn1 = 32'd11240
; 
32'd194691: dataIn1 = 32'd11241
; 
32'd194692: dataIn1 = 32'd11242
; 
32'd194693: dataIn1 = 32'd716
; 
32'd194694: dataIn1 = 32'd11241
; 
32'd194695: dataIn1 = 32'd11242
; 
32'd194696: dataIn1 = 32'd11243
; 
32'd194697: dataIn1 = 32'd716
; 
32'd194698: dataIn1 = 32'd1386
; 
32'd194699: dataIn1 = 32'd11242
; 
32'd194700: dataIn1 = 32'd11243
; 
32'd194701: dataIn1 = 32'd11244
; 
32'd194702: dataIn1 = 32'd1386
; 
32'd194703: dataIn1 = 32'd11243
; 
32'd194704: dataIn1 = 32'd11244
; 
32'd194705: dataIn1 = 32'd11245
; 
32'd194706: dataIn1 = 32'd717
; 
32'd194707: dataIn1 = 32'd1386
; 
32'd194708: dataIn1 = 32'd11244
; 
32'd194709: dataIn1 = 32'd11245
; 
32'd194710: dataIn1 = 32'd11246
; 
32'd194711: dataIn1 = 32'd717
; 
32'd194712: dataIn1 = 32'd11245
; 
32'd194713: dataIn1 = 32'd11246
; 
32'd194714: dataIn1 = 32'd11247
; 
32'd194715: dataIn1 = 32'd717
; 
32'd194716: dataIn1 = 32'd1388
; 
32'd194717: dataIn1 = 32'd11246
; 
32'd194718: dataIn1 = 32'd11247
; 
32'd194719: dataIn1 = 32'd11248
; 
32'd194720: dataIn1 = 32'd1388
; 
32'd194721: dataIn1 = 32'd11247
; 
32'd194722: dataIn1 = 32'd11248
; 
32'd194723: dataIn1 = 32'd11249
; 
32'd194724: dataIn1 = 32'd1388
; 
32'd194725: dataIn1 = 32'd11248
; 
32'd194726: dataIn1 = 32'd11249
; 
32'd194727: dataIn1 = 32'd11250
; 
32'd194728: dataIn1 = 32'd704
; 
32'd194729: dataIn1 = 32'd1388
; 
32'd194730: dataIn1 = 32'd11249
; 
32'd194731: dataIn1 = 32'd11250
; 
32'd194732: dataIn1 = 32'd11251
; 
32'd194733: dataIn1 = 32'd704
; 
32'd194734: dataIn1 = 32'd1379
; 
32'd194735: dataIn1 = 32'd11250
; 
32'd194736: dataIn1 = 32'd11251
; 
32'd194737: dataIn1 = 32'd11252
; 
32'd194738: dataIn1 = 32'd1379
; 
32'd194739: dataIn1 = 32'd11251
; 
32'd194740: dataIn1 = 32'd11252
; 
32'd194741: dataIn1 = 32'd11253
; 
32'd194742: dataIn1 = 32'd1379
; 
32'd194743: dataIn1 = 32'd11252
; 
32'd194744: dataIn1 = 32'd11253
; 
32'd194745: dataIn1 = 32'd11254
; 
32'd194746: dataIn1 = 32'd703
; 
32'd194747: dataIn1 = 32'd1379
; 
32'd194748: dataIn1 = 32'd11253
; 
32'd194749: dataIn1 = 32'd11254
; 
32'd194750: dataIn1 = 32'd11255
; 
32'd194751: dataIn1 = 32'd703
; 
32'd194752: dataIn1 = 32'd11254
; 
32'd194753: dataIn1 = 32'd11255
; 
32'd194754: dataIn1 = 32'd11256
; 
32'd194755: dataIn1 = 32'd703
; 
32'd194756: dataIn1 = 32'd1378
; 
32'd194757: dataIn1 = 32'd11255
; 
32'd194758: dataIn1 = 32'd11256
; 
32'd194759: dataIn1 = 32'd11257
; 
32'd194760: dataIn1 = 32'd1378
; 
32'd194761: dataIn1 = 32'd11256
; 
32'd194762: dataIn1 = 32'd11257
; 
32'd194763: dataIn1 = 32'd11258
; 
32'd194764: dataIn1 = 32'd701
; 
32'd194765: dataIn1 = 32'd1378
; 
32'd194766: dataIn1 = 32'd11257
; 
32'd194767: dataIn1 = 32'd11258
; 
32'd194768: dataIn1 = 32'd11259
; 
32'd194769: dataIn1 = 32'd701
; 
32'd194770: dataIn1 = 32'd1376
; 
32'd194771: dataIn1 = 32'd11258
; 
32'd194772: dataIn1 = 32'd11259
; 
32'd194773: dataIn1 = 32'd11260
; 
32'd194774: dataIn1 = 32'd1376
; 
32'd194775: dataIn1 = 32'd11259
; 
32'd194776: dataIn1 = 32'd11260
; 
32'd194777: dataIn1 = 32'd11261
; 
32'd194778: dataIn1 = 32'd1376
; 
32'd194779: dataIn1 = 32'd11260
; 
32'd194780: dataIn1 = 32'd11261
; 
32'd194781: dataIn1 = 32'd11262
; 
32'd194782: dataIn1 = 32'd700
; 
32'd194783: dataIn1 = 32'd1376
; 
32'd194784: dataIn1 = 32'd11261
; 
32'd194785: dataIn1 = 32'd11262
; 
32'd194786: dataIn1 = 32'd11263
; 
32'd194787: dataIn1 = 32'd700
; 
32'd194788: dataIn1 = 32'd11262
; 
32'd194789: dataIn1 = 32'd11263
; 
32'd194790: dataIn1 = 32'd11264
; 
32'd194791: dataIn1 = 32'd700
; 
32'd194792: dataIn1 = 32'd1377
; 
32'd194793: dataIn1 = 32'd11263
; 
32'd194794: dataIn1 = 32'd11264
; 
32'd194795: dataIn1 = 32'd11265
; 
32'd194796: dataIn1 = 32'd702
; 
32'd194797: dataIn1 = 32'd1377
; 
32'd194798: dataIn1 = 32'd11264
; 
32'd194799: dataIn1 = 32'd11265
; 
32'd194800: dataIn1 = 32'd11266
; 
32'd194801: dataIn1 = 32'd702
; 
32'd194802: dataIn1 = 32'd11265
; 
32'd194803: dataIn1 = 32'd11266
; 
32'd194804: dataIn1 = 32'd11267
; 
32'd194805: dataIn1 = 32'd702
; 
32'd194806: dataIn1 = 32'd11266
; 
32'd194807: dataIn1 = 32'd11267
; 
32'd194808: dataIn1 = 32'd11268
; 
32'd194809: dataIn1 = 32'd702
; 
32'd194810: dataIn1 = 32'd1380
; 
32'd194811: dataIn1 = 32'd11267
; 
32'd194812: dataIn1 = 32'd11268
; 
32'd194813: dataIn1 = 32'd11269
; 
32'd194814: dataIn1 = 32'd1380
; 
32'd194815: dataIn1 = 32'd11268
; 
32'd194816: dataIn1 = 32'd11269
; 
32'd194817: dataIn1 = 32'd11270
; 
32'd194818: dataIn1 = 32'd698
; 
32'd194819: dataIn1 = 32'd1380
; 
32'd194820: dataIn1 = 32'd11269
; 
32'd194821: dataIn1 = 32'd11270
; 
32'd194822: dataIn1 = 32'd11271
; 
32'd194823: dataIn1 = 32'd698
; 
32'd194824: dataIn1 = 32'd1374
; 
32'd194825: dataIn1 = 32'd11270
; 
32'd194826: dataIn1 = 32'd11271
; 
32'd194827: dataIn1 = 32'd11272
; 
32'd194828: dataIn1 = 32'd1374
; 
32'd194829: dataIn1 = 32'd11271
; 
32'd194830: dataIn1 = 32'd11272
; 
32'd194831: dataIn1 = 32'd11273
; 
32'd194832: dataIn1 = 32'd1374
; 
32'd194833: dataIn1 = 32'd11272
; 
32'd194834: dataIn1 = 32'd11273
; 
32'd194835: dataIn1 = 32'd11274
; 
32'd194836: dataIn1 = 32'd696
; 
32'd194837: dataIn1 = 32'd1374
; 
32'd194838: dataIn1 = 32'd11273
; 
32'd194839: dataIn1 = 32'd11274
; 
32'd194840: dataIn1 = 32'd11275
; 
32'd194841: dataIn1 = 32'd696
; 
32'd194842: dataIn1 = 32'd1373
; 
32'd194843: dataIn1 = 32'd11274
; 
32'd194844: dataIn1 = 32'd11275
; 
32'd194845: dataIn1 = 32'd11276
; 
32'd194846: dataIn1 = 32'd1373
; 
32'd194847: dataIn1 = 32'd11275
; 
32'd194848: dataIn1 = 32'd11276
; 
32'd194849: dataIn1 = 32'd11277
; 
32'd194850: dataIn1 = 32'd1373
; 
32'd194851: dataIn1 = 32'd11276
; 
32'd194852: dataIn1 = 32'd11277
; 
32'd194853: dataIn1 = 32'd11278
; 
32'd194854: dataIn1 = 32'd697
; 
32'd194855: dataIn1 = 32'd1373
; 
32'd194856: dataIn1 = 32'd11277
; 
32'd194857: dataIn1 = 32'd11278
; 
32'd194858: dataIn1 = 32'd11279
; 
32'd194859: dataIn1 = 32'd697
; 
32'd194860: dataIn1 = 32'd1375
; 
32'd194861: dataIn1 = 32'd11278
; 
32'd194862: dataIn1 = 32'd11279
; 
32'd194863: dataIn1 = 32'd11280
; 
32'd194864: dataIn1 = 32'd1375
; 
32'd194865: dataIn1 = 32'd11279
; 
32'd194866: dataIn1 = 32'd11280
; 
32'd194867: dataIn1 = 32'd11281
; 
32'd194868: dataIn1 = 32'd1375
; 
32'd194869: dataIn1 = 32'd11280
; 
32'd194870: dataIn1 = 32'd11281
; 
32'd194871: dataIn1 = 32'd11282
; 
32'd194872: dataIn1 = 32'd688
; 
32'd194873: dataIn1 = 32'd1375
; 
32'd194874: dataIn1 = 32'd11281
; 
32'd194875: dataIn1 = 32'd11282
; 
32'd194876: dataIn1 = 32'd11283
; 
32'd194877: dataIn1 = 32'd688
; 
32'd194878: dataIn1 = 32'd1368
; 
32'd194879: dataIn1 = 32'd11282
; 
32'd194880: dataIn1 = 32'd11283
; 
32'd194881: dataIn1 = 32'd11284
; 
32'd194882: dataIn1 = 32'd1368
; 
32'd194883: dataIn1 = 32'd11283
; 
32'd194884: dataIn1 = 32'd11284
; 
32'd194885: dataIn1 = 32'd11285
; 
32'd194886: dataIn1 = 32'd687
; 
32'd194887: dataIn1 = 32'd1368
; 
32'd194888: dataIn1 = 32'd11284
; 
32'd194889: dataIn1 = 32'd11285
; 
32'd194890: dataIn1 = 32'd11286
; 
32'd194891: dataIn1 = 32'd687
; 
32'd194892: dataIn1 = 32'd11285
; 
32'd194893: dataIn1 = 32'd11286
; 
32'd194894: dataIn1 = 32'd11287
; 
32'd194895: dataIn1 = 32'd687
; 
32'd194896: dataIn1 = 32'd11286
; 
32'd194897: dataIn1 = 32'd11287
; 
32'd194898: dataIn1 = 32'd11288
; 
32'd194899: dataIn1 = 32'd687
; 
32'd194900: dataIn1 = 32'd1367
; 
32'd194901: dataIn1 = 32'd11287
; 
32'd194902: dataIn1 = 32'd11288
; 
32'd194903: dataIn1 = 32'd11289
; 
32'd194904: dataIn1 = 32'd1367
; 
32'd194905: dataIn1 = 32'd11288
; 
32'd194906: dataIn1 = 32'd11289
; 
32'd194907: dataIn1 = 32'd11290
; 
32'd194908: dataIn1 = 32'd685
; 
32'd194909: dataIn1 = 32'd1367
; 
32'd194910: dataIn1 = 32'd11289
; 
32'd194911: dataIn1 = 32'd11290
; 
32'd194912: dataIn1 = 32'd11291
; 
32'd194913: dataIn1 = 32'd685
; 
32'd194914: dataIn1 = 32'd1365
; 
32'd194915: dataIn1 = 32'd11290
; 
32'd194916: dataIn1 = 32'd11291
; 
32'd194917: dataIn1 = 32'd11292
; 
32'd194918: dataIn1 = 32'd1365
; 
32'd194919: dataIn1 = 32'd11291
; 
32'd194920: dataIn1 = 32'd11292
; 
32'd194921: dataIn1 = 32'd11293
; 
32'd194922: dataIn1 = 32'd683
; 
32'd194923: dataIn1 = 32'd1365
; 
32'd194924: dataIn1 = 32'd11292
; 
32'd194925: dataIn1 = 32'd11293
; 
32'd194926: dataIn1 = 32'd11294
; 
32'd194927: dataIn1 = 32'd683
; 
32'd194928: dataIn1 = 32'd11293
; 
32'd194929: dataIn1 = 32'd11294
; 
32'd194930: dataIn1 = 32'd11295
; 
32'd194931: dataIn1 = 32'd683
; 
32'd194932: dataIn1 = 32'd1366
; 
32'd194933: dataIn1 = 32'd11294
; 
32'd194934: dataIn1 = 32'd11295
; 
32'd194935: dataIn1 = 32'd11296
; 
32'd194936: dataIn1 = 32'd1366
; 
32'd194937: dataIn1 = 32'd11295
; 
32'd194938: dataIn1 = 32'd11296
; 
32'd194939: dataIn1 = 32'd11297
; 
32'd194940: dataIn1 = 32'd1366
; 
32'd194941: dataIn1 = 32'd11296
; 
32'd194942: dataIn1 = 32'd11297
; 
32'd194943: dataIn1 = 32'd11298
; 
32'd194944: dataIn1 = 32'd686
; 
32'd194945: dataIn1 = 32'd1366
; 
32'd194946: dataIn1 = 32'd11297
; 
32'd194947: dataIn1 = 32'd11298
; 
32'd194948: dataIn1 = 32'd11299
; 
32'd194949: dataIn1 = 32'd686
; 
32'd194950: dataIn1 = 32'd1369
; 
32'd194951: dataIn1 = 32'd11298
; 
32'd194952: dataIn1 = 32'd11299
; 
32'd194953: dataIn1 = 32'd11300
; 
32'd194954: dataIn1 = 32'd1369
; 
32'd194955: dataIn1 = 32'd11299
; 
32'd194956: dataIn1 = 32'd11300
; 
32'd194957: dataIn1 = 32'd11301
; 
32'd194958: dataIn1 = 32'd1369
; 
32'd194959: dataIn1 = 32'd11300
; 
32'd194960: dataIn1 = 32'd11301
; 
32'd194961: dataIn1 = 32'd11302
; 
32'd194962: dataIn1 = 32'd691
; 
32'd194963: dataIn1 = 32'd1369
; 
32'd194964: dataIn1 = 32'd11301
; 
32'd194965: dataIn1 = 32'd11302
; 
32'd194966: dataIn1 = 32'd11303
; 
32'd194967: dataIn1 = 32'd691
; 
32'd194968: dataIn1 = 32'd1371
; 
32'd194969: dataIn1 = 32'd11302
; 
32'd194970: dataIn1 = 32'd11303
; 
32'd194971: dataIn1 = 32'd11304
; 
32'd194972: dataIn1 = 32'd1371
; 
32'd194973: dataIn1 = 32'd11303
; 
32'd194974: dataIn1 = 32'd11304
; 
32'd194975: dataIn1 = 32'd11305
; 
32'd194976: dataIn1 = 32'd1371
; 
32'd194977: dataIn1 = 32'd11304
; 
32'd194978: dataIn1 = 32'd11305
; 
32'd194979: dataIn1 = 32'd11306
; 
32'd194980: dataIn1 = 32'd692
; 
32'd194981: dataIn1 = 32'd1371
; 
32'd194982: dataIn1 = 32'd11305
; 
32'd194983: dataIn1 = 32'd11306
; 
32'd194984: dataIn1 = 32'd11307
; 
32'd194985: dataIn1 = 32'd692
; 
32'd194986: dataIn1 = 32'd1370
; 
32'd194987: dataIn1 = 32'd11306
; 
32'd194988: dataIn1 = 32'd11307
; 
32'd194989: dataIn1 = 32'd11308
; 
32'd194990: dataIn1 = 32'd1370
; 
32'd194991: dataIn1 = 32'd11307
; 
32'd194992: dataIn1 = 32'd11308
; 
32'd194993: dataIn1 = 32'd11309
; 
32'd194994: dataIn1 = 32'd693
; 
32'd194995: dataIn1 = 32'd1370
; 
32'd194996: dataIn1 = 32'd11308
; 
32'd194997: dataIn1 = 32'd11309
; 
32'd194998: dataIn1 = 32'd11310
; 
32'd194999: dataIn1 = 32'd693
; 
32'd195000: dataIn1 = 32'd11309
; 
32'd195001: dataIn1 = 32'd11310
; 
32'd195002: dataIn1 = 32'd11311
; 
32'd195003: dataIn1 = 32'd693
; 
32'd195004: dataIn1 = 32'd1372
; 
32'd195005: dataIn1 = 32'd11310
; 
32'd195006: dataIn1 = 32'd11311
; 
32'd195007: dataIn1 = 32'd11312
; 
32'd195008: dataIn1 = 32'd1372
; 
32'd195009: dataIn1 = 32'd11311
; 
32'd195010: dataIn1 = 32'd11312
; 
32'd195011: dataIn1 = 32'd11313
; 
32'd195012: dataIn1 = 32'd680
; 
32'd195013: dataIn1 = 32'd1372
; 
32'd195014: dataIn1 = 32'd11312
; 
32'd195015: dataIn1 = 32'd11313
; 
32'd195016: dataIn1 = 32'd11314
; 
32'd195017: dataIn1 = 32'd680
; 
32'd195018: dataIn1 = 32'd11313
; 
32'd195019: dataIn1 = 32'd11314
; 
32'd195020: dataIn1 = 32'd11315
; 
32'd195021: dataIn1 = 32'd680
; 
32'd195022: dataIn1 = 32'd1363
; 
32'd195023: dataIn1 = 32'd11314
; 
32'd195024: dataIn1 = 32'd11315
; 
32'd195025: dataIn1 = 32'd11316
; 
32'd195026: dataIn1 = 32'd1363
; 
32'd195027: dataIn1 = 32'd11315
; 
32'd195028: dataIn1 = 32'd11316
; 
32'd195029: dataIn1 = 32'd11317
; 
32'd195030: dataIn1 = 32'd679
; 
32'd195031: dataIn1 = 32'd1363
; 
32'd195032: dataIn1 = 32'd11316
; 
32'd195033: dataIn1 = 32'd11317
; 
32'd195034: dataIn1 = 32'd11318
; 
32'd195035: dataIn1 = 32'd679
; 
32'd195036: dataIn1 = 32'd11317
; 
32'd195037: dataIn1 = 32'd11318
; 
32'd195038: dataIn1 = 32'd11319
; 
32'd195039: dataIn1 = 32'd679
; 
32'd195040: dataIn1 = 32'd1362
; 
32'd195041: dataIn1 = 32'd11318
; 
32'd195042: dataIn1 = 32'd11319
; 
32'd195043: dataIn1 = 32'd11320
; 
32'd195044: dataIn1 = 32'd1362
; 
32'd195045: dataIn1 = 32'd11319
; 
32'd195046: dataIn1 = 32'd11320
; 
32'd195047: dataIn1 = 32'd11321
; 
32'd195048: dataIn1 = 32'd1362
; 
32'd195049: dataIn1 = 32'd11320
; 
32'd195050: dataIn1 = 32'd11321
; 
32'd195051: dataIn1 = 32'd11322
; 
32'd195052: dataIn1 = 32'd677
; 
32'd195053: dataIn1 = 32'd1362
; 
32'd195054: dataIn1 = 32'd11321
; 
32'd195055: dataIn1 = 32'd11322
; 
32'd195056: dataIn1 = 32'd11323
; 
32'd195057: dataIn1 = 32'd677
; 
32'd195058: dataIn1 = 32'd1360
; 
32'd195059: dataIn1 = 32'd11322
; 
32'd195060: dataIn1 = 32'd11323
; 
32'd195061: dataIn1 = 32'd11324
; 
32'd195062: dataIn1 = 32'd1360
; 
32'd195063: dataIn1 = 32'd11323
; 
32'd195064: dataIn1 = 32'd11324
; 
32'd195065: dataIn1 = 32'd11325
; 
32'd195066: dataIn1 = 32'd1360
; 
32'd195067: dataIn1 = 32'd11324
; 
32'd195068: dataIn1 = 32'd11325
; 
32'd195069: dataIn1 = 32'd11326
; 
32'd195070: dataIn1 = 32'd676
; 
32'd195071: dataIn1 = 32'd1360
; 
32'd195072: dataIn1 = 32'd11325
; 
32'd195073: dataIn1 = 32'd11326
; 
32'd195074: dataIn1 = 32'd11327
; 
32'd195075: dataIn1 = 32'd676
; 
32'd195076: dataIn1 = 32'd1361
; 
32'd195077: dataIn1 = 32'd11326
; 
32'd195078: dataIn1 = 32'd11327
; 
32'd195079: dataIn1 = 32'd11328
; 
32'd195080: dataIn1 = 32'd1361
; 
32'd195081: dataIn1 = 32'd11327
; 
32'd195082: dataIn1 = 32'd11328
; 
32'd195083: dataIn1 = 32'd11329
; 
32'd195084: dataIn1 = 32'd1361
; 
32'd195085: dataIn1 = 32'd11328
; 
32'd195086: dataIn1 = 32'd11329
; 
32'd195087: dataIn1 = 32'd11330
; 
32'd195088: dataIn1 = 32'd678
; 
32'd195089: dataIn1 = 32'd1361
; 
32'd195090: dataIn1 = 32'd11329
; 
32'd195091: dataIn1 = 32'd11330
; 
32'd195092: dataIn1 = 32'd11331
; 
32'd195093: dataIn1 = 32'd678
; 
32'd195094: dataIn1 = 32'd11330
; 
32'd195095: dataIn1 = 32'd11331
; 
32'd195096: dataIn1 = 32'd11332
; 
32'd195097: dataIn1 = 32'd678
; 
32'd195098: dataIn1 = 32'd1364
; 
32'd195099: dataIn1 = 32'd11331
; 
32'd195100: dataIn1 = 32'd11332
; 
32'd195101: dataIn1 = 32'd11333
; 
32'd195102: dataIn1 = 32'd1364
; 
32'd195103: dataIn1 = 32'd11332
; 
32'd195104: dataIn1 = 32'd11333
; 
32'd195105: dataIn1 = 32'd11334
; 
32'd195106: dataIn1 = 32'd674
; 
32'd195107: dataIn1 = 32'd1364
; 
32'd195108: dataIn1 = 32'd11333
; 
32'd195109: dataIn1 = 32'd11334
; 
32'd195110: dataIn1 = 32'd11335
; 
32'd195111: dataIn1 = 32'd674
; 
32'd195112: dataIn1 = 32'd1358
; 
32'd195113: dataIn1 = 32'd11334
; 
32'd195114: dataIn1 = 32'd11335
; 
32'd195115: dataIn1 = 32'd11336
; 
32'd195116: dataIn1 = 32'd1358
; 
32'd195117: dataIn1 = 32'd11335
; 
32'd195118: dataIn1 = 32'd11336
; 
32'd195119: dataIn1 = 32'd11337
; 
32'd195120: dataIn1 = 32'd672
; 
32'd195121: dataIn1 = 32'd1358
; 
32'd195122: dataIn1 = 32'd11336
; 
32'd195123: dataIn1 = 32'd11337
; 
32'd195124: dataIn1 = 32'd11338
; 
32'd195125: dataIn1 = 32'd672
; 
32'd195126: dataIn1 = 32'd11337
; 
32'd195127: dataIn1 = 32'd11338
; 
32'd195128: dataIn1 = 32'd11339
; 
32'd195129: dataIn1 = 32'd672
; 
32'd195130: dataIn1 = 32'd11338
; 
32'd195131: dataIn1 = 32'd11339
; 
32'd195132: dataIn1 = 32'd11340
; 
32'd195133: dataIn1 = 32'd672
; 
32'd195134: dataIn1 = 32'd1357
; 
32'd195135: dataIn1 = 32'd11339
; 
32'd195136: dataIn1 = 32'd11340
; 
32'd195137: dataIn1 = 32'd11341
; 
32'd195138: dataIn1 = 32'd1357
; 
32'd195139: dataIn1 = 32'd11340
; 
32'd195140: dataIn1 = 32'd11341
; 
32'd195141: dataIn1 = 32'd11342
; 
32'd195142: dataIn1 = 32'd673
; 
32'd195143: dataIn1 = 32'd1357
; 
32'd195144: dataIn1 = 32'd11341
; 
32'd195145: dataIn1 = 32'd11342
; 
32'd195146: dataIn1 = 32'd11343
; 
32'd195147: dataIn1 = 32'd673
; 
32'd195148: dataIn1 = 32'd11342
; 
32'd195149: dataIn1 = 32'd11343
; 
32'd195150: dataIn1 = 32'd11344
; 
32'd195151: dataIn1 = 32'd673
; 
32'd195152: dataIn1 = 32'd1359
; 
32'd195153: dataIn1 = 32'd11343
; 
32'd195154: dataIn1 = 32'd11344
; 
32'd195155: dataIn1 = 32'd11345
; 
32'd195156: dataIn1 = 32'd1359
; 
32'd195157: dataIn1 = 32'd11344
; 
32'd195158: dataIn1 = 32'd11345
; 
32'd195159: dataIn1 = 32'd11346
; 
32'd195160: dataIn1 = 32'd664
; 
32'd195161: dataIn1 = 32'd1359
; 
32'd195162: dataIn1 = 32'd11345
; 
32'd195163: dataIn1 = 32'd11346
; 
32'd195164: dataIn1 = 32'd11347
; 
32'd195165: dataIn1 = 32'd664
; 
32'd195166: dataIn1 = 32'd1352
; 
32'd195167: dataIn1 = 32'd11346
; 
32'd195168: dataIn1 = 32'd11347
; 
32'd195169: dataIn1 = 32'd11348
; 
32'd195170: dataIn1 = 32'd1352
; 
32'd195171: dataIn1 = 32'd11347
; 
32'd195172: dataIn1 = 32'd11348
; 
32'd195173: dataIn1 = 32'd11349
; 
32'd195174: dataIn1 = 32'd1352
; 
32'd195175: dataIn1 = 32'd11348
; 
32'd195176: dataIn1 = 32'd11349
; 
32'd195177: dataIn1 = 32'd11350
; 
32'd195178: dataIn1 = 32'd663
; 
32'd195179: dataIn1 = 32'd1352
; 
32'd195180: dataIn1 = 32'd11349
; 
32'd195181: dataIn1 = 32'd11350
; 
32'd195182: dataIn1 = 32'd11351
; 
32'd195183: dataIn1 = 32'd663
; 
32'd195184: dataIn1 = 32'd1351
; 
32'd195185: dataIn1 = 32'd11350
; 
32'd195186: dataIn1 = 32'd11351
; 
32'd195187: dataIn1 = 32'd11352
; 
32'd195188: dataIn1 = 32'd1351
; 
32'd195189: dataIn1 = 32'd11351
; 
32'd195190: dataIn1 = 32'd11352
; 
32'd195191: dataIn1 = 32'd11353
; 
32'd195192: dataIn1 = 32'd1351
; 
32'd195193: dataIn1 = 32'd11352
; 
32'd195194: dataIn1 = 32'd11353
; 
32'd195195: dataIn1 = 32'd11354
; 
32'd195196: dataIn1 = 32'd661
; 
32'd195197: dataIn1 = 32'd1351
; 
32'd195198: dataIn1 = 32'd11353
; 
32'd195199: dataIn1 = 32'd11354
; 
32'd195200: dataIn1 = 32'd11355
; 
32'd195201: dataIn1 = 32'd661
; 
32'd195202: dataIn1 = 32'd1349
; 
32'd195203: dataIn1 = 32'd11354
; 
32'd195204: dataIn1 = 32'd11355
; 
32'd195205: dataIn1 = 32'd11356
; 
32'd195206: dataIn1 = 32'd1349
; 
32'd195207: dataIn1 = 32'd11355
; 
32'd195208: dataIn1 = 32'd11356
; 
32'd195209: dataIn1 = 32'd11357
; 
32'd195210: dataIn1 = 32'd659
; 
32'd195211: dataIn1 = 32'd1349
; 
32'd195212: dataIn1 = 32'd11356
; 
32'd195213: dataIn1 = 32'd11357
; 
32'd195214: dataIn1 = 32'd11358
; 
32'd195215: dataIn1 = 32'd659
; 
32'd195216: dataIn1 = 32'd11357
; 
32'd195217: dataIn1 = 32'd11358
; 
32'd195218: dataIn1 = 32'd11359
; 
32'd195219: dataIn1 = 32'd659
; 
32'd195220: dataIn1 = 32'd11358
; 
32'd195221: dataIn1 = 32'd11359
; 
32'd195222: dataIn1 = 32'd11360
; 
32'd195223: dataIn1 = 32'd659
; 
32'd195224: dataIn1 = 32'd1350
; 
32'd195225: dataIn1 = 32'd11359
; 
32'd195226: dataIn1 = 32'd11360
; 
32'd195227: dataIn1 = 32'd11361
; 
32'd195228: dataIn1 = 32'd1350
; 
32'd195229: dataIn1 = 32'd11360
; 
32'd195230: dataIn1 = 32'd11361
; 
32'd195231: dataIn1 = 32'd11362
; 
32'd195232: dataIn1 = 32'd662
; 
32'd195233: dataIn1 = 32'd1350
; 
32'd195234: dataIn1 = 32'd11361
; 
32'd195235: dataIn1 = 32'd11362
; 
32'd195236: dataIn1 = 32'd11363
; 
32'd195237: dataIn1 = 32'd662
; 
32'd195238: dataIn1 = 32'd11362
; 
32'd195239: dataIn1 = 32'd11363
; 
32'd195240: dataIn1 = 32'd11364
; 
32'd195241: dataIn1 = 32'd662
; 
32'd195242: dataIn1 = 32'd1353
; 
32'd195243: dataIn1 = 32'd11363
; 
32'd195244: dataIn1 = 32'd11364
; 
32'd195245: dataIn1 = 32'd11365
; 
32'd195246: dataIn1 = 32'd667
; 
32'd195247: dataIn1 = 32'd1353
; 
32'd195248: dataIn1 = 32'd11364
; 
32'd195249: dataIn1 = 32'd11365
; 
32'd195250: dataIn1 = 32'd11366
; 
32'd195251: dataIn1 = 32'd667
; 
32'd195252: dataIn1 = 32'd11365
; 
32'd195253: dataIn1 = 32'd11366
; 
32'd195254: dataIn1 = 32'd11367
; 
32'd195255: dataIn1 = 32'd667
; 
32'd195256: dataIn1 = 32'd1355
; 
32'd195257: dataIn1 = 32'd11366
; 
32'd195258: dataIn1 = 32'd11367
; 
32'd195259: dataIn1 = 32'd11368
; 
32'd195260: dataIn1 = 32'd1355
; 
32'd195261: dataIn1 = 32'd11367
; 
32'd195262: dataIn1 = 32'd11368
; 
32'd195263: dataIn1 = 32'd11369
; 
32'd195264: dataIn1 = 32'd1355
; 
32'd195265: dataIn1 = 32'd11368
; 
32'd195266: dataIn1 = 32'd11369
; 
32'd195267: dataIn1 = 32'd11370
; 
32'd195268: dataIn1 = 32'd668
; 
32'd195269: dataIn1 = 32'd1355
; 
32'd195270: dataIn1 = 32'd11369
; 
32'd195271: dataIn1 = 32'd11370
; 
32'd195272: dataIn1 = 32'd11371
; 
32'd195273: dataIn1 = 32'd668
; 
32'd195274: dataIn1 = 32'd1354
; 
32'd195275: dataIn1 = 32'd11370
; 
32'd195276: dataIn1 = 32'd11371
; 
32'd195277: dataIn1 = 32'd11372
; 
32'd195278: dataIn1 = 32'd1354
; 
32'd195279: dataIn1 = 32'd11371
; 
32'd195280: dataIn1 = 32'd11372
; 
32'd195281: dataIn1 = 32'd11373
; 
32'd195282: dataIn1 = 32'd1354
; 
32'd195283: dataIn1 = 32'd11372
; 
32'd195284: dataIn1 = 32'd11373
; 
32'd195285: dataIn1 = 32'd11374
; 
32'd195286: dataIn1 = 32'd669
; 
32'd195287: dataIn1 = 32'd1354
; 
32'd195288: dataIn1 = 32'd11373
; 
32'd195289: dataIn1 = 32'd11374
; 
32'd195290: dataIn1 = 32'd11375
; 
32'd195291: dataIn1 = 32'd669
; 
32'd195292: dataIn1 = 32'd1356
; 
32'd195293: dataIn1 = 32'd11374
; 
32'd195294: dataIn1 = 32'd11375
; 
32'd195295: dataIn1 = 32'd11376
; 
32'd195296: dataIn1 = 32'd1356
; 
32'd195297: dataIn1 = 32'd11375
; 
32'd195298: dataIn1 = 32'd11376
; 
32'd195299: dataIn1 = 32'd11377
; 
32'd195300: dataIn1 = 32'd1356
; 
32'd195301: dataIn1 = 32'd11376
; 
32'd195302: dataIn1 = 32'd11377
; 
32'd195303: dataIn1 = 32'd11378
; 
32'd195304: dataIn1 = 32'd656
; 
32'd195305: dataIn1 = 32'd1356
; 
32'd195306: dataIn1 = 32'd11377
; 
32'd195307: dataIn1 = 32'd11378
; 
32'd195308: dataIn1 = 32'd11379
; 
32'd195309: dataIn1 = 32'd656
; 
32'd195310: dataIn1 = 32'd11378
; 
32'd195311: dataIn1 = 32'd11379
; 
32'd195312: dataIn1 = 32'd11380
; 
32'd195313: dataIn1 = 32'd656
; 
32'd195314: dataIn1 = 32'd1347
; 
32'd195315: dataIn1 = 32'd11379
; 
32'd195316: dataIn1 = 32'd11380
; 
32'd195317: dataIn1 = 32'd11381
; 
32'd195318: dataIn1 = 32'd655
; 
32'd195319: dataIn1 = 32'd1347
; 
32'd195320: dataIn1 = 32'd11380
; 
32'd195321: dataIn1 = 32'd11381
; 
32'd195322: dataIn1 = 32'd11382
; 
32'd195323: dataIn1 = 32'd655
; 
32'd195324: dataIn1 = 32'd11381
; 
32'd195325: dataIn1 = 32'd11382
; 
32'd195326: dataIn1 = 32'd11383
; 
32'd195327: dataIn1 = 32'd655
; 
32'd195328: dataIn1 = 32'd11382
; 
32'd195329: dataIn1 = 32'd11383
; 
32'd195330: dataIn1 = 32'd11384
; 
32'd195331: dataIn1 = 32'd655
; 
32'd195332: dataIn1 = 32'd1346
; 
32'd195333: dataIn1 = 32'd11383
; 
32'd195334: dataIn1 = 32'd11384
; 
32'd195335: dataIn1 = 32'd11385
; 
32'd195336: dataIn1 = 32'd653
; 
32'd195337: dataIn1 = 32'd1346
; 
32'd195338: dataIn1 = 32'd11384
; 
32'd195339: dataIn1 = 32'd11385
; 
32'd195340: dataIn1 = 32'd11386
; 
32'd195341: dataIn1 = 32'd653
; 
32'd195342: dataIn1 = 32'd11385
; 
32'd195343: dataIn1 = 32'd11386
; 
32'd195344: dataIn1 = 32'd11387
; 
32'd195345: dataIn1 = 32'd653
; 
32'd195346: dataIn1 = 32'd1344
; 
32'd195347: dataIn1 = 32'd11386
; 
32'd195348: dataIn1 = 32'd11387
; 
32'd195349: dataIn1 = 32'd11388
; 
32'd195350: dataIn1 = 32'd1344
; 
32'd195351: dataIn1 = 32'd11387
; 
32'd195352: dataIn1 = 32'd11388
; 
32'd195353: dataIn1 = 32'd11389
; 
32'd195354: dataIn1 = 32'd652
; 
32'd195355: dataIn1 = 32'd1344
; 
32'd195356: dataIn1 = 32'd11388
; 
32'd195357: dataIn1 = 32'd11389
; 
32'd195358: dataIn1 = 32'd11390
; 
32'd195359: dataIn1 = 32'd652
; 
32'd195360: dataIn1 = 32'd11389
; 
32'd195361: dataIn1 = 32'd11390
; 
32'd195362: dataIn1 = 32'd11391
; 
32'd195363: dataIn1 = 32'd652
; 
32'd195364: dataIn1 = 32'd1345
; 
32'd195365: dataIn1 = 32'd11390
; 
32'd195366: dataIn1 = 32'd11391
; 
32'd195367: dataIn1 = 32'd11392
; 
32'd195368: dataIn1 = 32'd1345
; 
32'd195369: dataIn1 = 32'd11391
; 
32'd195370: dataIn1 = 32'd11392
; 
32'd195371: dataIn1 = 32'd11393
; 
32'd195372: dataIn1 = 32'd1345
; 
32'd195373: dataIn1 = 32'd11392
; 
32'd195374: dataIn1 = 32'd11393
; 
32'd195375: dataIn1 = 32'd11394
; 
32'd195376: dataIn1 = 32'd654
; 
32'd195377: dataIn1 = 32'd1345
; 
32'd195378: dataIn1 = 32'd11393
; 
32'd195379: dataIn1 = 32'd11394
; 
32'd195380: dataIn1 = 32'd11395
; 
32'd195381: dataIn1 = 32'd654
; 
32'd195382: dataIn1 = 32'd1348
; 
32'd195383: dataIn1 = 32'd11394
; 
32'd195384: dataIn1 = 32'd11395
; 
32'd195385: dataIn1 = 32'd11396
; 
32'd195386: dataIn1 = 32'd1348
; 
32'd195387: dataIn1 = 32'd11395
; 
32'd195388: dataIn1 = 32'd11396
; 
32'd195389: dataIn1 = 32'd11397
; 
32'd195390: dataIn1 = 32'd650
; 
32'd195391: dataIn1 = 32'd1348
; 
32'd195392: dataIn1 = 32'd11396
; 
32'd195393: dataIn1 = 32'd11397
; 
32'd195394: dataIn1 = 32'd11398
; 
32'd195395: dataIn1 = 32'd650
; 
32'd195396: dataIn1 = 32'd11397
; 
32'd195397: dataIn1 = 32'd11398
; 
32'd195398: dataIn1 = 32'd11399
; 
32'd195399: dataIn1 = 32'd650
; 
32'd195400: dataIn1 = 32'd11398
; 
32'd195401: dataIn1 = 32'd11399
; 
32'd195402: dataIn1 = 32'd11400
; 
32'd195403: dataIn1 = 32'd650
; 
32'd195404: dataIn1 = 32'd1342
; 
32'd195405: dataIn1 = 32'd11399
; 
32'd195406: dataIn1 = 32'd11400
; 
32'd195407: dataIn1 = 32'd11401
; 
32'd195408: dataIn1 = 32'd1342
; 
32'd195409: dataIn1 = 32'd11400
; 
32'd195410: dataIn1 = 32'd11401
; 
32'd195411: dataIn1 = 32'd11402
; 
32'd195412: dataIn1 = 32'd648
; 
32'd195413: dataIn1 = 32'd1342
; 
32'd195414: dataIn1 = 32'd11401
; 
32'd195415: dataIn1 = 32'd11402
; 
32'd195416: dataIn1 = 32'd11403
; 
32'd195417: dataIn1 = 32'd648
; 
32'd195418: dataIn1 = 32'd1341
; 
32'd195419: dataIn1 = 32'd11402
; 
32'd195420: dataIn1 = 32'd11403
; 
32'd195421: dataIn1 = 32'd11404
; 
32'd195422: dataIn1 = 32'd1341
; 
32'd195423: dataIn1 = 32'd11403
; 
32'd195424: dataIn1 = 32'd11404
; 
32'd195425: dataIn1 = 32'd11405
; 
32'd195426: dataIn1 = 32'd649
; 
32'd195427: dataIn1 = 32'd1341
; 
32'd195428: dataIn1 = 32'd11404
; 
32'd195429: dataIn1 = 32'd11405
; 
32'd195430: dataIn1 = 32'd11406
; 
32'd195431: dataIn1 = 32'd649
; 
32'd195432: dataIn1 = 32'd11405
; 
32'd195433: dataIn1 = 32'd11406
; 
32'd195434: dataIn1 = 32'd11407
; 
32'd195435: dataIn1 = 32'd649
; 
32'd195436: dataIn1 = 32'd1343
; 
32'd195437: dataIn1 = 32'd11406
; 
32'd195438: dataIn1 = 32'd11407
; 
32'd195439: dataIn1 = 32'd11408
; 
32'd195440: dataIn1 = 32'd1343
; 
32'd195441: dataIn1 = 32'd11407
; 
32'd195442: dataIn1 = 32'd11408
; 
32'd195443: dataIn1 = 32'd11409
; 
32'd195444: dataIn1 = 32'd640
; 
32'd195445: dataIn1 = 32'd1343
; 
32'd195446: dataIn1 = 32'd11408
; 
32'd195447: dataIn1 = 32'd11409
; 
32'd195448: dataIn1 = 32'd11410
; 
32'd195449: dataIn1 = 32'd640
; 
32'd195450: dataIn1 = 32'd11409
; 
32'd195451: dataIn1 = 32'd11410
; 
32'd195452: dataIn1 = 32'd11411
; 
32'd195453: dataIn1 = 32'd640
; 
32'd195454: dataIn1 = 32'd1336
; 
32'd195455: dataIn1 = 32'd11410
; 
32'd195456: dataIn1 = 32'd11411
; 
32'd195457: dataIn1 = 32'd11412
; 
32'd195458: dataIn1 = 32'd1336
; 
32'd195459: dataIn1 = 32'd11411
; 
32'd195460: dataIn1 = 32'd11412
; 
32'd195461: dataIn1 = 32'd11413
; 
32'd195462: dataIn1 = 32'd1336
; 
32'd195463: dataIn1 = 32'd11412
; 
32'd195464: dataIn1 = 32'd11413
; 
32'd195465: dataIn1 = 32'd11414
; 
32'd195466: dataIn1 = 32'd639
; 
32'd195467: dataIn1 = 32'd1336
; 
32'd195468: dataIn1 = 32'd11413
; 
32'd195469: dataIn1 = 32'd11414
; 
32'd195470: dataIn1 = 32'd11415
; 
32'd195471: dataIn1 = 32'd639
; 
32'd195472: dataIn1 = 32'd1335
; 
32'd195473: dataIn1 = 32'd11414
; 
32'd195474: dataIn1 = 32'd11415
; 
32'd195475: dataIn1 = 32'd11416
; 
32'd195476: dataIn1 = 32'd1335
; 
32'd195477: dataIn1 = 32'd11415
; 
32'd195478: dataIn1 = 32'd11416
; 
32'd195479: dataIn1 = 32'd11417
; 
32'd195480: dataIn1 = 32'd637
; 
32'd195481: dataIn1 = 32'd1335
; 
32'd195482: dataIn1 = 32'd11416
; 
32'd195483: dataIn1 = 32'd11417
; 
32'd195484: dataIn1 = 32'd11418
; 
32'd195485: dataIn1 = 32'd637
; 
32'd195486: dataIn1 = 32'd11417
; 
32'd195487: dataIn1 = 32'd11418
; 
32'd195488: dataIn1 = 32'd11419
; 
32'd195489: dataIn1 = 32'd637
; 
32'd195490: dataIn1 = 32'd1333
; 
32'd195491: dataIn1 = 32'd11418
; 
32'd195492: dataIn1 = 32'd11419
; 
32'd195493: dataIn1 = 32'd11420
; 
32'd195494: dataIn1 = 32'd1333
; 
32'd195495: dataIn1 = 32'd11419
; 
32'd195496: dataIn1 = 32'd11420
; 
32'd195497: dataIn1 = 32'd11421
; 
32'd195498: dataIn1 = 32'd635
; 
32'd195499: dataIn1 = 32'd1333
; 
32'd195500: dataIn1 = 32'd11420
; 
32'd195501: dataIn1 = 32'd11421
; 
32'd195502: dataIn1 = 32'd11422
; 
32'd195503: dataIn1 = 32'd635
; 
32'd195504: dataIn1 = 32'd11421
; 
32'd195505: dataIn1 = 32'd11422
; 
32'd195506: dataIn1 = 32'd11423
; 
32'd195507: dataIn1 = 32'd635
; 
32'd195508: dataIn1 = 32'd1334
; 
32'd195509: dataIn1 = 32'd11422
; 
32'd195510: dataIn1 = 32'd11423
; 
32'd195511: dataIn1 = 32'd11424
; 
32'd195512: dataIn1 = 32'd1334
; 
32'd195513: dataIn1 = 32'd11423
; 
32'd195514: dataIn1 = 32'd11424
; 
32'd195515: dataIn1 = 32'd11425
; 
32'd195516: dataIn1 = 32'd1334
; 
32'd195517: dataIn1 = 32'd11424
; 
32'd195518: dataIn1 = 32'd11425
; 
32'd195519: dataIn1 = 32'd11426
; 
32'd195520: dataIn1 = 32'd638
; 
32'd195521: dataIn1 = 32'd1334
; 
32'd195522: dataIn1 = 32'd11425
; 
32'd195523: dataIn1 = 32'd11426
; 
32'd195524: dataIn1 = 32'd11427
; 
32'd195525: dataIn1 = 32'd638
; 
32'd195526: dataIn1 = 32'd11426
; 
32'd195527: dataIn1 = 32'd11427
; 
32'd195528: dataIn1 = 32'd11428
; 
32'd195529: dataIn1 = 32'd638
; 
32'd195530: dataIn1 = 32'd1337
; 
32'd195531: dataIn1 = 32'd11427
; 
32'd195532: dataIn1 = 32'd11428
; 
32'd195533: dataIn1 = 32'd11429
; 
32'd195534: dataIn1 = 32'd1337
; 
32'd195535: dataIn1 = 32'd11428
; 
32'd195536: dataIn1 = 32'd11429
; 
32'd195537: dataIn1 = 32'd11430
; 
32'd195538: dataIn1 = 32'd643
; 
32'd195539: dataIn1 = 32'd1337
; 
32'd195540: dataIn1 = 32'd11429
; 
32'd195541: dataIn1 = 32'd11430
; 
32'd195542: dataIn1 = 32'd11431
; 
32'd195543: dataIn1 = 32'd643
; 
32'd195544: dataIn1 = 32'd1339
; 
32'd195545: dataIn1 = 32'd11430
; 
32'd195546: dataIn1 = 32'd11431
; 
32'd195547: dataIn1 = 32'd11432
; 
32'd195548: dataIn1 = 32'd1339
; 
32'd195549: dataIn1 = 32'd11431
; 
32'd195550: dataIn1 = 32'd11432
; 
32'd195551: dataIn1 = 32'd11433
; 
32'd195552: dataIn1 = 32'd1339
; 
32'd195553: dataIn1 = 32'd11432
; 
32'd195554: dataIn1 = 32'd11433
; 
32'd195555: dataIn1 = 32'd11434
; 
32'd195556: dataIn1 = 32'd644
; 
32'd195557: dataIn1 = 32'd1339
; 
32'd195558: dataIn1 = 32'd11433
; 
32'd195559: dataIn1 = 32'd11434
; 
32'd195560: dataIn1 = 32'd11435
; 
32'd195561: dataIn1 = 32'd644
; 
32'd195562: dataIn1 = 32'd11434
; 
32'd195563: dataIn1 = 32'd11435
; 
32'd195564: dataIn1 = 32'd11436
; 
32'd195565: dataIn1 = 32'd644
; 
32'd195566: dataIn1 = 32'd1338
; 
32'd195567: dataIn1 = 32'd11435
; 
32'd195568: dataIn1 = 32'd11436
; 
32'd195569: dataIn1 = 32'd11437
; 
32'd195570: dataIn1 = 32'd1338
; 
32'd195571: dataIn1 = 32'd11436
; 
32'd195572: dataIn1 = 32'd11437
; 
32'd195573: dataIn1 = 32'd11438
; 
32'd195574: dataIn1 = 32'd645
; 
32'd195575: dataIn1 = 32'd1338
; 
32'd195576: dataIn1 = 32'd11437
; 
32'd195577: dataIn1 = 32'd11438
; 
32'd195578: dataIn1 = 32'd11439
; 
32'd195579: dataIn1 = 32'd645
; 
32'd195580: dataIn1 = 32'd1340
; 
32'd195581: dataIn1 = 32'd11438
; 
32'd195582: dataIn1 = 32'd11439
; 
32'd195583: dataIn1 = 32'd11440
; 
32'd195584: dataIn1 = 32'd1340
; 
32'd195585: dataIn1 = 32'd11439
; 
32'd195586: dataIn1 = 32'd11440
; 
32'd195587: dataIn1 = 32'd11441
; 
32'd195588: dataIn1 = 32'd632
; 
32'd195589: dataIn1 = 32'd1340
; 
32'd195590: dataIn1 = 32'd11440
; 
32'd195591: dataIn1 = 32'd11441
; 
32'd195592: dataIn1 = 32'd11442
; 
32'd195593: dataIn1 = 32'd632
; 
32'd195594: dataIn1 = 32'd11441
; 
32'd195595: dataIn1 = 32'd11442
; 
32'd195596: dataIn1 = 32'd11443
; 
32'd195597: dataIn1 = 32'd632
; 
32'd195598: dataIn1 = 32'd1331
; 
32'd195599: dataIn1 = 32'd11442
; 
32'd195600: dataIn1 = 32'd11443
; 
32'd195601: dataIn1 = 32'd11444
; 
32'd195602: dataIn1 = 32'd1331
; 
32'd195603: dataIn1 = 32'd11443
; 
32'd195604: dataIn1 = 32'd11444
; 
32'd195605: dataIn1 = 32'd11445
; 
32'd195606: dataIn1 = 32'd631
; 
32'd195607: dataIn1 = 32'd1331
; 
32'd195608: dataIn1 = 32'd11444
; 
32'd195609: dataIn1 = 32'd11445
; 
32'd195610: dataIn1 = 32'd11446
; 
32'd195611: dataIn1 = 32'd631
; 
32'd195612: dataIn1 = 32'd11445
; 
32'd195613: dataIn1 = 32'd11446
; 
32'd195614: dataIn1 = 32'd11447
; 
32'd195615: dataIn1 = 32'd631
; 
32'd195616: dataIn1 = 32'd1330
; 
32'd195617: dataIn1 = 32'd11446
; 
32'd195618: dataIn1 = 32'd11447
; 
32'd195619: dataIn1 = 32'd11448
; 
32'd195620: dataIn1 = 32'd1330
; 
32'd195621: dataIn1 = 32'd11447
; 
32'd195622: dataIn1 = 32'd11448
; 
32'd195623: dataIn1 = 32'd11449
; 
32'd195624: dataIn1 = 32'd629
; 
32'd195625: dataIn1 = 32'd1330
; 
32'd195626: dataIn1 = 32'd11448
; 
32'd195627: dataIn1 = 32'd11449
; 
32'd195628: dataIn1 = 32'd11450
; 
32'd195629: dataIn1 = 32'd629
; 
32'd195630: dataIn1 = 32'd11449
; 
32'd195631: dataIn1 = 32'd11450
; 
32'd195632: dataIn1 = 32'd11451
; 
32'd195633: dataIn1 = 32'd629
; 
32'd195634: dataIn1 = 32'd1328
; 
32'd195635: dataIn1 = 32'd11450
; 
32'd195636: dataIn1 = 32'd11451
; 
32'd195637: dataIn1 = 32'd11452
; 
32'd195638: dataIn1 = 32'd1328
; 
32'd195639: dataIn1 = 32'd11451
; 
32'd195640: dataIn1 = 32'd11452
; 
32'd195641: dataIn1 = 32'd11453
; 
32'd195642: dataIn1 = 32'd628
; 
32'd195643: dataIn1 = 32'd1328
; 
32'd195644: dataIn1 = 32'd11452
; 
32'd195645: dataIn1 = 32'd11453
; 
32'd195646: dataIn1 = 32'd11454
; 
32'd195647: dataIn1 = 32'd628
; 
32'd195648: dataIn1 = 32'd11453
; 
32'd195649: dataIn1 = 32'd11454
; 
32'd195650: dataIn1 = 32'd11455
; 
32'd195651: dataIn1 = 32'd628
; 
32'd195652: dataIn1 = 32'd1329
; 
32'd195653: dataIn1 = 32'd11454
; 
32'd195654: dataIn1 = 32'd11455
; 
32'd195655: dataIn1 = 32'd11456
; 
32'd195656: dataIn1 = 32'd1329
; 
32'd195657: dataIn1 = 32'd11455
; 
32'd195658: dataIn1 = 32'd11456
; 
32'd195659: dataIn1 = 32'd11457
; 
32'd195660: dataIn1 = 32'd630
; 
32'd195661: dataIn1 = 32'd1329
; 
32'd195662: dataIn1 = 32'd11456
; 
32'd195663: dataIn1 = 32'd11457
; 
32'd195664: dataIn1 = 32'd11458
; 
32'd195665: dataIn1 = 32'd630
; 
32'd195666: dataIn1 = 32'd11457
; 
32'd195667: dataIn1 = 32'd11458
; 
32'd195668: dataIn1 = 32'd11459
; 
32'd195669: dataIn1 = 32'd630
; 
32'd195670: dataIn1 = 32'd1332
; 
32'd195671: dataIn1 = 32'd11458
; 
32'd195672: dataIn1 = 32'd11459
; 
32'd195673: dataIn1 = 32'd11460
; 
32'd195674: dataIn1 = 32'd1332
; 
32'd195675: dataIn1 = 32'd11459
; 
32'd195676: dataIn1 = 32'd11460
; 
32'd195677: dataIn1 = 32'd11461
; 
32'd195678: dataIn1 = 32'd626
; 
32'd195679: dataIn1 = 32'd1332
; 
32'd195680: dataIn1 = 32'd11460
; 
32'd195681: dataIn1 = 32'd11461
; 
32'd195682: dataIn1 = 32'd11462
; 
32'd195683: dataIn1 = 32'd626
; 
32'd195684: dataIn1 = 32'd11461
; 
32'd195685: dataIn1 = 32'd11462
; 
32'd195686: dataIn1 = 32'd11463
; 
32'd195687: dataIn1 = 32'd626
; 
32'd195688: dataIn1 = 32'd1326
; 
32'd195689: dataIn1 = 32'd11462
; 
32'd195690: dataIn1 = 32'd11463
; 
32'd195691: dataIn1 = 32'd11464
; 
32'd195692: dataIn1 = 32'd1326
; 
32'd195693: dataIn1 = 32'd11463
; 
32'd195694: dataIn1 = 32'd11464
; 
32'd195695: dataIn1 = 32'd11465
; 
32'd195696: dataIn1 = 32'd1326
; 
32'd195697: dataIn1 = 32'd11464
; 
32'd195698: dataIn1 = 32'd11465
; 
32'd195699: dataIn1 = 32'd11466
; 
32'd195700: dataIn1 = 32'd624
; 
32'd195701: dataIn1 = 32'd1326
; 
32'd195702: dataIn1 = 32'd11465
; 
32'd195703: dataIn1 = 32'd11466
; 
32'd195704: dataIn1 = 32'd11467
; 
32'd195705: dataIn1 = 32'd624
; 
32'd195706: dataIn1 = 32'd11466
; 
32'd195707: dataIn1 = 32'd11467
; 
32'd195708: dataIn1 = 32'd11468
; 
32'd195709: dataIn1 = 32'd624
; 
32'd195710: dataIn1 = 32'd1325
; 
32'd195711: dataIn1 = 32'd11467
; 
32'd195712: dataIn1 = 32'd11468
; 
32'd195713: dataIn1 = 32'd11469
; 
32'd195714: dataIn1 = 32'd1325
; 
32'd195715: dataIn1 = 32'd11468
; 
32'd195716: dataIn1 = 32'd11469
; 
32'd195717: dataIn1 = 32'd11470
; 
32'd195718: dataIn1 = 32'd625
; 
32'd195719: dataIn1 = 32'd1325
; 
32'd195720: dataIn1 = 32'd11469
; 
32'd195721: dataIn1 = 32'd11470
; 
32'd195722: dataIn1 = 32'd11471
; 
32'd195723: dataIn1 = 32'd625
; 
32'd195724: dataIn1 = 32'd11470
; 
32'd195725: dataIn1 = 32'd11471
; 
32'd195726: dataIn1 = 32'd11472
; 
32'd195727: dataIn1 = 32'd625
; 
32'd195728: dataIn1 = 32'd1327
; 
32'd195729: dataIn1 = 32'd11471
; 
32'd195730: dataIn1 = 32'd11472
; 
32'd195731: dataIn1 = 32'd11473
; 
32'd195732: dataIn1 = 32'd1327
; 
32'd195733: dataIn1 = 32'd11472
; 
32'd195734: dataIn1 = 32'd11473
; 
32'd195735: dataIn1 = 32'd11474
; 
32'd195736: dataIn1 = 32'd616
; 
32'd195737: dataIn1 = 32'd1327
; 
32'd195738: dataIn1 = 32'd11473
; 
32'd195739: dataIn1 = 32'd11474
; 
32'd195740: dataIn1 = 32'd11475
; 
32'd195741: dataIn1 = 32'd616
; 
32'd195742: dataIn1 = 32'd11474
; 
32'd195743: dataIn1 = 32'd11475
; 
32'd195744: dataIn1 = 32'd11476
; 
32'd195745: dataIn1 = 32'd616
; 
32'd195746: dataIn1 = 32'd1320
; 
32'd195747: dataIn1 = 32'd11475
; 
32'd195748: dataIn1 = 32'd11476
; 
32'd195749: dataIn1 = 32'd11477
; 
32'd195750: dataIn1 = 32'd1320
; 
32'd195751: dataIn1 = 32'd11476
; 
32'd195752: dataIn1 = 32'd11477
; 
32'd195753: dataIn1 = 32'd11478
; 
32'd195754: dataIn1 = 32'd615
; 
32'd195755: dataIn1 = 32'd1320
; 
32'd195756: dataIn1 = 32'd11477
; 
32'd195757: dataIn1 = 32'd11478
; 
32'd195758: dataIn1 = 32'd11479
; 
32'd195759: dataIn1 = 32'd615
; 
32'd195760: dataIn1 = 32'd11478
; 
32'd195761: dataIn1 = 32'd11479
; 
32'd195762: dataIn1 = 32'd11480
; 
32'd195763: dataIn1 = 32'd615
; 
32'd195764: dataIn1 = 32'd1319
; 
32'd195765: dataIn1 = 32'd11479
; 
32'd195766: dataIn1 = 32'd11480
; 
32'd195767: dataIn1 = 32'd11481
; 
32'd195768: dataIn1 = 32'd1319
; 
32'd195769: dataIn1 = 32'd11480
; 
32'd195770: dataIn1 = 32'd11481
; 
32'd195771: dataIn1 = 32'd11482
; 
32'd195772: dataIn1 = 32'd613
; 
32'd195773: dataIn1 = 32'd1319
; 
32'd195774: dataIn1 = 32'd11481
; 
32'd195775: dataIn1 = 32'd11482
; 
32'd195776: dataIn1 = 32'd11483
; 
32'd195777: dataIn1 = 32'd613
; 
32'd195778: dataIn1 = 32'd11482
; 
32'd195779: dataIn1 = 32'd11483
; 
32'd195780: dataIn1 = 32'd11484
; 
32'd195781: dataIn1 = 32'd613
; 
32'd195782: dataIn1 = 32'd1317
; 
32'd195783: dataIn1 = 32'd11483
; 
32'd195784: dataIn1 = 32'd11484
; 
32'd195785: dataIn1 = 32'd11485
; 
32'd195786: dataIn1 = 32'd1317
; 
32'd195787: dataIn1 = 32'd11484
; 
32'd195788: dataIn1 = 32'd11485
; 
32'd195789: dataIn1 = 32'd11486
; 
32'd195790: dataIn1 = 32'd611
; 
32'd195791: dataIn1 = 32'd1317
; 
32'd195792: dataIn1 = 32'd11485
; 
32'd195793: dataIn1 = 32'd11486
; 
32'd195794: dataIn1 = 32'd11487
; 
32'd195795: dataIn1 = 32'd611
; 
32'd195796: dataIn1 = 32'd11486
; 
32'd195797: dataIn1 = 32'd11487
; 
32'd195798: dataIn1 = 32'd11488
; 
32'd195799: dataIn1 = 32'd611
; 
32'd195800: dataIn1 = 32'd1318
; 
32'd195801: dataIn1 = 32'd11487
; 
32'd195802: dataIn1 = 32'd11488
; 
32'd195803: dataIn1 = 32'd11489
; 
32'd195804: dataIn1 = 32'd1318
; 
32'd195805: dataIn1 = 32'd11488
; 
32'd195806: dataIn1 = 32'd11489
; 
32'd195807: dataIn1 = 32'd11490
; 
32'd195808: dataIn1 = 32'd614
; 
32'd195809: dataIn1 = 32'd1318
; 
32'd195810: dataIn1 = 32'd11489
; 
32'd195811: dataIn1 = 32'd11490
; 
32'd195812: dataIn1 = 32'd11491
; 
32'd195813: dataIn1 = 32'd614
; 
32'd195814: dataIn1 = 32'd11490
; 
32'd195815: dataIn1 = 32'd11491
; 
32'd195816: dataIn1 = 32'd11492
; 
32'd195817: dataIn1 = 32'd614
; 
32'd195818: dataIn1 = 32'd1321
; 
32'd195819: dataIn1 = 32'd11491
; 
32'd195820: dataIn1 = 32'd11492
; 
32'd195821: dataIn1 = 32'd11493
; 
32'd195822: dataIn1 = 32'd1321
; 
32'd195823: dataIn1 = 32'd11492
; 
32'd195824: dataIn1 = 32'd11493
; 
32'd195825: dataIn1 = 32'd11494
; 
32'd195826: dataIn1 = 32'd619
; 
32'd195827: dataIn1 = 32'd1321
; 
32'd195828: dataIn1 = 32'd11493
; 
32'd195829: dataIn1 = 32'd11494
; 
32'd195830: dataIn1 = 32'd11495
; 
32'd195831: dataIn1 = 32'd619
; 
32'd195832: dataIn1 = 32'd11494
; 
32'd195833: dataIn1 = 32'd11495
; 
32'd195834: dataIn1 = 32'd11496
; 
32'd195835: dataIn1 = 32'd619
; 
32'd195836: dataIn1 = 32'd1323
; 
32'd195837: dataIn1 = 32'd11495
; 
32'd195838: dataIn1 = 32'd11496
; 
32'd195839: dataIn1 = 32'd11497
; 
32'd195840: dataIn1 = 32'd1323
; 
32'd195841: dataIn1 = 32'd11496
; 
32'd195842: dataIn1 = 32'd11497
; 
32'd195843: dataIn1 = 32'd11498
; 
32'd195844: dataIn1 = 32'd620
; 
32'd195845: dataIn1 = 32'd1323
; 
32'd195846: dataIn1 = 32'd11497
; 
32'd195847: dataIn1 = 32'd11498
; 
32'd195848: dataIn1 = 32'd11499
; 
32'd195849: dataIn1 = 32'd620
; 
32'd195850: dataIn1 = 32'd1322
; 
32'd195851: dataIn1 = 32'd11498
; 
32'd195852: dataIn1 = 32'd11499
; 
32'd195853: dataIn1 = 32'd11500
; 
32'd195854: dataIn1 = 32'd1322
; 
32'd195855: dataIn1 = 32'd11499
; 
32'd195856: dataIn1 = 32'd11500
; 
32'd195857: dataIn1 = 32'd11501
; 
32'd195858: dataIn1 = 32'd621
; 
32'd195859: dataIn1 = 32'd1322
; 
32'd195860: dataIn1 = 32'd11500
; 
32'd195861: dataIn1 = 32'd11501
; 
32'd195862: dataIn1 = 32'd11502
; 
32'd195863: dataIn1 = 32'd621
; 
32'd195864: dataIn1 = 32'd11501
; 
32'd195865: dataIn1 = 32'd11502
; 
32'd195866: dataIn1 = 32'd11503
; 
32'd195867: dataIn1 = 32'd621
; 
32'd195868: dataIn1 = 32'd1324
; 
32'd195869: dataIn1 = 32'd11502
; 
32'd195870: dataIn1 = 32'd11503
; 
32'd195871: dataIn1 = 32'd11504
; 
32'd195872: dataIn1 = 32'd1324
; 
32'd195873: dataIn1 = 32'd11503
; 
32'd195874: dataIn1 = 32'd11504
; 
32'd195875: dataIn1 = 32'd11505
; 
32'd195876: dataIn1 = 32'd608
; 
32'd195877: dataIn1 = 32'd1324
; 
32'd195878: dataIn1 = 32'd11504
; 
32'd195879: dataIn1 = 32'd11505
; 
32'd195880: dataIn1 = 32'd11506
; 
32'd195881: dataIn1 = 32'd608
; 
32'd195882: dataIn1 = 32'd11505
; 
32'd195883: dataIn1 = 32'd11506
; 
32'd195884: dataIn1 = 32'd11507
; 
32'd195885: dataIn1 = 32'd608
; 
32'd195886: dataIn1 = 32'd1315
; 
32'd195887: dataIn1 = 32'd11506
; 
32'd195888: dataIn1 = 32'd11507
; 
32'd195889: dataIn1 = 32'd11508
; 
32'd195890: dataIn1 = 32'd1315
; 
32'd195891: dataIn1 = 32'd11507
; 
32'd195892: dataIn1 = 32'd11508
; 
32'd195893: dataIn1 = 32'd11509
; 
32'd195894: dataIn1 = 32'd607
; 
32'd195895: dataIn1 = 32'd1315
; 
32'd195896: dataIn1 = 32'd11508
; 
32'd195897: dataIn1 = 32'd11509
; 
32'd195898: dataIn1 = 32'd11510
; 
32'd195899: dataIn1 = 32'd607
; 
32'd195900: dataIn1 = 32'd11509
; 
32'd195901: dataIn1 = 32'd11510
; 
32'd195902: dataIn1 = 32'd11511
; 
32'd195903: dataIn1 = 32'd607
; 
32'd195904: dataIn1 = 32'd1314
; 
32'd195905: dataIn1 = 32'd11510
; 
32'd195906: dataIn1 = 32'd11511
; 
32'd195907: dataIn1 = 32'd11512
; 
32'd195908: dataIn1 = 32'd1314
; 
32'd195909: dataIn1 = 32'd11511
; 
32'd195910: dataIn1 = 32'd11512
; 
32'd195911: dataIn1 = 32'd11513
; 
32'd195912: dataIn1 = 32'd605
; 
32'd195913: dataIn1 = 32'd1314
; 
32'd195914: dataIn1 = 32'd11512
; 
32'd195915: dataIn1 = 32'd11513
; 
32'd195916: dataIn1 = 32'd11514
; 
32'd195917: dataIn1 = 32'd605
; 
32'd195918: dataIn1 = 32'd11513
; 
32'd195919: dataIn1 = 32'd11514
; 
32'd195920: dataIn1 = 32'd11515
; 
32'd195921: dataIn1 = 32'd605
; 
32'd195922: dataIn1 = 32'd1312
; 
32'd195923: dataIn1 = 32'd11514
; 
32'd195924: dataIn1 = 32'd11515
; 
32'd195925: dataIn1 = 32'd11516
; 
32'd195926: dataIn1 = 32'd1312
; 
32'd195927: dataIn1 = 32'd11515
; 
32'd195928: dataIn1 = 32'd11516
; 
32'd195929: dataIn1 = 32'd11517
; 
32'd195930: dataIn1 = 32'd604
; 
32'd195931: dataIn1 = 32'd1312
; 
32'd195932: dataIn1 = 32'd11516
; 
32'd195933: dataIn1 = 32'd11517
; 
32'd195934: dataIn1 = 32'd11518
; 
32'd195935: dataIn1 = 32'd604
; 
32'd195936: dataIn1 = 32'd11517
; 
32'd195937: dataIn1 = 32'd11518
; 
32'd195938: dataIn1 = 32'd11519
; 
32'd195939: dataIn1 = 32'd604
; 
32'd195940: dataIn1 = 32'd1313
; 
32'd195941: dataIn1 = 32'd11518
; 
32'd195942: dataIn1 = 32'd11519
; 
32'd195943: dataIn1 = 32'd11520
; 
32'd195944: dataIn1 = 32'd1313
; 
32'd195945: dataIn1 = 32'd11519
; 
32'd195946: dataIn1 = 32'd11520
; 
32'd195947: dataIn1 = 32'd11521
; 
32'd195948: dataIn1 = 32'd606
; 
32'd195949: dataIn1 = 32'd1313
; 
32'd195950: dataIn1 = 32'd11520
; 
32'd195951: dataIn1 = 32'd11521
; 
32'd195952: dataIn1 = 32'd11522
; 
32'd195953: dataIn1 = 32'd606
; 
32'd195954: dataIn1 = 32'd11521
; 
32'd195955: dataIn1 = 32'd11522
; 
32'd195956: dataIn1 = 32'd11523
; 
32'd195957: dataIn1 = 32'd606
; 
32'd195958: dataIn1 = 32'd11522
; 
32'd195959: dataIn1 = 32'd11523
; 
32'd195960: dataIn1 = 32'd11524
; 
32'd195961: dataIn1 = 32'd606
; 
32'd195962: dataIn1 = 32'd1316
; 
32'd195963: dataIn1 = 32'd11523
; 
32'd195964: dataIn1 = 32'd11524
; 
32'd195965: dataIn1 = 32'd11525
; 
32'd195966: dataIn1 = 32'd1316
; 
32'd195967: dataIn1 = 32'd11524
; 
32'd195968: dataIn1 = 32'd11525
; 
32'd195969: dataIn1 = 32'd11526
; 
32'd195970: dataIn1 = 32'd602
; 
32'd195971: dataIn1 = 32'd1316
; 
32'd195972: dataIn1 = 32'd11525
; 
32'd195973: dataIn1 = 32'd11526
; 
32'd195974: dataIn1 = 32'd11527
; 
32'd195975: dataIn1 = 32'd602
; 
32'd195976: dataIn1 = 32'd11526
; 
32'd195977: dataIn1 = 32'd11527
; 
32'd195978: dataIn1 = 32'd11528
; 
32'd195979: dataIn1 = 32'd602
; 
32'd195980: dataIn1 = 32'd1310
; 
32'd195981: dataIn1 = 32'd11527
; 
32'd195982: dataIn1 = 32'd11528
; 
32'd195983: dataIn1 = 32'd11529
; 
32'd195984: dataIn1 = 32'd1310
; 
32'd195985: dataIn1 = 32'd11528
; 
32'd195986: dataIn1 = 32'd11529
; 
32'd195987: dataIn1 = 32'd11530
; 
32'd195988: dataIn1 = 32'd600
; 
32'd195989: dataIn1 = 32'd1310
; 
32'd195990: dataIn1 = 32'd11529
; 
32'd195991: dataIn1 = 32'd11530
; 
32'd195992: dataIn1 = 32'd11531
; 
32'd195993: dataIn1 = 32'd600
; 
32'd195994: dataIn1 = 32'd11530
; 
32'd195995: dataIn1 = 32'd11531
; 
32'd195996: dataIn1 = 32'd11532
; 
32'd195997: dataIn1 = 32'd600
; 
32'd195998: dataIn1 = 32'd1309
; 
32'd195999: dataIn1 = 32'd11531
; 
32'd196000: dataIn1 = 32'd11532
; 
32'd196001: dataIn1 = 32'd11533
; 
32'd196002: dataIn1 = 32'd1309
; 
32'd196003: dataIn1 = 32'd11532
; 
32'd196004: dataIn1 = 32'd11533
; 
32'd196005: dataIn1 = 32'd11534
; 
32'd196006: dataIn1 = 32'd601
; 
32'd196007: dataIn1 = 32'd1309
; 
32'd196008: dataIn1 = 32'd11533
; 
32'd196009: dataIn1 = 32'd11534
; 
32'd196010: dataIn1 = 32'd11535
; 
32'd196011: dataIn1 = 32'd601
; 
32'd196012: dataIn1 = 32'd11534
; 
32'd196013: dataIn1 = 32'd11535
; 
32'd196014: dataIn1 = 32'd11536
; 
32'd196015: dataIn1 = 32'd601
; 
32'd196016: dataIn1 = 32'd1311
; 
32'd196017: dataIn1 = 32'd11535
; 
32'd196018: dataIn1 = 32'd11536
; 
32'd196019: dataIn1 = 32'd11537
; 
32'd196020: dataIn1 = 32'd592
; 
32'd196021: dataIn1 = 32'd1311
; 
32'd196022: dataIn1 = 32'd11536
; 
32'd196023: dataIn1 = 32'd11537
; 
32'd196024: dataIn1 = 32'd11538
; 
32'd196025: dataIn1 = 32'd592
; 
32'd196026: dataIn1 = 32'd11537
; 
32'd196027: dataIn1 = 32'd11538
; 
32'd196028: dataIn1 = 32'd11539
; 
32'd196029: dataIn1 = 32'd592
; 
32'd196030: dataIn1 = 32'd1304
; 
32'd196031: dataIn1 = 32'd11538
; 
32'd196032: dataIn1 = 32'd11539
; 
32'd196033: dataIn1 = 32'd11540
; 
32'd196034: dataIn1 = 32'd1304
; 
32'd196035: dataIn1 = 32'd11539
; 
32'd196036: dataIn1 = 32'd11540
; 
32'd196037: dataIn1 = 32'd11541
; 
32'd196038: dataIn1 = 32'd1304
; 
32'd196039: dataIn1 = 32'd11540
; 
32'd196040: dataIn1 = 32'd11541
; 
32'd196041: dataIn1 = 32'd11542
; 
32'd196042: dataIn1 = 32'd591
; 
32'd196043: dataIn1 = 32'd1304
; 
32'd196044: dataIn1 = 32'd11541
; 
32'd196045: dataIn1 = 32'd11542
; 
32'd196046: dataIn1 = 32'd11543
; 
32'd196047: dataIn1 = 32'd591
; 
32'd196048: dataIn1 = 32'd11542
; 
32'd196049: dataIn1 = 32'd11543
; 
32'd196050: dataIn1 = 32'd11544
; 
32'd196051: dataIn1 = 32'd591
; 
32'd196052: dataIn1 = 32'd1303
; 
32'd196053: dataIn1 = 32'd11543
; 
32'd196054: dataIn1 = 32'd11544
; 
32'd196055: dataIn1 = 32'd11545
; 
32'd196056: dataIn1 = 32'd1303
; 
32'd196057: dataIn1 = 32'd11544
; 
32'd196058: dataIn1 = 32'd11545
; 
32'd196059: dataIn1 = 32'd11546
; 
32'd196060: dataIn1 = 32'd589
; 
32'd196061: dataIn1 = 32'd1303
; 
32'd196062: dataIn1 = 32'd11545
; 
32'd196063: dataIn1 = 32'd11546
; 
32'd196064: dataIn1 = 32'd11547
; 
32'd196065: dataIn1 = 32'd589
; 
32'd196066: dataIn1 = 32'd11546
; 
32'd196067: dataIn1 = 32'd11547
; 
32'd196068: dataIn1 = 32'd11548
; 
32'd196069: dataIn1 = 32'd589
; 
32'd196070: dataIn1 = 32'd1301
; 
32'd196071: dataIn1 = 32'd11547
; 
32'd196072: dataIn1 = 32'd11548
; 
32'd196073: dataIn1 = 32'd11549
; 
32'd196074: dataIn1 = 32'd587
; 
32'd196075: dataIn1 = 32'd1301
; 
32'd196076: dataIn1 = 32'd11548
; 
32'd196077: dataIn1 = 32'd11549
; 
32'd196078: dataIn1 = 32'd11550
; 
32'd196079: dataIn1 = 32'd587
; 
32'd196080: dataIn1 = 32'd11549
; 
32'd196081: dataIn1 = 32'd11550
; 
32'd196082: dataIn1 = 32'd11551
; 
32'd196083: dataIn1 = 32'd587
; 
32'd196084: dataIn1 = 32'd1302
; 
32'd196085: dataIn1 = 32'd11550
; 
32'd196086: dataIn1 = 32'd11551
; 
32'd196087: dataIn1 = 32'd11552
; 
32'd196088: dataIn1 = 32'd1302
; 
32'd196089: dataIn1 = 32'd11551
; 
32'd196090: dataIn1 = 32'd11552
; 
32'd196091: dataIn1 = 32'd11553
; 
32'd196092: dataIn1 = 32'd590
; 
32'd196093: dataIn1 = 32'd1302
; 
32'd196094: dataIn1 = 32'd11552
; 
32'd196095: dataIn1 = 32'd11553
; 
32'd196096: dataIn1 = 32'd11554
; 
32'd196097: dataIn1 = 32'd590
; 
32'd196098: dataIn1 = 32'd11553
; 
32'd196099: dataIn1 = 32'd11554
; 
32'd196100: dataIn1 = 32'd11555
; 
32'd196101: dataIn1 = 32'd590
; 
32'd196102: dataIn1 = 32'd11554
; 
32'd196103: dataIn1 = 32'd11555
; 
32'd196104: dataIn1 = 32'd11556
; 
32'd196105: dataIn1 = 32'd590
; 
32'd196106: dataIn1 = 32'd1305
; 
32'd196107: dataIn1 = 32'd11555
; 
32'd196108: dataIn1 = 32'd11556
; 
32'd196109: dataIn1 = 32'd11557
; 
32'd196110: dataIn1 = 32'd1305
; 
32'd196111: dataIn1 = 32'd11556
; 
32'd196112: dataIn1 = 32'd11557
; 
32'd196113: dataIn1 = 32'd11558
; 
32'd196114: dataIn1 = 32'd595
; 
32'd196115: dataIn1 = 32'd1305
; 
32'd196116: dataIn1 = 32'd11557
; 
32'd196117: dataIn1 = 32'd11558
; 
32'd196118: dataIn1 = 32'd11559
; 
32'd196119: dataIn1 = 32'd595
; 
32'd196120: dataIn1 = 32'd11558
; 
32'd196121: dataIn1 = 32'd11559
; 
32'd196122: dataIn1 = 32'd11560
; 
32'd196123: dataIn1 = 32'd595
; 
32'd196124: dataIn1 = 32'd1307
; 
32'd196125: dataIn1 = 32'd11559
; 
32'd196126: dataIn1 = 32'd11560
; 
32'd196127: dataIn1 = 32'd11561
; 
32'd196128: dataIn1 = 32'd1307
; 
32'd196129: dataIn1 = 32'd11560
; 
32'd196130: dataIn1 = 32'd11561
; 
32'd196131: dataIn1 = 32'd11562
; 
32'd196132: dataIn1 = 32'd596
; 
32'd196133: dataIn1 = 32'd1307
; 
32'd196134: dataIn1 = 32'd11561
; 
32'd196135: dataIn1 = 32'd11562
; 
32'd196136: dataIn1 = 32'd11563
; 
32'd196137: dataIn1 = 32'd596
; 
32'd196138: dataIn1 = 32'd11562
; 
32'd196139: dataIn1 = 32'd11563
; 
32'd196140: dataIn1 = 32'd11564
; 
32'd196141: dataIn1 = 32'd596
; 
32'd196142: dataIn1 = 32'd1306
; 
32'd196143: dataIn1 = 32'd11563
; 
32'd196144: dataIn1 = 32'd11564
; 
32'd196145: dataIn1 = 32'd11565
; 
32'd196146: dataIn1 = 32'd1306
; 
32'd196147: dataIn1 = 32'd11564
; 
32'd196148: dataIn1 = 32'd11565
; 
32'd196149: dataIn1 = 32'd11566
; 
32'd196150: dataIn1 = 32'd597
; 
32'd196151: dataIn1 = 32'd1306
; 
32'd196152: dataIn1 = 32'd11565
; 
32'd196153: dataIn1 = 32'd11566
; 
32'd196154: dataIn1 = 32'd11567
; 
32'd196155: dataIn1 = 32'd597
; 
32'd196156: dataIn1 = 32'd1308
; 
32'd196157: dataIn1 = 32'd11566
; 
32'd196158: dataIn1 = 32'd11567
; 
32'd196159: dataIn1 = 32'd11568
; 
32'd196160: dataIn1 = 32'd1308
; 
32'd196161: dataIn1 = 32'd11567
; 
32'd196162: dataIn1 = 32'd11568
; 
32'd196163: dataIn1 = 32'd11569
; 
32'd196164: dataIn1 = 32'd580
; 
32'd196165: dataIn1 = 32'd1308
; 
32'd196166: dataIn1 = 32'd11568
; 
32'd196167: dataIn1 = 32'd11569
; 
32'd196168: dataIn1 = 32'd11570
; 
32'd196169: dataIn1 = 32'd580
; 
32'd196170: dataIn1 = 32'd11569
; 
32'd196171: dataIn1 = 32'd11570
; 
32'd196172: dataIn1 = 32'd11571
; 
32'd196173: dataIn1 = 32'd580
; 
32'd196174: dataIn1 = 32'd1297
; 
32'd196175: dataIn1 = 32'd11570
; 
32'd196176: dataIn1 = 32'd11571
; 
32'd196177: dataIn1 = 32'd11572
; 
32'd196178: dataIn1 = 32'd1297
; 
32'd196179: dataIn1 = 32'd11571
; 
32'd196180: dataIn1 = 32'd11572
; 
32'd196181: dataIn1 = 32'd11573
; 
32'd196182: dataIn1 = 32'd579
; 
32'd196183: dataIn1 = 32'd1297
; 
32'd196184: dataIn1 = 32'd11572
; 
32'd196185: dataIn1 = 32'd11573
; 
32'd196186: dataIn1 = 32'd11574
; 
32'd196187: dataIn1 = 32'd579
; 
32'd196188: dataIn1 = 32'd11573
; 
32'd196189: dataIn1 = 32'd11574
; 
32'd196190: dataIn1 = 32'd11575
; 
32'd196191: dataIn1 = 32'd579
; 
32'd196192: dataIn1 = 32'd1296
; 
32'd196193: dataIn1 = 32'd11574
; 
32'd196194: dataIn1 = 32'd11575
; 
32'd196195: dataIn1 = 32'd11576
; 
32'd196196: dataIn1 = 32'd1296
; 
32'd196197: dataIn1 = 32'd11575
; 
32'd196198: dataIn1 = 32'd11576
; 
32'd196199: dataIn1 = 32'd11577
; 
32'd196200: dataIn1 = 32'd577
; 
32'd196201: dataIn1 = 32'd1296
; 
32'd196202: dataIn1 = 32'd11576
; 
32'd196203: dataIn1 = 32'd11577
; 
32'd196204: dataIn1 = 32'd11578
; 
32'd196205: dataIn1 = 32'd577
; 
32'd196206: dataIn1 = 32'd11577
; 
32'd196207: dataIn1 = 32'd11578
; 
32'd196208: dataIn1 = 32'd11579
; 
32'd196209: dataIn1 = 32'd577
; 
32'd196210: dataIn1 = 32'd1294
; 
32'd196211: dataIn1 = 32'd11578
; 
32'd196212: dataIn1 = 32'd11579
; 
32'd196213: dataIn1 = 32'd11580
; 
32'd196214: dataIn1 = 32'd1294
; 
32'd196215: dataIn1 = 32'd11579
; 
32'd196216: dataIn1 = 32'd11580
; 
32'd196217: dataIn1 = 32'd11581
; 
32'd196218: dataIn1 = 32'd576
; 
32'd196219: dataIn1 = 32'd1294
; 
32'd196220: dataIn1 = 32'd11580
; 
32'd196221: dataIn1 = 32'd11581
; 
32'd196222: dataIn1 = 32'd11582
; 
32'd196223: dataIn1 = 32'd576
; 
32'd196224: dataIn1 = 32'd11581
; 
32'd196225: dataIn1 = 32'd11582
; 
32'd196226: dataIn1 = 32'd11583
; 
32'd196227: dataIn1 = 32'd576
; 
32'd196228: dataIn1 = 32'd1295
; 
32'd196229: dataIn1 = 32'd11582
; 
32'd196230: dataIn1 = 32'd11583
; 
32'd196231: dataIn1 = 32'd11584
; 
32'd196232: dataIn1 = 32'd1295
; 
32'd196233: dataIn1 = 32'd11583
; 
32'd196234: dataIn1 = 32'd11584
; 
32'd196235: dataIn1 = 32'd11585
; 
32'd196236: dataIn1 = 32'd578
; 
32'd196237: dataIn1 = 32'd1295
; 
32'd196238: dataIn1 = 32'd11584
; 
32'd196239: dataIn1 = 32'd11585
; 
32'd196240: dataIn1 = 32'd11586
; 
32'd196241: dataIn1 = 32'd578
; 
32'd196242: dataIn1 = 32'd11585
; 
32'd196243: dataIn1 = 32'd11586
; 
32'd196244: dataIn1 = 32'd11587
; 
32'd196245: dataIn1 = 32'd578
; 
32'd196246: dataIn1 = 32'd1298
; 
32'd196247: dataIn1 = 32'd11586
; 
32'd196248: dataIn1 = 32'd11587
; 
32'd196249: dataIn1 = 32'd11588
; 
32'd196250: dataIn1 = 32'd1298
; 
32'd196251: dataIn1 = 32'd11587
; 
32'd196252: dataIn1 = 32'd11588
; 
32'd196253: dataIn1 = 32'd11589
; 
32'd196254: dataIn1 = 32'd574
; 
32'd196255: dataIn1 = 32'd1298
; 
32'd196256: dataIn1 = 32'd11588
; 
32'd196257: dataIn1 = 32'd11589
; 
32'd196258: dataIn1 = 32'd11590
; 
32'd196259: dataIn1 = 32'd574
; 
32'd196260: dataIn1 = 32'd11589
; 
32'd196261: dataIn1 = 32'd11590
; 
32'd196262: dataIn1 = 32'd11591
; 
32'd196263: dataIn1 = 32'd574
; 
32'd196264: dataIn1 = 32'd1293
; 
32'd196265: dataIn1 = 32'd11590
; 
32'd196266: dataIn1 = 32'd11591
; 
32'd196267: dataIn1 = 32'd11592
; 
32'd196268: dataIn1 = 32'd1293
; 
32'd196269: dataIn1 = 32'd11591
; 
32'd196270: dataIn1 = 32'd11592
; 
32'd196271: dataIn1 = 32'd11593
; 
32'd196272: dataIn1 = 32'd1293
; 
32'd196273: dataIn1 = 32'd11592
; 
32'd196274: dataIn1 = 32'd11593
; 
32'd196275: dataIn1 = 32'd11594
; 
32'd196276: dataIn1 = 32'd573
; 
32'd196277: dataIn1 = 32'd1293
; 
32'd196278: dataIn1 = 32'd11593
; 
32'd196279: dataIn1 = 32'd11594
; 
32'd196280: dataIn1 = 32'd11595
; 
32'd196281: dataIn1 = 32'd573
; 
32'd196282: dataIn1 = 32'd11594
; 
32'd196283: dataIn1 = 32'd11595
; 
32'd196284: dataIn1 = 32'd11596
; 
32'd196285: dataIn1 = 32'd573
; 
32'd196286: dataIn1 = 32'd1289
; 
32'd196287: dataIn1 = 32'd1290
; 
32'd196288: dataIn1 = 32'd11595
; 
32'd196289: dataIn1 = 32'd11596
; 
32'd196290: dataIn1 = 32'd11597
; 
32'd196291: dataIn1 = 32'd1289
; 
32'd196292: dataIn1 = 32'd11596
; 
32'd196293: dataIn1 = 32'd11597
; 
32'd196294: dataIn1 = 32'd11598
; 
32'd196295: dataIn1 = 32'd1289
; 
32'd196296: dataIn1 = 32'd1291
; 
32'd196297: dataIn1 = 32'd11597
; 
32'd196298: dataIn1 = 32'd11598
; 
32'd196299: dataIn1 = 32'd11599
; 
32'd196300: dataIn1 = 32'd1291
; 
32'd196301: dataIn1 = 32'd11598
; 
32'd196302: dataIn1 = 32'd11599
; 
32'd196303: dataIn1 = 32'd11600
; 
32'd196304: dataIn1 = 32'd273
; 
32'd196305: dataIn1 = 32'd1277
; 
32'd196306: dataIn1 = 32'd1291
; 
32'd196307: dataIn1 = 32'd11599
; 
32'd196308: dataIn1 = 32'd11600
; 
32'd196309: dataIn1 = 32'd11601
; 
32'd196310: dataIn1 = 32'd1277
; 
32'd196311: dataIn1 = 32'd11600
; 
32'd196312: dataIn1 = 32'd11601
; 
32'd196313: dataIn1 = 32'd11602
; 
32'd196314: dataIn1 = 32'd1275
; 
32'd196315: dataIn1 = 32'd1277
; 
32'd196316: dataIn1 = 32'd11601
; 
32'd196317: dataIn1 = 32'd11602
; 
32'd196318: dataIn1 = 32'd11603
; 
32'd196319: dataIn1 = 32'd1275
; 
32'd196320: dataIn1 = 32'd11602
; 
32'd196321: dataIn1 = 32'd11603
; 
32'd196322: dataIn1 = 32'd11604
; 
32'd196323: dataIn1 = 32'd1275
; 
32'd196324: dataIn1 = 32'd11603
; 
32'd196325: dataIn1 = 32'd11604
; 
32'd196326: dataIn1 = 32'd11605
; 
32'd196327: dataIn1 = 32'd562
; 
32'd196328: dataIn1 = 32'd1275
; 
32'd196329: dataIn1 = 32'd1276
; 
32'd196330: dataIn1 = 32'd11604
; 
32'd196331: dataIn1 = 32'd11605
; 
32'd196332: dataIn1 = 32'd11606
; 
32'd196333: dataIn1 = 32'd562
; 
32'd196334: dataIn1 = 32'd11605
; 
32'd196335: dataIn1 = 32'd11606
; 
32'd196336: dataIn1 = 32'd11607
; 
32'd196337: dataIn1 = 32'd562
; 
32'd196338: dataIn1 = 32'd1279
; 
32'd196339: dataIn1 = 32'd11606
; 
32'd196340: dataIn1 = 32'd11607
; 
32'd196341: dataIn1 = 32'd11608
; 
32'd196342: dataIn1 = 32'd1279
; 
32'd196343: dataIn1 = 32'd11607
; 
32'd196344: dataIn1 = 32'd11608
; 
32'd196345: dataIn1 = 32'd11609
; 
32'd196346: dataIn1 = 32'd1279
; 
32'd196347: dataIn1 = 32'd11608
; 
32'd196348: dataIn1 = 32'd11609
; 
32'd196349: dataIn1 = 32'd11610
; 
32'd196350: dataIn1 = 32'd563
; 
32'd196351: dataIn1 = 32'd1279
; 
32'd196352: dataIn1 = 32'd11609
; 
32'd196353: dataIn1 = 32'd11610
; 
32'd196354: dataIn1 = 32'd11611
; 
32'd196355: dataIn1 = 32'd563
; 
32'd196356: dataIn1 = 32'd11610
; 
32'd196357: dataIn1 = 32'd11611
; 
32'd196358: dataIn1 = 32'd11612
; 
32'd196359: dataIn1 = 32'd563
; 
32'd196360: dataIn1 = 32'd1285
; 
32'd196361: dataIn1 = 32'd11611
; 
32'd196362: dataIn1 = 32'd11612
; 
32'd196363: dataIn1 = 32'd11613
; 
32'd196364: dataIn1 = 32'd1285
; 
32'd196365: dataIn1 = 32'd11612
; 
32'd196366: dataIn1 = 32'd11613
; 
32'd196367: dataIn1 = 32'd11614
; 
32'd196368: dataIn1 = 32'd1282
; 
32'd196369: dataIn1 = 32'd1285
; 
32'd196370: dataIn1 = 32'd11613
; 
32'd196371: dataIn1 = 32'd11614
; 
32'd196372: dataIn1 = 32'd11615
; 
32'd196373: dataIn1 = 32'd1282
; 
32'd196374: dataIn1 = 32'd11614
; 
32'd196375: dataIn1 = 32'd11615
; 
32'd196376: dataIn1 = 32'd11616
; 
32'd196377: dataIn1 = 32'd1281
; 
32'd196378: dataIn1 = 32'd1282
; 
32'd196379: dataIn1 = 32'd11615
; 
32'd196380: dataIn1 = 32'd11616
; 
32'd196381: dataIn1 = 32'd11617
; 
32'd196382: dataIn1 = 32'd1281
; 
32'd196383: dataIn1 = 32'd11616
; 
32'd196384: dataIn1 = 32'd11617
; 
32'd196385: dataIn1 = 32'd11618
; 
32'd196386: dataIn1 = 32'd1280
; 
32'd196387: dataIn1 = 32'd1281
; 
32'd196388: dataIn1 = 32'd11617
; 
32'd196389: dataIn1 = 32'd11618
; 
32'd196390: dataIn1 = 32'd11619
; 
32'd196391: dataIn1 = 32'd564
; 
32'd196392: dataIn1 = 32'd1280
; 
32'd196393: dataIn1 = 32'd11618
; 
32'd196394: dataIn1 = 32'd11619
; 
32'd196395: dataIn1 = 32'd11620
; 
32'd196396: dataIn1 = 32'd564
; 
32'd196397: dataIn1 = 32'd11619
; 
32'd196398: dataIn1 = 32'd11620
; 
32'd196399: dataIn1 = 32'd11621
; 
32'd196400: dataIn1 = 32'd564
; 
32'd196401: dataIn1 = 32'd1283
; 
32'd196402: dataIn1 = 32'd1284
; 
32'd196403: dataIn1 = 32'd11620
; 
32'd196404: dataIn1 = 32'd11621
; 
32'd196405: dataIn1 = 32'd11622
; 
32'd196406: dataIn1 = 32'd1284
; 
32'd196407: dataIn1 = 32'd11621
; 
32'd196408: dataIn1 = 32'd11622
; 
32'd196409: dataIn1 = 32'd11623
; 
32'd196410: dataIn1 = 32'd1284
; 
32'd196411: dataIn1 = 32'd1288
; 
32'd196412: dataIn1 = 32'd11622
; 
32'd196413: dataIn1 = 32'd11623
; 
32'd196414: dataIn1 = 32'd11624
; 
32'd196415: dataIn1 = 32'd570
; 
32'd196416: dataIn1 = 32'd1286
; 
32'd196417: dataIn1 = 32'd1288
; 
32'd196418: dataIn1 = 32'd11623
; 
32'd196419: dataIn1 = 32'd11624
; 
32'd196420: dataIn1 = 32'd11625
; 
32'd196421: dataIn1 = 32'd568
; 
32'd196422: dataIn1 = 32'd1286
; 
32'd196423: dataIn1 = 32'd11624
; 
32'd196424: dataIn1 = 32'd11625
; 
32'd196425: dataIn1 = 32'd11626
; 
32'd196426: dataIn1 = 32'd568
; 
32'd196427: dataIn1 = 32'd11625
; 
32'd196428: dataIn1 = 32'd11626
; 
32'd196429: dataIn1 = 32'd11627
; 
32'd196430: dataIn1 = 32'd568
; 
32'd196431: dataIn1 = 32'd1287
; 
32'd196432: dataIn1 = 32'd11626
; 
32'd196433: dataIn1 = 32'd11627
; 
32'd196434: dataIn1 = 32'd11628
; 
32'd196435: dataIn1 = 32'd1287
; 
32'd196436: dataIn1 = 32'd11627
; 
32'd196437: dataIn1 = 32'd11628
; 
32'd196438: dataIn1 = 32'd11629
; 
32'd196439: dataIn1 = 32'd560
; 
32'd196440: dataIn1 = 32'd1287
; 
32'd196441: dataIn1 = 32'd11628
; 
32'd196442: dataIn1 = 32'd11629
; 
32'd196443: dataIn1 = 32'd11630
; 
32'd196444: dataIn1 = 32'd560
; 
32'd196445: dataIn1 = 32'd11629
; 
32'd196446: dataIn1 = 32'd11630
; 
32'd196447: dataIn1 = 32'd11631
; 
32'd196448: dataIn1 = 32'd560
; 
32'd196449: dataIn1 = 32'd1274
; 
32'd196450: dataIn1 = 32'd11630
; 
32'd196451: dataIn1 = 32'd11631
; 
32'd196452: dataIn1 = 32'd11632
; 
32'd196453: dataIn1 = 32'd1274
; 
32'd196454: dataIn1 = 32'd11631
; 
32'd196455: dataIn1 = 32'd11632
; 
32'd196456: dataIn1 = 32'd11633
; 
32'd196457: dataIn1 = 32'd554
; 
32'd196458: dataIn1 = 32'd1274
; 
32'd196459: dataIn1 = 32'd11632
; 
32'd196460: dataIn1 = 32'd11633
; 
32'd196461: dataIn1 = 32'd11634
; 
32'd196462: dataIn1 = 32'd554
; 
32'd196463: dataIn1 = 32'd11633
; 
32'd196464: dataIn1 = 32'd11634
; 
32'd196465: dataIn1 = 32'd11635
; 
32'd196466: dataIn1 = 32'd554
; 
32'd196467: dataIn1 = 32'd1269
; 
32'd196468: dataIn1 = 32'd11634
; 
32'd196469: dataIn1 = 32'd11635
; 
32'd196470: dataIn1 = 32'd11636
; 
32'd196471: dataIn1 = 32'd1269
; 
32'd196472: dataIn1 = 32'd11635
; 
32'd196473: dataIn1 = 32'd11636
; 
32'd196474: dataIn1 = 32'd11637
; 
32'd196475: dataIn1 = 32'd1269
; 
32'd196476: dataIn1 = 32'd11636
; 
32'd196477: dataIn1 = 32'd11637
; 
32'd196478: dataIn1 = 32'd11638
; 
32'd196479: dataIn1 = 32'd551
; 
32'd196480: dataIn1 = 32'd1269
; 
32'd196481: dataIn1 = 32'd11637
; 
32'd196482: dataIn1 = 32'd11638
; 
32'd196483: dataIn1 = 32'd11639
; 
32'd196484: dataIn1 = 32'd551
; 
32'd196485: dataIn1 = 32'd11638
; 
32'd196486: dataIn1 = 32'd11639
; 
32'd196487: dataIn1 = 32'd11640
; 
32'd196488: dataIn1 = 32'd551
; 
32'd196489: dataIn1 = 32'd1268
; 
32'd196490: dataIn1 = 32'd11639
; 
32'd196491: dataIn1 = 32'd11640
; 
32'd196492: dataIn1 = 32'd11641
; 
32'd196493: dataIn1 = 32'd1268
; 
32'd196494: dataIn1 = 32'd11640
; 
32'd196495: dataIn1 = 32'd11641
; 
32'd196496: dataIn1 = 32'd11642
; 
32'd196497: dataIn1 = 32'd553
; 
32'd196498: dataIn1 = 32'd1268
; 
32'd196499: dataIn1 = 32'd11641
; 
32'd196500: dataIn1 = 32'd11642
; 
32'd196501: dataIn1 = 32'd11643
; 
32'd196502: dataIn1 = 32'd553
; 
32'd196503: dataIn1 = 32'd11642
; 
32'd196504: dataIn1 = 32'd11643
; 
32'd196505: dataIn1 = 32'd11644
; 
32'd196506: dataIn1 = 32'd553
; 
32'd196507: dataIn1 = 32'd1270
; 
32'd196508: dataIn1 = 32'd11643
; 
32'd196509: dataIn1 = 32'd11644
; 
32'd196510: dataIn1 = 32'd11645
; 
32'd196511: dataIn1 = 32'd555
; 
32'd196512: dataIn1 = 32'd1270
; 
32'd196513: dataIn1 = 32'd11644
; 
32'd196514: dataIn1 = 32'd11645
; 
32'd196515: dataIn1 = 32'd11646
; 
32'd196516: dataIn1 = 32'd555
; 
32'd196517: dataIn1 = 32'd11645
; 
32'd196518: dataIn1 = 32'd11646
; 
32'd196519: dataIn1 = 32'd11647
; 
32'd196520: dataIn1 = 32'd555
; 
32'd196521: dataIn1 = 32'd1273
; 
32'd196522: dataIn1 = 32'd11646
; 
32'd196523: dataIn1 = 32'd11647
; 
32'd196524: dataIn1 = 32'd11648
; 
32'd196525: dataIn1 = 32'd1273
; 
32'd196526: dataIn1 = 32'd11647
; 
32'd196527: dataIn1 = 32'd11648
; 
32'd196528: dataIn1 = 32'd11649
; 
32'd196529: dataIn1 = 32'd1273
; 
32'd196530: dataIn1 = 32'd11648
; 
32'd196531: dataIn1 = 32'd11649
; 
32'd196532: dataIn1 = 32'd11650
; 
32'd196533: dataIn1 = 32'd557
; 
32'd196534: dataIn1 = 32'd1273
; 
32'd196535: dataIn1 = 32'd11649
; 
32'd196536: dataIn1 = 32'd11650
; 
32'd196537: dataIn1 = 32'd11651
; 
32'd196538: dataIn1 = 32'd557
; 
32'd196539: dataIn1 = 32'd11650
; 
32'd196540: dataIn1 = 32'd11651
; 
32'd196541: dataIn1 = 32'd11652
; 
32'd196542: dataIn1 = 32'd557
; 
32'd196543: dataIn1 = 32'd11651
; 
32'd196544: dataIn1 = 32'd11652
; 
32'd196545: dataIn1 = 32'd11653
; 
32'd196546: dataIn1 = 32'd11654
; 
32'd196547: dataIn1 = 32'd11652
; 
32'd196548: dataIn1 = 32'd11653
; 
32'd196549: dataIn1 = 32'd11654
; 
32'd196550: dataIn1 = 32'd557
; 
32'd196551: dataIn1 = 32'd2101
; 
32'd196552: dataIn1 = 32'd11652
; 
32'd196553: dataIn1 = 32'd11653
; 
32'd196554: dataIn1 = 32'd11654
; 
32'd196555: dataIn1 = 32'd11655
; 
32'd196556: dataIn1 = 32'd2101
; 
32'd196557: dataIn1 = 32'd11654
; 
32'd196558: dataIn1 = 32'd11655
; 
32'd196559: dataIn1 = 32'd11656
; 
32'd196560: dataIn1 = 32'd2101
; 
32'd196561: dataIn1 = 32'd10247
; 
32'd196562: dataIn1 = 32'd11655
; 
32'd196563: dataIn1 = 32'd11656
; 
32'd196564: dataIn1 = 32'd11657
; 
32'd196565: dataIn1 = 32'd1272
; 
32'd196566: dataIn1 = 32'd10247
; 
32'd196567: dataIn1 = 32'd11656
; 
32'd196568: dataIn1 = 32'd11657
; 
32'd196569: dataIn1 = 32'd11658
; 
32'd196570: dataIn1 = 32'd1272
; 
32'd196571: dataIn1 = 32'd11657
; 
32'd196572: dataIn1 = 32'd11658
; 
32'd196573: dataIn1 = 32'd11659
; 
32'd196574: dataIn1 = 32'd556
; 
32'd196575: dataIn1 = 32'd1272
; 
32'd196576: dataIn1 = 32'd11658
; 
32'd196577: dataIn1 = 32'd11659
; 
32'd196578: dataIn1 = 32'd11660
; 
32'd196579: dataIn1 = 32'd556
; 
32'd196580: dataIn1 = 32'd1271
; 
32'd196581: dataIn1 = 32'd11659
; 
32'd196582: dataIn1 = 32'd11660
; 
32'd196583: dataIn1 = 32'd11661
; 
32'd196584: dataIn1 = 32'd1271
; 
32'd196585: dataIn1 = 32'd11660
; 
32'd196586: dataIn1 = 32'd11661
; 
32'd196587: dataIn1 = 32'd11662
; 
32'd196588: dataIn1 = 32'd1271
; 
32'd196589: dataIn1 = 32'd10564
; 
32'd196590: dataIn1 = 32'd11661
; 
32'd196591: dataIn1 = 32'd11662
; 
32'd196592: dataIn1 = 32'd11663
; 
32'd196593: dataIn1 = 32'd1488
; 
32'd196594: dataIn1 = 32'd10564
; 
32'd196595: dataIn1 = 32'd11662
; 
32'd196596: dataIn1 = 32'd11663
; 
32'd196597: dataIn1 = 32'd11664
; 
32'd196598: dataIn1 = 32'd1488
; 
32'd196599: dataIn1 = 32'd11663
; 
32'd196600: dataIn1 = 32'd11664
; 
32'd196601: dataIn1 = 32'd11665
; 
32'd196602: dataIn1 = 32'd782
; 
32'd196603: dataIn1 = 32'd1488
; 
32'd196604: dataIn1 = 32'd11664
; 
32'd196605: dataIn1 = 32'd11665
; 
32'd196606: dataIn1 = 32'd11666
; 
32'd196607: dataIn1 = 32'd782
; 
32'd196608: dataIn1 = 32'd1489
; 
32'd196609: dataIn1 = 32'd11665
; 
32'd196610: dataIn1 = 32'd11666
; 
32'd196611: dataIn1 = 32'd11667
; 
32'd196612: dataIn1 = 32'd1489
; 
32'd196613: dataIn1 = 32'd11666
; 
32'd196614: dataIn1 = 32'd11667
; 
32'd196615: dataIn1 = 32'd11668
; 
32'd196616: dataIn1 = 32'd1489
; 
32'd196617: dataIn1 = 32'd3439
; 
32'd196618: dataIn1 = 32'd11667
; 
32'd196619: dataIn1 = 32'd11668
; 
32'd196620: dataIn1 = 32'd11669
; 
32'd196621: dataIn1 = 32'd1462
; 
32'd196622: dataIn1 = 32'd3439
; 
32'd196623: dataIn1 = 32'd11668
; 
32'd196624: dataIn1 = 32'd11669
; 
32'd196625: dataIn1 = 32'd11670
; 
32'd196626: dataIn1 = 32'd1462
; 
32'd196627: dataIn1 = 32'd11669
; 
32'd196628: dataIn1 = 32'd11670
; 
32'd196629: dataIn1 = 32'd11671
; 
32'd196630: dataIn1 = 32'd1461
; 
32'd196631: dataIn1 = 32'd1462
; 
32'd196632: dataIn1 = 32'd11670
; 
32'd196633: dataIn1 = 32'd11671
; 
32'd196634: dataIn1 = 32'd11672
; 
32'd196635: dataIn1 = 32'd1461
; 
32'd196636: dataIn1 = 32'd10684
; 
32'd196637: dataIn1 = 32'd11671
; 
32'd196638: dataIn1 = 32'd11672
; 
32'd196639: dataIn1 = 32'd1170
; 
32'd196640: dataIn1 = 32'd1172
; 
32'd196641: dataIn1 = 32'd10565
; 
32'd196642: dataIn1 = 32'd11673
; 
32'd196643: dataIn1 = 32'd516
; 
32'd196644: dataIn1 = 32'd1174
; 
32'd196645: dataIn1 = 32'd10683
; 
32'd196646: dataIn1 = 32'd11674
; 
32'd196647: dataIn1 = 32'd11675
; 
32'd196648: dataIn1 = 32'd514
; 
32'd196649: dataIn1 = 32'd1174
; 
32'd196650: dataIn1 = 32'd11674
; 
32'd196651: dataIn1 = 32'd11675
; 
32'd196652: dataIn1 = 32'd11676
; 
32'd196653: dataIn1 = 32'd514
; 
32'd196654: dataIn1 = 32'd1168
; 
32'd196655: dataIn1 = 32'd11675
; 
32'd196656: dataIn1 = 32'd11676
; 
32'd196657: dataIn1 = 32'd11677
; 
32'd196658: dataIn1 = 32'd515
; 
32'd196659: dataIn1 = 32'd1168
; 
32'd196660: dataIn1 = 32'd1175
; 
32'd196661: dataIn1 = 32'd11676
; 
32'd196662: dataIn1 = 32'd11677
; 
32'd196663: dataIn1 = 32'd11678
; 
32'd196664: dataIn1 = 32'd508
; 
32'd196665: dataIn1 = 32'd1175
; 
32'd196666: dataIn1 = 32'd11677
; 
32'd196667: dataIn1 = 32'd11678
; 
32'd196668: dataIn1 = 32'd11679
; 
32'd196669: dataIn1 = 32'd508
; 
32'd196670: dataIn1 = 32'd1160
; 
32'd196671: dataIn1 = 32'd11678
; 
32'd196672: dataIn1 = 32'd11679
; 
32'd196673: dataIn1 = 32'd11680
; 
32'd196674: dataIn1 = 32'd509
; 
32'd196675: dataIn1 = 32'd1160
; 
32'd196676: dataIn1 = 32'd11679
; 
32'd196677: dataIn1 = 32'd11680
; 
32'd196678: dataIn1 = 32'd11681
; 
32'd196679: dataIn1 = 32'd509
; 
32'd196680: dataIn1 = 32'd1167
; 
32'd196681: dataIn1 = 32'd11680
; 
32'd196682: dataIn1 = 32'd11681
; 
32'd196683: dataIn1 = 32'd11682
; 
32'd196684: dataIn1 = 32'd512
; 
32'd196685: dataIn1 = 32'd1167
; 
32'd196686: dataIn1 = 32'd11681
; 
32'd196687: dataIn1 = 32'd11682
; 
32'd196688: dataIn1 = 32'd11683
; 
32'd196689: dataIn1 = 32'd512
; 
32'd196690: dataIn1 = 32'd1161
; 
32'd196691: dataIn1 = 32'd11682
; 
32'd196692: dataIn1 = 32'd11683
; 
32'd196693: dataIn1 = 32'd11684
; 
32'd196694: dataIn1 = 32'd510
; 
32'd196695: dataIn1 = 32'd1161
; 
32'd196696: dataIn1 = 32'd11683
; 
32'd196697: dataIn1 = 32'd11684
; 
32'd196698: dataIn1 = 32'd11685
; 
32'd196699: dataIn1 = 32'd510
; 
32'd196700: dataIn1 = 32'd1162
; 
32'd196701: dataIn1 = 32'd11684
; 
32'd196702: dataIn1 = 32'd11685
; 
32'd196703: dataIn1 = 32'd11686
; 
32'd196704: dataIn1 = 32'd505
; 
32'd196705: dataIn1 = 32'd1162
; 
32'd196706: dataIn1 = 32'd11685
; 
32'd196707: dataIn1 = 32'd11686
; 
32'd196708: dataIn1 = 32'd11687
; 
32'd196709: dataIn1 = 32'd505
; 
32'd196710: dataIn1 = 32'd1149
; 
32'd196711: dataIn1 = 32'd11686
; 
32'd196712: dataIn1 = 32'd11687
; 
32'd196713: dataIn1 = 32'd11688
; 
32'd196714: dataIn1 = 32'd506
; 
32'd196715: dataIn1 = 32'd1149
; 
32'd196716: dataIn1 = 32'd11687
; 
32'd196717: dataIn1 = 32'd11688
; 
32'd196718: dataIn1 = 32'd11689
; 
32'd196719: dataIn1 = 32'd506
; 
32'd196720: dataIn1 = 32'd1186
; 
32'd196721: dataIn1 = 32'd11688
; 
32'd196722: dataIn1 = 32'd11689
; 
32'd196723: dataIn1 = 32'd11690
; 
32'd196724: dataIn1 = 32'd520
; 
32'd196725: dataIn1 = 32'd1186
; 
32'd196726: dataIn1 = 32'd11689
; 
32'd196727: dataIn1 = 32'd11690
; 
32'd196728: dataIn1 = 32'd11691
; 
32'd196729: dataIn1 = 32'd520
; 
32'd196730: dataIn1 = 32'd1185
; 
32'd196731: dataIn1 = 32'd11690
; 
32'd196732: dataIn1 = 32'd11691
; 
32'd196733: dataIn1 = 32'd11692
; 
32'd196734: dataIn1 = 32'd521
; 
32'd196735: dataIn1 = 32'd1185
; 
32'd196736: dataIn1 = 32'd11691
; 
32'd196737: dataIn1 = 32'd11692
; 
32'd196738: dataIn1 = 32'd11693
; 
32'd196739: dataIn1 = 32'd521
; 
32'd196740: dataIn1 = 32'd1187
; 
32'd196741: dataIn1 = 32'd11692
; 
32'd196742: dataIn1 = 32'd11693
; 
32'd196743: dataIn1 = 32'd11694
; 
32'd196744: dataIn1 = 32'd519
; 
32'd196745: dataIn1 = 32'd1187
; 
32'd196746: dataIn1 = 32'd11693
; 
32'd196747: dataIn1 = 32'd11694
; 
32'd196748: dataIn1 = 32'd11695
; 
32'd196749: dataIn1 = 32'd519
; 
32'd196750: dataIn1 = 32'd11694
; 
32'd196751: dataIn1 = 32'd11695
; 
32'd196752: dataIn1 = 32'd11696
; 
32'd196753: dataIn1 = 32'd519
; 
32'd196754: dataIn1 = 32'd1183
; 
32'd196755: dataIn1 = 32'd11695
; 
32'd196756: dataIn1 = 32'd11696
; 
32'd196757: dataIn1 = 32'd11697
; 
32'd196758: dataIn1 = 32'd518
; 
32'd196759: dataIn1 = 32'd1183
; 
32'd196760: dataIn1 = 32'd11696
; 
32'd196761: dataIn1 = 32'd11697
; 
32'd196762: dataIn1 = 32'd11698
; 
32'd196763: dataIn1 = 32'd518
; 
32'd196764: dataIn1 = 32'd1198
; 
32'd196765: dataIn1 = 32'd11697
; 
32'd196766: dataIn1 = 32'd11698
; 
32'd196767: dataIn1 = 32'd11699
; 
32'd196768: dataIn1 = 32'd524
; 
32'd196769: dataIn1 = 32'd1198
; 
32'd196770: dataIn1 = 32'd11698
; 
32'd196771: dataIn1 = 32'd11699
; 
32'd196772: dataIn1 = 32'd11700
; 
32'd196773: dataIn1 = 32'd524
; 
32'd196774: dataIn1 = 32'd1192
; 
32'd196775: dataIn1 = 32'd11699
; 
32'd196776: dataIn1 = 32'd11700
; 
32'd196777: dataIn1 = 32'd11701
; 
32'd196778: dataIn1 = 32'd525
; 
32'd196779: dataIn1 = 32'd1192
; 
32'd196780: dataIn1 = 32'd11700
; 
32'd196781: dataIn1 = 32'd11701
; 
32'd196782: dataIn1 = 32'd11702
; 
32'd196783: dataIn1 = 32'd525
; 
32'd196784: dataIn1 = 32'd1199
; 
32'd196785: dataIn1 = 32'd11701
; 
32'd196786: dataIn1 = 32'd11702
; 
32'd196787: dataIn1 = 32'd11703
; 
32'd196788: dataIn1 = 32'd526
; 
32'd196789: dataIn1 = 32'd1199
; 
32'd196790: dataIn1 = 32'd11702
; 
32'd196791: dataIn1 = 32'd11703
; 
32'd196792: dataIn1 = 32'd11704
; 
32'd196793: dataIn1 = 32'd526
; 
32'd196794: dataIn1 = 32'd1206
; 
32'd196795: dataIn1 = 32'd11703
; 
32'd196796: dataIn1 = 32'd11704
; 
32'd196797: dataIn1 = 32'd11705
; 
32'd196798: dataIn1 = 32'd528
; 
32'd196799: dataIn1 = 32'd1206
; 
32'd196800: dataIn1 = 32'd11704
; 
32'd196801: dataIn1 = 32'd11705
; 
32'd196802: dataIn1 = 32'd11706
; 
32'd196803: dataIn1 = 32'd528
; 
32'd196804: dataIn1 = 32'd1238
; 
32'd196805: dataIn1 = 32'd11705
; 
32'd196806: dataIn1 = 32'd11706
; 
32'd196807: dataIn1 = 32'd11707
; 
32'd196808: dataIn1 = 32'd539
; 
32'd196809: dataIn1 = 32'd1238
; 
32'd196810: dataIn1 = 32'd11706
; 
32'd196811: dataIn1 = 32'd11707
; 
32'd196812: dataIn1 = 32'd11708
; 
32'd196813: dataIn1 = 32'd539
; 
32'd196814: dataIn1 = 32'd1233
; 
32'd196815: dataIn1 = 32'd11707
; 
32'd196816: dataIn1 = 32'd11708
; 
32'd196817: dataIn1 = 32'd11709
; 
32'd196818: dataIn1 = 32'd540
; 
32'd196819: dataIn1 = 32'd1233
; 
32'd196820: dataIn1 = 32'd11708
; 
32'd196821: dataIn1 = 32'd11709
; 
32'd196822: dataIn1 = 32'd11710
; 
32'd196823: dataIn1 = 32'd540
; 
32'd196824: dataIn1 = 32'd1239
; 
32'd196825: dataIn1 = 32'd11709
; 
32'd196826: dataIn1 = 32'd11710
; 
32'd196827: dataIn1 = 32'd11711
; 
32'd196828: dataIn1 = 32'd533
; 
32'd196829: dataIn1 = 32'd1239
; 
32'd196830: dataIn1 = 32'd11710
; 
32'd196831: dataIn1 = 32'd11711
; 
32'd196832: dataIn1 = 32'd11712
; 
32'd196833: dataIn1 = 32'd533
; 
32'd196834: dataIn1 = 32'd1225
; 
32'd196835: dataIn1 = 32'd11711
; 
32'd196836: dataIn1 = 32'd11712
; 
32'd196837: dataIn1 = 32'd11713
; 
32'd196838: dataIn1 = 32'd534
; 
32'd196839: dataIn1 = 32'd1225
; 
32'd196840: dataIn1 = 32'd11712
; 
32'd196841: dataIn1 = 32'd11713
; 
32'd196842: dataIn1 = 32'd11714
; 
32'd196843: dataIn1 = 32'd534
; 
32'd196844: dataIn1 = 32'd1232
; 
32'd196845: dataIn1 = 32'd11713
; 
32'd196846: dataIn1 = 32'd11714
; 
32'd196847: dataIn1 = 32'd11715
; 
32'd196848: dataIn1 = 32'd537
; 
32'd196849: dataIn1 = 32'd1232
; 
32'd196850: dataIn1 = 32'd11714
; 
32'd196851: dataIn1 = 32'd11715
; 
32'd196852: dataIn1 = 32'd11716
; 
32'd196853: dataIn1 = 32'd537
; 
32'd196854: dataIn1 = 32'd1226
; 
32'd196855: dataIn1 = 32'd11715
; 
32'd196856: dataIn1 = 32'd11716
; 
32'd196857: dataIn1 = 32'd11717
; 
32'd196858: dataIn1 = 32'd535
; 
32'd196859: dataIn1 = 32'd1226
; 
32'd196860: dataIn1 = 32'd11716
; 
32'd196861: dataIn1 = 32'd11717
; 
32'd196862: dataIn1 = 32'd11718
; 
32'd196863: dataIn1 = 32'd535
; 
32'd196864: dataIn1 = 32'd1227
; 
32'd196865: dataIn1 = 32'd11717
; 
32'd196866: dataIn1 = 32'd11718
; 
32'd196867: dataIn1 = 32'd11719
; 
32'd196868: dataIn1 = 32'd530
; 
32'd196869: dataIn1 = 32'd1227
; 
32'd196870: dataIn1 = 32'd11718
; 
32'd196871: dataIn1 = 32'd11719
; 
32'd196872: dataIn1 = 32'd11720
; 
32'd196873: dataIn1 = 32'd530
; 
32'd196874: dataIn1 = 32'd1214
; 
32'd196875: dataIn1 = 32'd11719
; 
32'd196876: dataIn1 = 32'd11720
; 
32'd196877: dataIn1 = 32'd11721
; 
32'd196878: dataIn1 = 32'd531
; 
32'd196879: dataIn1 = 32'd1214
; 
32'd196880: dataIn1 = 32'd11720
; 
32'd196881: dataIn1 = 32'd11721
; 
32'd196882: dataIn1 = 32'd11722
; 
32'd196883: dataIn1 = 32'd531
; 
32'd196884: dataIn1 = 32'd1252
; 
32'd196885: dataIn1 = 32'd11721
; 
32'd196886: dataIn1 = 32'd11722
; 
32'd196887: dataIn1 = 32'd11723
; 
32'd196888: dataIn1 = 32'd544
; 
32'd196889: dataIn1 = 32'd1252
; 
32'd196890: dataIn1 = 32'd11722
; 
32'd196891: dataIn1 = 32'd11723
; 
32'd196892: dataIn1 = 32'd11724
; 
32'd196893: dataIn1 = 32'd544
; 
32'd196894: dataIn1 = 32'd1251
; 
32'd196895: dataIn1 = 32'd11723
; 
32'd196896: dataIn1 = 32'd11724
; 
32'd196897: dataIn1 = 32'd11725
; 
32'd196898: dataIn1 = 32'd545
; 
32'd196899: dataIn1 = 32'd1251
; 
32'd196900: dataIn1 = 32'd11724
; 
32'd196901: dataIn1 = 32'd11725
; 
32'd196902: dataIn1 = 32'd11726
; 
32'd196903: dataIn1 = 32'd545
; 
32'd196904: dataIn1 = 32'd1253
; 
32'd196905: dataIn1 = 32'd11725
; 
32'd196906: dataIn1 = 32'd11726
; 
32'd196907: dataIn1 = 32'd11727
; 
32'd196908: dataIn1 = 32'd543
; 
32'd196909: dataIn1 = 32'd1247
; 
32'd196910: dataIn1 = 32'd1253
; 
32'd196911: dataIn1 = 32'd11726
; 
32'd196912: dataIn1 = 32'd11727
; 
32'd196913: dataIn1 = 32'd11728
; 
32'd196914: dataIn1 = 32'd1247
; 
32'd196915: dataIn1 = 32'd11727
; 
32'd196916: dataIn1 = 32'd11728
; 
32'd196917: dataIn1 = 32'd11729
; 
32'd196918: dataIn1 = 32'd1247
; 
32'd196919: dataIn1 = 32'd1249
; 
32'd196920: dataIn1 = 32'd11728
; 
32'd196921: dataIn1 = 32'd11729
; 
32'd196922: dataIn1 = 32'd11730
; 
32'd196923: dataIn1 = 32'd1249
; 
32'd196924: dataIn1 = 32'd1261
; 
32'd196925: dataIn1 = 32'd11729
; 
32'd196926: dataIn1 = 32'd11730
; 
32'd196927: dataIn1 = 32'd11731
; 
32'd196928: dataIn1 = 32'd1261
; 
32'd196929: dataIn1 = 32'd11730
; 
32'd196930: dataIn1 = 32'd11731
; 
32'd196931: dataIn1 = 32'd11732
; 
32'd196932: dataIn1 = 32'd744
; 
32'd196933: dataIn1 = 32'd1261
; 
32'd196934: dataIn1 = 32'd1432
; 
32'd196935: dataIn1 = 32'd11731
; 
32'd196936: dataIn1 = 32'd11732
; 
32'd196937: dataIn1 = 32'd11733
; 
32'd196938: dataIn1 = 32'd744
; 
32'd196939: dataIn1 = 32'd11732
; 
32'd196940: dataIn1 = 32'd11733
; 
32'd196941: dataIn1 = 32'd11734
; 
32'd196942: dataIn1 = 32'd744
; 
32'd196943: dataIn1 = 32'd1422
; 
32'd196944: dataIn1 = 32'd1423
; 
32'd196945: dataIn1 = 32'd11733
; 
32'd196946: dataIn1 = 32'd11734
; 
32'd196947: dataIn1 = 32'd11735
; 
32'd196948: dataIn1 = 32'd1422
; 
32'd196949: dataIn1 = 32'd11734
; 
32'd196950: dataIn1 = 32'd11735
; 
32'd196951: dataIn1 = 32'd11736
; 
32'd196952: dataIn1 = 32'd1421
; 
32'd196953: dataIn1 = 32'd1422
; 
32'd196954: dataIn1 = 32'd11735
; 
32'd196955: dataIn1 = 32'd11736
; 
32'd196956: dataIn1 = 32'd11737
; 
32'd196957: dataIn1 = 32'd743
; 
32'd196958: dataIn1 = 32'd1421
; 
32'd196959: dataIn1 = 32'd11736
; 
32'd196960: dataIn1 = 32'd11737
; 
32'd196961: dataIn1 = 32'd11738
; 
32'd196962: dataIn1 = 32'd743
; 
32'd196963: dataIn1 = 32'd10707
; 
32'd196964: dataIn1 = 32'd11737
; 
32'd196965: dataIn1 = 32'd11738
; 
default:  
	dataIn1 = 32'd99999; 
endcase 
case(addr2) 
32'd2: dataIn2 = 32'd1; 
32'd3: dataIn2 = 32'd1; 
32'd4: dataIn2 = 32'd1; 
32'd5: dataIn2 = 32'd1; 
32'd6: dataIn2 = 32'd0; 
32'd7: dataIn2 = 32'd0; 
32'd8: dataIn2 = 32'd1; 
32'd9: dataIn2 = 32'd1; 
32'd10: dataIn2 = 32'd1; 
32'd11: dataIn2 = 32'd0; 
32'd12: dataIn2 = 32'd1; 
32'd13: dataIn2 = 32'd0; 
32'd14: dataIn2 = 32'd1; 
32'd15: dataIn2 = 32'd1; 
32'd16: dataIn2 = 32'd1; 
32'd17: dataIn2 = 32'd0; 
32'd18: dataIn2 = 32'd0; 
32'd19: dataIn2 = 32'd1; 
32'd20: dataIn2 = 32'd0; 
32'd21: dataIn2 = 32'd1; 
32'd22: dataIn2 = 32'd0; 
32'd23: dataIn2 = 32'd0; 
32'd24: dataIn2 = 32'd1; 
32'd25: dataIn2 = 32'd0; 
32'd26: dataIn2 = 32'd1; 
32'd27: dataIn2 = 32'd1; 
32'd28: dataIn2 = 32'd1; 
32'd29: dataIn2 = 32'd0; 
32'd30: dataIn2 = 32'd0; 
32'd31: dataIn2 = 32'd0; 
32'd32: dataIn2 = 32'd0; 
32'd33: dataIn2 = 32'd0; 
32'd34: dataIn2 = 32'd0; 
32'd35: dataIn2 = 32'd0; 
32'd36: dataIn2 = 32'd1; 
32'd37: dataIn2 = 32'd1; 
32'd38: dataIn2 = 32'd1; 
32'd39: dataIn2 = 32'd0; 
32'd40: dataIn2 = 32'd1; 
32'd41: dataIn2 = 32'd0; 
32'd42: dataIn2 = 32'd0; 
32'd43: dataIn2 = 32'd1; 
32'd44: dataIn2 = 32'd0; 
32'd45: dataIn2 = 32'd1; 
32'd46: dataIn2 = 32'd0; 
32'd47: dataIn2 = 32'd0; 
32'd48: dataIn2 = 32'd0; 
32'd49: dataIn2 = 32'd0; 
32'd50: dataIn2 = 32'd0; 
32'd51: dataIn2 = 32'd0; 
32'd52: dataIn2 = 32'd0; 
32'd53: dataIn2 = 32'd0; 
32'd54: dataIn2 = 32'd1; 
32'd55: dataIn2 = 32'd0; 
32'd56: dataIn2 = 32'd0; 
32'd57: dataIn2 = 32'd0; 
32'd58: dataIn2 = 32'd1; 
32'd59: dataIn2 = 32'd1; 
32'd60: dataIn2 = 32'd0; 
32'd61: dataIn2 = 32'd0; 
32'd62: dataIn2 = 32'd0; 
32'd63: dataIn2 = 32'd1; 
32'd64: dataIn2 = 32'd0; 
32'd65: dataIn2 = 32'd0; 
32'd66: dataIn2 = 32'd1; 
32'd67: dataIn2 = 32'd1; 
32'd68: dataIn2 = 32'd0; 
32'd69: dataIn2 = 32'd1; 
32'd70: dataIn2 = 32'd1; 
32'd71: dataIn2 = 32'd1; 
32'd72: dataIn2 = 32'd1; 
32'd73: dataIn2 = 32'd0; 
32'd74: dataIn2 = 32'd1; 
32'd75: dataIn2 = 32'd1; 
32'd76: dataIn2 = 32'd1; 
32'd77: dataIn2 = 32'd1; 
32'd78: dataIn2 = 32'd1; 
32'd79: dataIn2 = 32'd0; 
32'd80: dataIn2 = 32'd0; 
32'd81: dataIn2 = 32'd0; 
32'd82: dataIn2 = 32'd0; 
32'd83: dataIn2 = 32'd1; 
32'd84: dataIn2 = 32'd1; 
32'd85: dataIn2 = 32'd0; 
32'd86: dataIn2 = 32'd0; 
32'd87: dataIn2 = 32'd1; 
32'd88: dataIn2 = 32'd0; 
32'd89: dataIn2 = 32'd0; 
32'd90: dataIn2 = 32'd0; 
32'd91: dataIn2 = 32'd1; 
32'd92: dataIn2 = 32'd1; 
32'd93: dataIn2 = 32'd0; 
32'd94: dataIn2 = 32'd1; 
32'd95: dataIn2 = 32'd1; 
32'd96: dataIn2 = 32'd0; 
32'd97: dataIn2 = 32'd1; 
32'd98: dataIn2 = 32'd0; 
32'd99: dataIn2 = 32'd0; 
32'd100: dataIn2 = 32'd1; 
32'd101: dataIn2 = 32'd0; 
32'd102: dataIn2 = 32'd0; 
32'd103: dataIn2 = 32'd0; 
32'd104: dataIn2 = 32'd1; 
32'd105: dataIn2 = 32'd1; 
32'd106: dataIn2 = 32'd0; 
32'd107: dataIn2 = 32'd1; 
32'd108: dataIn2 = 32'd0; 
32'd109: dataIn2 = 32'd1; 
32'd110: dataIn2 = 32'd0; 
32'd111: dataIn2 = 32'd0; 
32'd112: dataIn2 = 32'd1; 
32'd113: dataIn2 = 32'd0; 
32'd114: dataIn2 = 32'd1; 
32'd115: dataIn2 = 32'd0; 
32'd116: dataIn2 = 32'd1; 
32'd117: dataIn2 = 32'd0; 
32'd118: dataIn2 = 32'd1; 
32'd119: dataIn2 = 32'd1; 
32'd120: dataIn2 = 32'd0; 
32'd121: dataIn2 = 32'd1; 
32'd122: dataIn2 = 32'd1; 
32'd123: dataIn2 = 32'd0; 
32'd124: dataIn2 = 32'd1; 
32'd125: dataIn2 = 32'd1; 
32'd126: dataIn2 = 32'd1; 
32'd127: dataIn2 = 32'd0; 
32'd128: dataIn2 = 32'd0; 
32'd129: dataIn2 = 32'd0; 
32'd130: dataIn2 = 32'd1; 
32'd131: dataIn2 = 32'd0; 
32'd132: dataIn2 = 32'd0; 
32'd133: dataIn2 = 32'd0; 
32'd134: dataIn2 = 32'd0; 
32'd135: dataIn2 = 32'd1; 
32'd136: dataIn2 = 32'd1; 
32'd137: dataIn2 = 32'd0; 
32'd138: dataIn2 = 32'd1; 
32'd139: dataIn2 = 32'd1; 
32'd140: dataIn2 = 32'd1; 
32'd141: dataIn2 = 32'd0; 
32'd142: dataIn2 = 32'd1; 
32'd143: dataIn2 = 32'd0; 
32'd144: dataIn2 = 32'd0; 
32'd145: dataIn2 = 32'd1; 
32'd146: dataIn2 = 32'd1; 
32'd147: dataIn2 = 32'd1; 
32'd148: dataIn2 = 32'd0; 
32'd149: dataIn2 = 32'd0; 
32'd150: dataIn2 = 32'd1; 
32'd151: dataIn2 = 32'd0; 
32'd152: dataIn2 = 32'd0; 
32'd153: dataIn2 = 32'd0; 
32'd154: dataIn2 = 32'd0; 
32'd155: dataIn2 = 32'd1; 
32'd156: dataIn2 = 32'd0; 
32'd157: dataIn2 = 32'd0; 
32'd158: dataIn2 = 32'd1; 
32'd159: dataIn2 = 32'd0; 
32'd160: dataIn2 = 32'd0; 
32'd161: dataIn2 = 32'd0; 
32'd162: dataIn2 = 32'd1; 
32'd163: dataIn2 = 32'd0; 
32'd164: dataIn2 = 32'd0; 
32'd165: dataIn2 = 32'd0; 
32'd166: dataIn2 = 32'd0; 
32'd167: dataIn2 = 32'd0; 
32'd168: dataIn2 = 32'd1; 
32'd169: dataIn2 = 32'd0; 
32'd170: dataIn2 = 32'd0; 
32'd171: dataIn2 = 32'd0; 
32'd172: dataIn2 = 32'd0; 
32'd173: dataIn2 = 32'd1; 
32'd174: dataIn2 = 32'd1; 
32'd175: dataIn2 = 32'd0; 
32'd176: dataIn2 = 32'd1; 
32'd177: dataIn2 = 32'd0; 
32'd178: dataIn2 = 32'd1; 
32'd179: dataIn2 = 32'd0; 
32'd180: dataIn2 = 32'd0; 
32'd181: dataIn2 = 32'd1; 
32'd182: dataIn2 = 32'd0; 
32'd183: dataIn2 = 32'd1; 
32'd184: dataIn2 = 32'd1; 
32'd185: dataIn2 = 32'd0; 
32'd186: dataIn2 = 32'd1; 
32'd187: dataIn2 = 32'd1; 
32'd188: dataIn2 = 32'd1; 
32'd189: dataIn2 = 32'd1; 
32'd190: dataIn2 = 32'd1; 
32'd191: dataIn2 = 32'd1; 
32'd192: dataIn2 = 32'd1; 
32'd193: dataIn2 = 32'd0; 
32'd194: dataIn2 = 32'd1; 
32'd195: dataIn2 = 32'd0; 
32'd196: dataIn2 = 32'd1; 
32'd197: dataIn2 = 32'd0; 
32'd198: dataIn2 = 32'd0; 
32'd199: dataIn2 = 32'd1; 
32'd200: dataIn2 = 32'd0; 
32'd201: dataIn2 = 32'd1; 
32'd202: dataIn2 = 32'd0; 
32'd203: dataIn2 = 32'd0; 
32'd204: dataIn2 = 32'd0; 
32'd205: dataIn2 = 32'd0; 
32'd206: dataIn2 = 32'd1; 
32'd207: dataIn2 = 32'd0; 
32'd208: dataIn2 = 32'd0; 
32'd209: dataIn2 = 32'd0; 
32'd210: dataIn2 = 32'd0; 
32'd211: dataIn2 = 32'd1; 
32'd212: dataIn2 = 32'd1; 
32'd213: dataIn2 = 32'd1; 
32'd214: dataIn2 = 32'd0; 
32'd215: dataIn2 = 32'd1; 
32'd216: dataIn2 = 32'd0; 
32'd217: dataIn2 = 32'd0; 
32'd218: dataIn2 = 32'd0; 
32'd219: dataIn2 = 32'd1; 
32'd220: dataIn2 = 32'd0; 
32'd221: dataIn2 = 32'd1; 
32'd222: dataIn2 = 32'd1; 
32'd223: dataIn2 = 32'd1; 
32'd224: dataIn2 = 32'd1; 
32'd225: dataIn2 = 32'd1; 
32'd226: dataIn2 = 32'd0; 
32'd227: dataIn2 = 32'd1; 
32'd228: dataIn2 = 32'd1; 
32'd229: dataIn2 = 32'd0; 
32'd230: dataIn2 = 32'd0; 
32'd231: dataIn2 = 32'd0; 
32'd232: dataIn2 = 32'd1; 
32'd233: dataIn2 = 32'd1; 
32'd234: dataIn2 = 32'd0; 
32'd235: dataIn2 = 32'd1; 
32'd236: dataIn2 = 32'd1; 
32'd237: dataIn2 = 32'd1; 
32'd238: dataIn2 = 32'd0; 
32'd239: dataIn2 = 32'd1; 
32'd240: dataIn2 = 32'd0; 
32'd241: dataIn2 = 32'd1; 
32'd242: dataIn2 = 32'd1; 
32'd243: dataIn2 = 32'd1; 
32'd244: dataIn2 = 32'd0; 
32'd245: dataIn2 = 32'd0; 
32'd246: dataIn2 = 32'd0; 
32'd247: dataIn2 = 32'd1; 
32'd248: dataIn2 = 32'd1; 
32'd249: dataIn2 = 32'd0; 
32'd250: dataIn2 = 32'd1; 
32'd251: dataIn2 = 32'd0; 
32'd252: dataIn2 = 32'd0; 
32'd253: dataIn2 = 32'd1; 
32'd254: dataIn2 = 32'd1; 
32'd255: dataIn2 = 32'd1; 
32'd256: dataIn2 = 32'd0; 
32'd257: dataIn2 = 32'd1; 
32'd258: dataIn2 = 32'd0; 
32'd259: dataIn2 = 32'd0; 
32'd260: dataIn2 = 32'd1; 
32'd261: dataIn2 = 32'd0; 
32'd262: dataIn2 = 32'd0; 
32'd263: dataIn2 = 32'd1; 
32'd264: dataIn2 = 32'd0; 
32'd265: dataIn2 = 32'd0; 
32'd266: dataIn2 = 32'd1; 
32'd267: dataIn2 = 32'd1; 
32'd268: dataIn2 = 32'd1; 
32'd269: dataIn2 = 32'd1; 
32'd270: dataIn2 = 32'd0; 
32'd271: dataIn2 = 32'd0; 
32'd272: dataIn2 = 32'd0; 
32'd273: dataIn2 = 32'd0; 
32'd274: dataIn2 = 32'd1; 
32'd275: dataIn2 = 32'd1; 
32'd276: dataIn2 = 32'd1; 
32'd277: dataIn2 = 32'd0; 
32'd278: dataIn2 = 32'd0; 
32'd279: dataIn2 = 32'd0; 
32'd280: dataIn2 = 32'd1; 
32'd281: dataIn2 = 32'd0; 
32'd282: dataIn2 = 32'd1; 
32'd283: dataIn2 = 32'd1; 
32'd284: dataIn2 = 32'd1; 
32'd285: dataIn2 = 32'd0; 
32'd286: dataIn2 = 32'd1; 
32'd287: dataIn2 = 32'd0; 
32'd288: dataIn2 = 32'd1; 
32'd289: dataIn2 = 32'd0; 
32'd290: dataIn2 = 32'd0; 
32'd291: dataIn2 = 32'd1; 
32'd292: dataIn2 = 32'd1; 
32'd293: dataIn2 = 32'd1; 
32'd294: dataIn2 = 32'd1; 
32'd295: dataIn2 = 32'd1; 
32'd296: dataIn2 = 32'd1; 
32'd297: dataIn2 = 32'd0; 
32'd298: dataIn2 = 32'd0; 
32'd299: dataIn2 = 32'd1; 
32'd300: dataIn2 = 32'd0; 
32'd301: dataIn2 = 32'd1; 
32'd302: dataIn2 = 32'd0; 
32'd303: dataIn2 = 32'd1; 
32'd304: dataIn2 = 32'd1; 
32'd305: dataIn2 = 32'd0; 
32'd306: dataIn2 = 32'd0; 
32'd307: dataIn2 = 32'd1; 
32'd308: dataIn2 = 32'd0; 
32'd309: dataIn2 = 32'd1; 
32'd310: dataIn2 = 32'd0; 
32'd311: dataIn2 = 32'd0; 
32'd312: dataIn2 = 32'd0; 
32'd313: dataIn2 = 32'd0; 
32'd314: dataIn2 = 32'd1; 
32'd315: dataIn2 = 32'd1; 
32'd316: dataIn2 = 32'd0; 
32'd317: dataIn2 = 32'd1; 
32'd318: dataIn2 = 32'd1; 
32'd319: dataIn2 = 32'd1; 
32'd320: dataIn2 = 32'd0; 
32'd321: dataIn2 = 32'd0; 
32'd322: dataIn2 = 32'd0; 
32'd323: dataIn2 = 32'd0; 
32'd324: dataIn2 = 32'd1; 
32'd325: dataIn2 = 32'd1; 
32'd326: dataIn2 = 32'd0; 
32'd327: dataIn2 = 32'd1; 
32'd328: dataIn2 = 32'd1; 
32'd329: dataIn2 = 32'd0; 
32'd330: dataIn2 = 32'd0; 
32'd331: dataIn2 = 32'd1; 
32'd332: dataIn2 = 32'd1; 
32'd333: dataIn2 = 32'd1; 
32'd334: dataIn2 = 32'd0; 
32'd335: dataIn2 = 32'd0; 
32'd336: dataIn2 = 32'd1; 
32'd337: dataIn2 = 32'd1; 
32'd338: dataIn2 = 32'd1; 
32'd339: dataIn2 = 32'd1; 
32'd340: dataIn2 = 32'd1; 
32'd341: dataIn2 = 32'd1; 
32'd342: dataIn2 = 32'd1; 
32'd343: dataIn2 = 32'd0; 
32'd344: dataIn2 = 32'd0; 
32'd345: dataIn2 = 32'd0; 
32'd346: dataIn2 = 32'd0; 
32'd347: dataIn2 = 32'd1; 
32'd348: dataIn2 = 32'd1; 
32'd349: dataIn2 = 32'd1; 
32'd350: dataIn2 = 32'd0; 
32'd351: dataIn2 = 32'd1; 
32'd352: dataIn2 = 32'd1; 
32'd353: dataIn2 = 32'd1; 
32'd354: dataIn2 = 32'd0; 
32'd355: dataIn2 = 32'd1; 
32'd356: dataIn2 = 32'd0; 
32'd357: dataIn2 = 32'd0; 
32'd358: dataIn2 = 32'd1; 
32'd359: dataIn2 = 32'd0; 
32'd360: dataIn2 = 32'd0; 
32'd361: dataIn2 = 32'd0; 
32'd362: dataIn2 = 32'd0; 
32'd363: dataIn2 = 32'd1; 
32'd364: dataIn2 = 32'd0; 
32'd365: dataIn2 = 32'd1; 
32'd366: dataIn2 = 32'd0; 
32'd367: dataIn2 = 32'd1; 
32'd368: dataIn2 = 32'd0; 
32'd369: dataIn2 = 32'd1; 
32'd370: dataIn2 = 32'd1; 
32'd371: dataIn2 = 32'd1; 
32'd372: dataIn2 = 32'd1; 
32'd373: dataIn2 = 32'd0; 
32'd374: dataIn2 = 32'd0; 
32'd375: dataIn2 = 32'd1; 
32'd376: dataIn2 = 32'd0; 
32'd377: dataIn2 = 32'd1; 
32'd378: dataIn2 = 32'd0; 
32'd379: dataIn2 = 32'd0; 
32'd380: dataIn2 = 32'd0; 
32'd381: dataIn2 = 32'd0; 
32'd382: dataIn2 = 32'd0; 
32'd383: dataIn2 = 32'd1; 
32'd384: dataIn2 = 32'd1; 
32'd385: dataIn2 = 32'd1; 
32'd386: dataIn2 = 32'd0; 
32'd387: dataIn2 = 32'd1; 
32'd388: dataIn2 = 32'd1; 
32'd389: dataIn2 = 32'd0; 
32'd390: dataIn2 = 32'd1; 
32'd391: dataIn2 = 32'd1; 
32'd392: dataIn2 = 32'd0; 
32'd393: dataIn2 = 32'd0; 
32'd394: dataIn2 = 32'd0; 
32'd395: dataIn2 = 32'd1; 
32'd396: dataIn2 = 32'd0; 
32'd397: dataIn2 = 32'd0; 
32'd398: dataIn2 = 32'd1; 
32'd399: dataIn2 = 32'd0; 
32'd400: dataIn2 = 32'd0; 
32'd401: dataIn2 = 32'd0; 
32'd402: dataIn2 = 32'd0; 
32'd403: dataIn2 = 32'd0; 
32'd404: dataIn2 = 32'd0; 
32'd405: dataIn2 = 32'd0; 
32'd406: dataIn2 = 32'd0; 
32'd407: dataIn2 = 32'd1; 
32'd408: dataIn2 = 32'd1; 
32'd409: dataIn2 = 32'd1; 
32'd410: dataIn2 = 32'd0; 
32'd411: dataIn2 = 32'd1; 
32'd412: dataIn2 = 32'd1; 
32'd413: dataIn2 = 32'd1; 
32'd414: dataIn2 = 32'd0; 
32'd415: dataIn2 = 32'd1; 
32'd416: dataIn2 = 32'd1; 
32'd417: dataIn2 = 32'd0; 
32'd418: dataIn2 = 32'd1; 
32'd419: dataIn2 = 32'd1; 
32'd420: dataIn2 = 32'd1; 
32'd421: dataIn2 = 32'd0; 
32'd422: dataIn2 = 32'd1; 
32'd423: dataIn2 = 32'd1; 
32'd424: dataIn2 = 32'd1; 
32'd425: dataIn2 = 32'd1; 
32'd426: dataIn2 = 32'd0; 
32'd427: dataIn2 = 32'd1; 
32'd428: dataIn2 = 32'd1; 
32'd429: dataIn2 = 32'd1; 
32'd430: dataIn2 = 32'd0; 
32'd431: dataIn2 = 32'd0; 
32'd432: dataIn2 = 32'd0; 
32'd433: dataIn2 = 32'd0; 
32'd434: dataIn2 = 32'd0; 
32'd435: dataIn2 = 32'd0; 
32'd436: dataIn2 = 32'd0; 
32'd437: dataIn2 = 32'd0; 
32'd438: dataIn2 = 32'd0; 
32'd439: dataIn2 = 32'd1; 
32'd440: dataIn2 = 32'd0; 
32'd441: dataIn2 = 32'd0; 
32'd442: dataIn2 = 32'd0; 
32'd443: dataIn2 = 32'd0; 
32'd444: dataIn2 = 32'd1; 
32'd445: dataIn2 = 32'd0; 
32'd446: dataIn2 = 32'd1; 
32'd447: dataIn2 = 32'd0; 
32'd448: dataIn2 = 32'd0; 
32'd449: dataIn2 = 32'd1; 
32'd450: dataIn2 = 32'd1; 
32'd451: dataIn2 = 32'd1; 
32'd452: dataIn2 = 32'd0; 
32'd453: dataIn2 = 32'd1; 
32'd454: dataIn2 = 32'd0; 
32'd455: dataIn2 = 32'd0; 
32'd456: dataIn2 = 32'd0; 
32'd457: dataIn2 = 32'd1; 
32'd458: dataIn2 = 32'd0; 
32'd459: dataIn2 = 32'd0; 
32'd460: dataIn2 = 32'd0; 
32'd461: dataIn2 = 32'd0; 
32'd462: dataIn2 = 32'd1; 
32'd463: dataIn2 = 32'd1; 
32'd464: dataIn2 = 32'd1; 
32'd465: dataIn2 = 32'd0; 
32'd466: dataIn2 = 32'd1; 
32'd467: dataIn2 = 32'd1; 
32'd468: dataIn2 = 32'd0; 
32'd469: dataIn2 = 32'd1; 
32'd470: dataIn2 = 32'd1; 
32'd471: dataIn2 = 32'd0; 
32'd472: dataIn2 = 32'd0; 
32'd473: dataIn2 = 32'd1; 
32'd474: dataIn2 = 32'd1; 
32'd475: dataIn2 = 32'd0; 
32'd476: dataIn2 = 32'd0; 
32'd477: dataIn2 = 32'd0; 
32'd478: dataIn2 = 32'd1; 
32'd479: dataIn2 = 32'd1; 
32'd480: dataIn2 = 32'd1; 
32'd481: dataIn2 = 32'd1; 
32'd482: dataIn2 = 32'd0; 
32'd483: dataIn2 = 32'd1; 
32'd484: dataIn2 = 32'd0; 
32'd485: dataIn2 = 32'd1; 
32'd486: dataIn2 = 32'd0; 
32'd487: dataIn2 = 32'd1; 
32'd488: dataIn2 = 32'd0; 
32'd489: dataIn2 = 32'd1; 
32'd490: dataIn2 = 32'd1; 
32'd491: dataIn2 = 32'd1; 
32'd492: dataIn2 = 32'd1; 
32'd493: dataIn2 = 32'd0; 
32'd494: dataIn2 = 32'd1; 
32'd495: dataIn2 = 32'd1; 
32'd496: dataIn2 = 32'd1; 
32'd497: dataIn2 = 32'd0; 
32'd498: dataIn2 = 32'd1; 
32'd499: dataIn2 = 32'd1; 
32'd500: dataIn2 = 32'd0; 
32'd501: dataIn2 = 32'd1; 
32'd502: dataIn2 = 32'd1; 
32'd503: dataIn2 = 32'd0; 
32'd504: dataIn2 = 32'd1; 
32'd505: dataIn2 = 32'd1; 
32'd506: dataIn2 = 32'd0; 
32'd507: dataIn2 = 32'd1; 
32'd508: dataIn2 = 32'd0; 
32'd509: dataIn2 = 32'd1; 
32'd510: dataIn2 = 32'd1; 
32'd511: dataIn2 = 32'd1; 
32'd512: dataIn2 = 32'd0; 
32'd513: dataIn2 = 32'd1; 
32'd514: dataIn2 = 32'd1; 
32'd515: dataIn2 = 32'd1; 
32'd516: dataIn2 = 32'd0; 
32'd517: dataIn2 = 32'd0; 
32'd518: dataIn2 = 32'd1; 
32'd519: dataIn2 = 32'd0; 
32'd520: dataIn2 = 32'd1; 
32'd521: dataIn2 = 32'd0; 
32'd522: dataIn2 = 32'd0; 
32'd523: dataIn2 = 32'd0; 
32'd524: dataIn2 = 32'd1; 
32'd525: dataIn2 = 32'd0; 
32'd526: dataIn2 = 32'd0; 
32'd527: dataIn2 = 32'd1; 
32'd528: dataIn2 = 32'd1; 
32'd529: dataIn2 = 32'd1; 
32'd530: dataIn2 = 32'd1; 
32'd531: dataIn2 = 32'd0; 
32'd532: dataIn2 = 32'd1; 
32'd533: dataIn2 = 32'd0; 
32'd534: dataIn2 = 32'd1; 
32'd535: dataIn2 = 32'd0; 
32'd536: dataIn2 = 32'd0; 
32'd537: dataIn2 = 32'd1; 
32'd538: dataIn2 = 32'd1; 
32'd539: dataIn2 = 32'd1; 
32'd540: dataIn2 = 32'd0; 
32'd541: dataIn2 = 32'd1; 
32'd542: dataIn2 = 32'd1; 
32'd543: dataIn2 = 32'd1; 
32'd544: dataIn2 = 32'd0; 
32'd545: dataIn2 = 32'd0; 
32'd546: dataIn2 = 32'd0; 
32'd547: dataIn2 = 32'd1; 
32'd548: dataIn2 = 32'd1; 
32'd549: dataIn2 = 32'd1; 
32'd550: dataIn2 = 32'd0; 
32'd551: dataIn2 = 32'd0; 
32'd552: dataIn2 = 32'd1; 
32'd553: dataIn2 = 32'd1; 
32'd554: dataIn2 = 32'd0; 
32'd555: dataIn2 = 32'd1; 
32'd556: dataIn2 = 32'd0; 
32'd557: dataIn2 = 32'd1; 
32'd558: dataIn2 = 32'd0; 
32'd559: dataIn2 = 32'd0; 
32'd560: dataIn2 = 32'd1; 
32'd561: dataIn2 = 32'd1; 
32'd562: dataIn2 = 32'd1; 
32'd563: dataIn2 = 32'd0; 
32'd564: dataIn2 = 32'd1; 
32'd565: dataIn2 = 32'd1; 
32'd566: dataIn2 = 32'd1; 
32'd567: dataIn2 = 32'd0; 
32'd568: dataIn2 = 32'd1; 
32'd569: dataIn2 = 32'd1; 
32'd570: dataIn2 = 32'd1; 
32'd571: dataIn2 = 32'd0; 
32'd572: dataIn2 = 32'd0; 
32'd573: dataIn2 = 32'd1; 
32'd574: dataIn2 = 32'd1; 
32'd575: dataIn2 = 32'd1; 
32'd576: dataIn2 = 32'd1; 
32'd577: dataIn2 = 32'd0; 
32'd578: dataIn2 = 32'd0; 
32'd579: dataIn2 = 32'd1; 
32'd580: dataIn2 = 32'd0; 
32'd581: dataIn2 = 32'd0; 
32'd582: dataIn2 = 32'd1; 
32'd583: dataIn2 = 32'd0; 
32'd584: dataIn2 = 32'd1; 
32'd585: dataIn2 = 32'd1; 
32'd586: dataIn2 = 32'd1; 
32'd587: dataIn2 = 32'd1; 
32'd588: dataIn2 = 32'd0; 
32'd589: dataIn2 = 32'd0; 
32'd590: dataIn2 = 32'd1; 
32'd591: dataIn2 = 32'd0; 
32'd592: dataIn2 = 32'd1; 
32'd593: dataIn2 = 32'd0; 
32'd594: dataIn2 = 32'd1; 
32'd595: dataIn2 = 32'd0; 
32'd596: dataIn2 = 32'd1; 
32'd597: dataIn2 = 32'd0; 
32'd598: dataIn2 = 32'd1; 
32'd599: dataIn2 = 32'd0; 
32'd600: dataIn2 = 32'd1; 
32'd601: dataIn2 = 32'd1; 
32'd602: dataIn2 = 32'd1; 
32'd603: dataIn2 = 32'd1; 
32'd604: dataIn2 = 32'd1; 
32'd605: dataIn2 = 32'd0; 
32'd606: dataIn2 = 32'd1; 
32'd607: dataIn2 = 32'd1; 
32'd608: dataIn2 = 32'd1; 
32'd609: dataIn2 = 32'd1; 
32'd610: dataIn2 = 32'd0; 
32'd611: dataIn2 = 32'd0; 
32'd612: dataIn2 = 32'd0; 
32'd613: dataIn2 = 32'd1; 
32'd614: dataIn2 = 32'd1; 
32'd615: dataIn2 = 32'd1; 
32'd616: dataIn2 = 32'd0; 
32'd617: dataIn2 = 32'd1; 
32'd618: dataIn2 = 32'd1; 
32'd619: dataIn2 = 32'd0; 
32'd620: dataIn2 = 32'd1; 
32'd621: dataIn2 = 32'd1; 
32'd622: dataIn2 = 32'd1; 
32'd623: dataIn2 = 32'd1; 
32'd624: dataIn2 = 32'd0; 
32'd625: dataIn2 = 32'd0; 
32'd626: dataIn2 = 32'd1; 
32'd627: dataIn2 = 32'd0; 
32'd628: dataIn2 = 32'd0; 
32'd629: dataIn2 = 32'd0; 
32'd630: dataIn2 = 32'd0; 
32'd631: dataIn2 = 32'd1; 
32'd632: dataIn2 = 32'd0; 
32'd633: dataIn2 = 32'd1; 
32'd634: dataIn2 = 32'd1; 
32'd635: dataIn2 = 32'd1; 
32'd636: dataIn2 = 32'd1; 
32'd637: dataIn2 = 32'd0; 
32'd638: dataIn2 = 32'd1; 
32'd639: dataIn2 = 32'd0; 
32'd640: dataIn2 = 32'd1; 
32'd641: dataIn2 = 32'd0; 
32'd642: dataIn2 = 32'd0; 
32'd643: dataIn2 = 32'd1; 
32'd644: dataIn2 = 32'd0; 
32'd645: dataIn2 = 32'd0; 
32'd646: dataIn2 = 32'd0; 
32'd647: dataIn2 = 32'd0; 
32'd648: dataIn2 = 32'd1; 
32'd649: dataIn2 = 32'd0; 
32'd650: dataIn2 = 32'd1; 
32'd651: dataIn2 = 32'd0; 
32'd652: dataIn2 = 32'd1; 
32'd653: dataIn2 = 32'd0; 
32'd654: dataIn2 = 32'd0; 
32'd655: dataIn2 = 32'd1; 
32'd656: dataIn2 = 32'd0; 
32'd657: dataIn2 = 32'd1; 
32'd658: dataIn2 = 32'd1; 
32'd659: dataIn2 = 32'd1; 
32'd660: dataIn2 = 32'd0; 
32'd661: dataIn2 = 32'd1; 
32'd662: dataIn2 = 32'd1; 
32'd663: dataIn2 = 32'd1; 
32'd664: dataIn2 = 32'd0; 
32'd665: dataIn2 = 32'd1; 
32'd666: dataIn2 = 32'd1; 
32'd667: dataIn2 = 32'd1; 
32'd668: dataIn2 = 32'd0; 
32'd669: dataIn2 = 32'd1; 
32'd670: dataIn2 = 32'd0; 
32'd671: dataIn2 = 32'd0; 
32'd672: dataIn2 = 32'd0; 
32'd673: dataIn2 = 32'd1; 
32'd674: dataIn2 = 32'd0; 
32'd675: dataIn2 = 32'd1; 
32'd676: dataIn2 = 32'd0; 
32'd677: dataIn2 = 32'd0; 
32'd678: dataIn2 = 32'd1; 
32'd679: dataIn2 = 32'd1; 
32'd680: dataIn2 = 32'd1; 
32'd681: dataIn2 = 32'd0; 
32'd682: dataIn2 = 32'd1; 
32'd683: dataIn2 = 32'd0; 
32'd684: dataIn2 = 32'd1; 
32'd685: dataIn2 = 32'd0; 
32'd686: dataIn2 = 32'd0; 
32'd687: dataIn2 = 32'd1; 
32'd688: dataIn2 = 32'd1; 
32'd689: dataIn2 = 32'd1; 
32'd690: dataIn2 = 32'd0; 
32'd691: dataIn2 = 32'd0; 
32'd692: dataIn2 = 32'd1; 
32'd693: dataIn2 = 32'd0; 
32'd694: dataIn2 = 32'd1; 
32'd695: dataIn2 = 32'd1; 
32'd696: dataIn2 = 32'd0; 
32'd697: dataIn2 = 32'd0; 
32'd698: dataIn2 = 32'd0; 
32'd699: dataIn2 = 32'd0; 
32'd700: dataIn2 = 32'd0; 
32'd701: dataIn2 = 32'd0; 
32'd702: dataIn2 = 32'd1; 
32'd703: dataIn2 = 32'd1; 
32'd704: dataIn2 = 32'd0; 
32'd705: dataIn2 = 32'd0; 
32'd706: dataIn2 = 32'd1; 
32'd707: dataIn2 = 32'd1; 
32'd708: dataIn2 = 32'd1; 
32'd709: dataIn2 = 32'd0; 
32'd710: dataIn2 = 32'd1; 
32'd711: dataIn2 = 32'd0; 
32'd712: dataIn2 = 32'd0; 
32'd713: dataIn2 = 32'd0; 
32'd714: dataIn2 = 32'd0; 
32'd715: dataIn2 = 32'd1; 
32'd716: dataIn2 = 32'd0; 
32'd717: dataIn2 = 32'd0; 
32'd718: dataIn2 = 32'd1; 
32'd719: dataIn2 = 32'd0; 
32'd720: dataIn2 = 32'd1; 
32'd721: dataIn2 = 32'd1; 
32'd722: dataIn2 = 32'd0; 
32'd723: dataIn2 = 32'd1; 
32'd724: dataIn2 = 32'd0; 
32'd725: dataIn2 = 32'd0; 
32'd726: dataIn2 = 32'd0; 
32'd727: dataIn2 = 32'd1; 
32'd728: dataIn2 = 32'd1; 
32'd729: dataIn2 = 32'd1; 
32'd730: dataIn2 = 32'd0; 
32'd731: dataIn2 = 32'd0; 
32'd732: dataIn2 = 32'd1; 
32'd733: dataIn2 = 32'd0; 
32'd734: dataIn2 = 32'd0; 
32'd735: dataIn2 = 32'd0; 
32'd736: dataIn2 = 32'd0; 
32'd737: dataIn2 = 32'd1; 
32'd738: dataIn2 = 32'd0; 
32'd739: dataIn2 = 32'd1; 
32'd740: dataIn2 = 32'd1; 
32'd741: dataIn2 = 32'd1; 
32'd742: dataIn2 = 32'd0; 
32'd743: dataIn2 = 32'd0; 
32'd744: dataIn2 = 32'd1; 
32'd745: dataIn2 = 32'd1; 
32'd746: dataIn2 = 32'd0; 
32'd747: dataIn2 = 32'd1; 
32'd748: dataIn2 = 32'd1; 
32'd749: dataIn2 = 32'd1; 
32'd750: dataIn2 = 32'd1; 
32'd751: dataIn2 = 32'd1; 
32'd752: dataIn2 = 32'd0; 
32'd753: dataIn2 = 32'd0; 
32'd754: dataIn2 = 32'd1; 
32'd755: dataIn2 = 32'd1; 
32'd756: dataIn2 = 32'd1; 
32'd757: dataIn2 = 32'd1; 
32'd758: dataIn2 = 32'd0; 
32'd759: dataIn2 = 32'd0; 
32'd760: dataIn2 = 32'd0; 
32'd761: dataIn2 = 32'd1; 
32'd762: dataIn2 = 32'd0; 
32'd763: dataIn2 = 32'd0; 
32'd764: dataIn2 = 32'd1; 
32'd765: dataIn2 = 32'd1; 
32'd766: dataIn2 = 32'd0; 
32'd767: dataIn2 = 32'd0; 
32'd768: dataIn2 = 32'd1; 
32'd769: dataIn2 = 32'd1; 
32'd770: dataIn2 = 32'd0; 
32'd771: dataIn2 = 32'd0; 
32'd772: dataIn2 = 32'd1; 
32'd773: dataIn2 = 32'd0; 
32'd774: dataIn2 = 32'd0; 
32'd775: dataIn2 = 32'd1; 
32'd776: dataIn2 = 32'd0; 
32'd777: dataIn2 = 32'd1; 
32'd778: dataIn2 = 32'd0; 
32'd779: dataIn2 = 32'd0; 
32'd780: dataIn2 = 32'd1; 
32'd781: dataIn2 = 32'd1; 
32'd782: dataIn2 = 32'd0; 
32'd783: dataIn2 = 32'd0; 
32'd784: dataIn2 = 32'd0; 
32'd785: dataIn2 = 32'd1; 
32'd786: dataIn2 = 32'd0; 
32'd787: dataIn2 = 32'd1; 
32'd788: dataIn2 = 32'd1; 
32'd789: dataIn2 = 32'd1; 
32'd790: dataIn2 = 32'd0; 
32'd791: dataIn2 = 32'd0; 
32'd792: dataIn2 = 32'd1; 
32'd793: dataIn2 = 32'd1; 
32'd794: dataIn2 = 32'd0; 
32'd795: dataIn2 = 32'd0; 
32'd796: dataIn2 = 32'd1; 
32'd797: dataIn2 = 32'd1; 
32'd798: dataIn2 = 32'd1; 
32'd799: dataIn2 = 32'd0; 
32'd800: dataIn2 = 32'd1; 
32'd801: dataIn2 = 32'd0; 
32'd802: dataIn2 = 32'd0; 
32'd803: dataIn2 = 32'd1; 
32'd804: dataIn2 = 32'd1; 
32'd805: dataIn2 = 32'd1; 
32'd806: dataIn2 = 32'd0; 
32'd807: dataIn2 = 32'd0; 
32'd808: dataIn2 = 32'd0; 
32'd809: dataIn2 = 32'd0; 
32'd810: dataIn2 = 32'd1; 
32'd811: dataIn2 = 32'd1; 
32'd812: dataIn2 = 32'd1; 
32'd813: dataIn2 = 32'd1; 
32'd814: dataIn2 = 32'd1; 
32'd815: dataIn2 = 32'd1; 
32'd816: dataIn2 = 32'd1; 
32'd817: dataIn2 = 32'd1; 
32'd818: dataIn2 = 32'd1; 
32'd819: dataIn2 = 32'd0; 
32'd820: dataIn2 = 32'd0; 
32'd821: dataIn2 = 32'd0; 
32'd822: dataIn2 = 32'd0; 
32'd823: dataIn2 = 32'd0; 
32'd824: dataIn2 = 32'd0; 
32'd825: dataIn2 = 32'd0; 
32'd826: dataIn2 = 32'd1; 
32'd827: dataIn2 = 32'd0; 
32'd828: dataIn2 = 32'd0; 
32'd829: dataIn2 = 32'd0; 
32'd830: dataIn2 = 32'd0; 
32'd831: dataIn2 = 32'd1; 
32'd832: dataIn2 = 32'd1; 
32'd833: dataIn2 = 32'd1; 
32'd834: dataIn2 = 32'd0; 
32'd835: dataIn2 = 32'd0; 
32'd836: dataIn2 = 32'd0; 
32'd837: dataIn2 = 32'd0; 
32'd838: dataIn2 = 32'd1; 
32'd839: dataIn2 = 32'd0; 
32'd840: dataIn2 = 32'd1; 
32'd841: dataIn2 = 32'd1; 
32'd842: dataIn2 = 32'd1; 
32'd843: dataIn2 = 32'd0; 
32'd844: dataIn2 = 32'd0; 
32'd845: dataIn2 = 32'd0; 
32'd846: dataIn2 = 32'd1; 
32'd847: dataIn2 = 32'd0; 
32'd848: dataIn2 = 32'd1; 
32'd849: dataIn2 = 32'd0; 
32'd850: dataIn2 = 32'd1; 
32'd851: dataIn2 = 32'd0; 
32'd852: dataIn2 = 32'd1; 
32'd853: dataIn2 = 32'd1; 
32'd854: dataIn2 = 32'd1; 
32'd855: dataIn2 = 32'd1; 
32'd856: dataIn2 = 32'd1; 
32'd857: dataIn2 = 32'd1; 
32'd858: dataIn2 = 32'd0; 
32'd859: dataIn2 = 32'd1; 
32'd860: dataIn2 = 32'd1; 
32'd861: dataIn2 = 32'd0; 
32'd862: dataIn2 = 32'd1; 
32'd863: dataIn2 = 32'd1; 
32'd864: dataIn2 = 32'd0; 
32'd865: dataIn2 = 32'd0; 
32'd866: dataIn2 = 32'd0; 
32'd867: dataIn2 = 32'd1; 
32'd868: dataIn2 = 32'd1; 
32'd869: dataIn2 = 32'd0; 
32'd870: dataIn2 = 32'd1; 
32'd871: dataIn2 = 32'd0; 
32'd872: dataIn2 = 32'd0; 
32'd873: dataIn2 = 32'd1; 
32'd874: dataIn2 = 32'd1; 
32'd875: dataIn2 = 32'd1; 
32'd876: dataIn2 = 32'd1; 
32'd877: dataIn2 = 32'd0; 
32'd878: dataIn2 = 32'd0; 
32'd879: dataIn2 = 32'd0; 
32'd880: dataIn2 = 32'd0; 
32'd881: dataIn2 = 32'd0; 
32'd882: dataIn2 = 32'd0; 
32'd883: dataIn2 = 32'd0; 
32'd884: dataIn2 = 32'd0; 
32'd885: dataIn2 = 32'd1; 
32'd886: dataIn2 = 32'd1; 
32'd887: dataIn2 = 32'd1; 
32'd888: dataIn2 = 32'd0; 
32'd889: dataIn2 = 32'd1; 
32'd890: dataIn2 = 32'd1; 
32'd891: dataIn2 = 32'd0; 
32'd892: dataIn2 = 32'd0; 
32'd893: dataIn2 = 32'd0; 
32'd894: dataIn2 = 32'd1; 
32'd895: dataIn2 = 32'd0; 
32'd896: dataIn2 = 32'd1; 
32'd897: dataIn2 = 32'd1; 
32'd898: dataIn2 = 32'd0; 
32'd899: dataIn2 = 32'd0; 
32'd900: dataIn2 = 32'd0; 
32'd901: dataIn2 = 32'd0; 
32'd902: dataIn2 = 32'd0; 
32'd903: dataIn2 = 32'd1; 
32'd904: dataIn2 = 32'd0; 
32'd905: dataIn2 = 32'd1; 
32'd906: dataIn2 = 32'd0; 
32'd907: dataIn2 = 32'd0; 
32'd908: dataIn2 = 32'd1; 
32'd909: dataIn2 = 32'd1; 
32'd910: dataIn2 = 32'd0; 
32'd911: dataIn2 = 32'd1; 
32'd912: dataIn2 = 32'd1; 
32'd913: dataIn2 = 32'd0; 
32'd914: dataIn2 = 32'd0; 
32'd915: dataIn2 = 32'd0; 
32'd916: dataIn2 = 32'd1; 
32'd917: dataIn2 = 32'd1; 
32'd918: dataIn2 = 32'd1; 
32'd919: dataIn2 = 32'd0; 
32'd920: dataIn2 = 32'd0; 
32'd921: dataIn2 = 32'd1; 
32'd922: dataIn2 = 32'd1; 
32'd923: dataIn2 = 32'd0; 
32'd924: dataIn2 = 32'd1; 
32'd925: dataIn2 = 32'd1; 
32'd926: dataIn2 = 32'd1; 
32'd927: dataIn2 = 32'd0; 
32'd928: dataIn2 = 32'd1; 
32'd929: dataIn2 = 32'd0; 
32'd930: dataIn2 = 32'd1; 
32'd931: dataIn2 = 32'd0; 
32'd932: dataIn2 = 32'd0; 
32'd933: dataIn2 = 32'd1; 
32'd934: dataIn2 = 32'd1; 
32'd935: dataIn2 = 32'd0; 
32'd936: dataIn2 = 32'd0; 
32'd937: dataIn2 = 32'd1; 
32'd938: dataIn2 = 32'd1; 
32'd939: dataIn2 = 32'd1; 
32'd940: dataIn2 = 32'd0; 
32'd941: dataIn2 = 32'd1; 
32'd942: dataIn2 = 32'd1; 
32'd943: dataIn2 = 32'd1; 
32'd944: dataIn2 = 32'd1; 
32'd945: dataIn2 = 32'd0; 
32'd946: dataIn2 = 32'd0; 
32'd947: dataIn2 = 32'd0; 
32'd948: dataIn2 = 32'd0; 
32'd949: dataIn2 = 32'd1; 
32'd950: dataIn2 = 32'd0; 
32'd951: dataIn2 = 32'd0; 
32'd952: dataIn2 = 32'd0; 
32'd953: dataIn2 = 32'd1; 
32'd954: dataIn2 = 32'd0; 
32'd955: dataIn2 = 32'd1; 
32'd956: dataIn2 = 32'd1; 
32'd957: dataIn2 = 32'd1; 
32'd958: dataIn2 = 32'd0; 
32'd959: dataIn2 = 32'd0; 
32'd960: dataIn2 = 32'd0; 
32'd961: dataIn2 = 32'd0; 
32'd962: dataIn2 = 32'd0; 
32'd963: dataIn2 = 32'd0; 
32'd964: dataIn2 = 32'd0; 
32'd965: dataIn2 = 32'd1; 
32'd966: dataIn2 = 32'd1; 
32'd967: dataIn2 = 32'd1; 
32'd968: dataIn2 = 32'd0; 
32'd969: dataIn2 = 32'd1; 
32'd970: dataIn2 = 32'd1; 
32'd971: dataIn2 = 32'd1; 
32'd972: dataIn2 = 32'd0; 
32'd973: dataIn2 = 32'd0; 
32'd974: dataIn2 = 32'd1; 
32'd975: dataIn2 = 32'd0; 
32'd976: dataIn2 = 32'd0; 
32'd977: dataIn2 = 32'd1; 
32'd978: dataIn2 = 32'd0; 
32'd979: dataIn2 = 32'd1; 
32'd980: dataIn2 = 32'd1; 
32'd981: dataIn2 = 32'd1; 
32'd982: dataIn2 = 32'd1; 
32'd983: dataIn2 = 32'd1; 
32'd984: dataIn2 = 32'd0; 
32'd985: dataIn2 = 32'd0; 
32'd986: dataIn2 = 32'd1; 
32'd987: dataIn2 = 32'd1; 
32'd988: dataIn2 = 32'd1; 
32'd989: dataIn2 = 32'd0; 
32'd990: dataIn2 = 32'd1; 
32'd991: dataIn2 = 32'd1; 
32'd992: dataIn2 = 32'd0; 
32'd993: dataIn2 = 32'd0; 
32'd994: dataIn2 = 32'd0; 
32'd995: dataIn2 = 32'd1; 
32'd996: dataIn2 = 32'd1; 
32'd997: dataIn2 = 32'd0; 
32'd998: dataIn2 = 32'd0; 
32'd999: dataIn2 = 32'd0; 
32'd1000: dataIn2 = 32'd0; 
32'd1001: dataIn2 = 32'd1; 
32'd1002: dataIn2 = 32'd0; 
32'd1003: dataIn2 = 32'd1; 
32'd1004: dataIn2 = 32'd0; 
32'd1005: dataIn2 = 32'd0; 
32'd1006: dataIn2 = 32'd1; 
32'd1007: dataIn2 = 32'd1; 
32'd1008: dataIn2 = 32'd1; 
32'd1009: dataIn2 = 32'd1; 
32'd1010: dataIn2 = 32'd0; 
32'd1011: dataIn2 = 32'd1; 
32'd1012: dataIn2 = 32'd1; 
32'd1013: dataIn2 = 32'd1; 
32'd1014: dataIn2 = 32'd1; 
32'd1015: dataIn2 = 32'd1; 
32'd1016: dataIn2 = 32'd0; 
32'd1017: dataIn2 = 32'd1; 
32'd1018: dataIn2 = 32'd0; 
32'd1019: dataIn2 = 32'd0; 
32'd1020: dataIn2 = 32'd1; 
32'd1021: dataIn2 = 32'd0; 
32'd1022: dataIn2 = 32'd0; 
32'd1023: dataIn2 = 32'd0; 
32'd1024: dataIn2 = 32'd0; 
32'd1025: dataIn2 = 32'd0; 
32'd1026: dataIn2 = 32'd0; 
32'd1027: dataIn2 = 32'd1; 
32'd1028: dataIn2 = 32'd0; 
32'd1029: dataIn2 = 32'd0; 
32'd1030: dataIn2 = 32'd1; 
32'd1031: dataIn2 = 32'd1; 
32'd1032: dataIn2 = 32'd0; 
32'd1033: dataIn2 = 32'd0; 
32'd1034: dataIn2 = 32'd1; 
32'd1035: dataIn2 = 32'd1; 
32'd1036: dataIn2 = 32'd0; 
32'd1037: dataIn2 = 32'd0; 
32'd1038: dataIn2 = 32'd0; 
32'd1039: dataIn2 = 32'd0; 
32'd1040: dataIn2 = 32'd1; 
32'd1041: dataIn2 = 32'd0; 
32'd1042: dataIn2 = 32'd1; 
32'd1043: dataIn2 = 32'd1; 
32'd1044: dataIn2 = 32'd0; 
32'd1045: dataIn2 = 32'd0; 
32'd1046: dataIn2 = 32'd0; 
32'd1047: dataIn2 = 32'd0; 
32'd1048: dataIn2 = 32'd0; 
32'd1049: dataIn2 = 32'd0; 
32'd1050: dataIn2 = 32'd1; 
32'd1051: dataIn2 = 32'd0; 
32'd1052: dataIn2 = 32'd1; 
32'd1053: dataIn2 = 32'd1; 
32'd1054: dataIn2 = 32'd1; 
32'd1055: dataIn2 = 32'd0; 
32'd1056: dataIn2 = 32'd0; 
32'd1057: dataIn2 = 32'd1; 
32'd1058: dataIn2 = 32'd1; 
32'd1059: dataIn2 = 32'd0; 
32'd1060: dataIn2 = 32'd1; 
32'd1061: dataIn2 = 32'd1; 
32'd1062: dataIn2 = 32'd1; 
32'd1063: dataIn2 = 32'd0; 
32'd1064: dataIn2 = 32'd0; 
32'd1065: dataIn2 = 32'd0; 
32'd1066: dataIn2 = 32'd1; 
32'd1067: dataIn2 = 32'd0; 
32'd1068: dataIn2 = 32'd1; 
32'd1069: dataIn2 = 32'd0; 
32'd1070: dataIn2 = 32'd0; 
32'd1071: dataIn2 = 32'd0; 
32'd1072: dataIn2 = 32'd0; 
32'd1073: dataIn2 = 32'd1; 
32'd1074: dataIn2 = 32'd1; 
32'd1075: dataIn2 = 32'd1; 
32'd1076: dataIn2 = 32'd1; 
32'd1077: dataIn2 = 32'd0; 
32'd1078: dataIn2 = 32'd0; 
32'd1079: dataIn2 = 32'd1; 
32'd1080: dataIn2 = 32'd0; 
32'd1081: dataIn2 = 32'd1; 
32'd1082: dataIn2 = 32'd1; 
32'd1083: dataIn2 = 32'd0; 
32'd1084: dataIn2 = 32'd0; 
32'd1085: dataIn2 = 32'd0; 
32'd1086: dataIn2 = 32'd1; 
32'd1087: dataIn2 = 32'd1; 
32'd1088: dataIn2 = 32'd1; 
32'd1089: dataIn2 = 32'd0; 
32'd1090: dataIn2 = 32'd0; 
32'd1091: dataIn2 = 32'd1; 
32'd1092: dataIn2 = 32'd0; 
32'd1093: dataIn2 = 32'd1; 
32'd1094: dataIn2 = 32'd1; 
32'd1095: dataIn2 = 32'd0; 
32'd1096: dataIn2 = 32'd0; 
32'd1097: dataIn2 = 32'd1; 
32'd1098: dataIn2 = 32'd1; 
32'd1099: dataIn2 = 32'd0; 
32'd1100: dataIn2 = 32'd0; 
32'd1101: dataIn2 = 32'd0; 
32'd1102: dataIn2 = 32'd0; 
32'd1103: dataIn2 = 32'd0; 
32'd1104: dataIn2 = 32'd1; 
32'd1105: dataIn2 = 32'd0; 
32'd1106: dataIn2 = 32'd0; 
32'd1107: dataIn2 = 32'd1; 
32'd1108: dataIn2 = 32'd0; 
32'd1109: dataIn2 = 32'd1; 
32'd1110: dataIn2 = 32'd1; 
32'd1111: dataIn2 = 32'd0; 
32'd1112: dataIn2 = 32'd1; 
32'd1113: dataIn2 = 32'd0; 
32'd1114: dataIn2 = 32'd1; 
32'd1115: dataIn2 = 32'd0; 
32'd1116: dataIn2 = 32'd1; 
32'd1117: dataIn2 = 32'd1; 
32'd1118: dataIn2 = 32'd0; 
32'd1119: dataIn2 = 32'd0; 
32'd1120: dataIn2 = 32'd0; 
32'd1121: dataIn2 = 32'd0; 
32'd1122: dataIn2 = 32'd0; 
32'd1123: dataIn2 = 32'd0; 
32'd1124: dataIn2 = 32'd1; 
32'd1125: dataIn2 = 32'd1; 
32'd1126: dataIn2 = 32'd0; 
32'd1127: dataIn2 = 32'd0; 
32'd1128: dataIn2 = 32'd0; 
32'd1129: dataIn2 = 32'd0; 
32'd1130: dataIn2 = 32'd1; 
32'd1131: dataIn2 = 32'd1; 
32'd1132: dataIn2 = 32'd0; 
32'd1133: dataIn2 = 32'd0; 
32'd1134: dataIn2 = 32'd0; 
32'd1135: dataIn2 = 32'd0; 
32'd1136: dataIn2 = 32'd0; 
32'd1137: dataIn2 = 32'd0; 
32'd1138: dataIn2 = 32'd0; 
32'd1139: dataIn2 = 32'd0; 
32'd1140: dataIn2 = 32'd1; 
32'd1141: dataIn2 = 32'd1; 
32'd1142: dataIn2 = 32'd0; 
32'd1143: dataIn2 = 32'd1; 
32'd1144: dataIn2 = 32'd0; 
32'd1145: dataIn2 = 32'd0; 
32'd1146: dataIn2 = 32'd1; 
32'd1147: dataIn2 = 32'd0; 
32'd1148: dataIn2 = 32'd1; 
32'd1149: dataIn2 = 32'd1; 
32'd1150: dataIn2 = 32'd1; 
32'd1151: dataIn2 = 32'd0; 
32'd1152: dataIn2 = 32'd1; 
32'd1153: dataIn2 = 32'd0; 
32'd1154: dataIn2 = 32'd1; 
32'd1155: dataIn2 = 32'd1; 
32'd1156: dataIn2 = 32'd1; 
32'd1157: dataIn2 = 32'd0; 
32'd1158: dataIn2 = 32'd1; 
32'd1159: dataIn2 = 32'd1; 
32'd1160: dataIn2 = 32'd0; 
32'd1161: dataIn2 = 32'd0; 
32'd1162: dataIn2 = 32'd1; 
32'd1163: dataIn2 = 32'd1; 
32'd1164: dataIn2 = 32'd0; 
32'd1165: dataIn2 = 32'd0; 
32'd1166: dataIn2 = 32'd0; 
32'd1167: dataIn2 = 32'd1; 
32'd1168: dataIn2 = 32'd1; 
32'd1169: dataIn2 = 32'd0; 
32'd1170: dataIn2 = 32'd0; 
32'd1171: dataIn2 = 32'd0; 
32'd1172: dataIn2 = 32'd0; 
32'd1173: dataIn2 = 32'd0; 
32'd1174: dataIn2 = 32'd0; 
32'd1175: dataIn2 = 32'd1; 
32'd1176: dataIn2 = 32'd0; 
32'd1177: dataIn2 = 32'd0; 
32'd1178: dataIn2 = 32'd1; 
32'd1179: dataIn2 = 32'd0; 
32'd1180: dataIn2 = 32'd0; 
32'd1181: dataIn2 = 32'd0; 
32'd1182: dataIn2 = 32'd0; 
32'd1183: dataIn2 = 32'd0; 
32'd1184: dataIn2 = 32'd0; 
32'd1185: dataIn2 = 32'd0; 
32'd1186: dataIn2 = 32'd0; 
32'd1187: dataIn2 = 32'd0; 
32'd1188: dataIn2 = 32'd1; 
32'd1189: dataIn2 = 32'd1; 
32'd1190: dataIn2 = 32'd1; 
32'd1191: dataIn2 = 32'd0; 
32'd1192: dataIn2 = 32'd1; 
32'd1193: dataIn2 = 32'd0; 
32'd1194: dataIn2 = 32'd1; 
32'd1195: dataIn2 = 32'd0; 
32'd1196: dataIn2 = 32'd0; 
32'd1197: dataIn2 = 32'd1; 
32'd1198: dataIn2 = 32'd0; 
32'd1199: dataIn2 = 32'd0; 
32'd1200: dataIn2 = 32'd0; 
32'd1201: dataIn2 = 32'd1; 
32'd1202: dataIn2 = 32'd0; 
32'd1203: dataIn2 = 32'd1; 
32'd1204: dataIn2 = 32'd0; 
32'd1205: dataIn2 = 32'd1; 
32'd1206: dataIn2 = 32'd0; 
32'd1207: dataIn2 = 32'd0; 
32'd1208: dataIn2 = 32'd0; 
32'd1209: dataIn2 = 32'd1; 
32'd1210: dataIn2 = 32'd1; 
32'd1211: dataIn2 = 32'd1; 
32'd1212: dataIn2 = 32'd1; 
32'd1213: dataIn2 = 32'd0; 
32'd1214: dataIn2 = 32'd1; 
32'd1215: dataIn2 = 32'd0; 
32'd1216: dataIn2 = 32'd0; 
32'd1217: dataIn2 = 32'd0; 
32'd1218: dataIn2 = 32'd0; 
32'd1219: dataIn2 = 32'd1; 
32'd1220: dataIn2 = 32'd1; 
32'd1221: dataIn2 = 32'd0; 
32'd1222: dataIn2 = 32'd0; 
32'd1223: dataIn2 = 32'd0; 
32'd1224: dataIn2 = 32'd0; 
32'd1225: dataIn2 = 32'd1; 
32'd1226: dataIn2 = 32'd0; 
32'd1227: dataIn2 = 32'd0; 
32'd1228: dataIn2 = 32'd1; 
32'd1229: dataIn2 = 32'd0; 
32'd1230: dataIn2 = 32'd1; 
32'd1231: dataIn2 = 32'd0; 
32'd1232: dataIn2 = 32'd0; 
32'd1233: dataIn2 = 32'd0; 
32'd1234: dataIn2 = 32'd1; 
32'd1235: dataIn2 = 32'd0; 
32'd1236: dataIn2 = 32'd0; 
32'd1237: dataIn2 = 32'd0; 
32'd1238: dataIn2 = 32'd0; 
32'd1239: dataIn2 = 32'd1; 
32'd1240: dataIn2 = 32'd0; 
32'd1241: dataIn2 = 32'd1; 
32'd1242: dataIn2 = 32'd0; 
32'd1243: dataIn2 = 32'd0; 
32'd1244: dataIn2 = 32'd0; 
32'd1245: dataIn2 = 32'd0; 
32'd1246: dataIn2 = 32'd1; 
32'd1247: dataIn2 = 32'd0; 
32'd1248: dataIn2 = 32'd0; 
32'd1249: dataIn2 = 32'd1; 
32'd1250: dataIn2 = 32'd1; 
32'd1251: dataIn2 = 32'd0; 
32'd1252: dataIn2 = 32'd0; 
32'd1253: dataIn2 = 32'd1; 
32'd1254: dataIn2 = 32'd0; 
32'd1255: dataIn2 = 32'd0; 
32'd1256: dataIn2 = 32'd0; 
32'd1257: dataIn2 = 32'd0; 
32'd1258: dataIn2 = 32'd1; 
32'd1259: dataIn2 = 32'd0; 
32'd1260: dataIn2 = 32'd0; 
32'd1261: dataIn2 = 32'd0; 
32'd1262: dataIn2 = 32'd1; 
32'd1263: dataIn2 = 32'd1; 
32'd1264: dataIn2 = 32'd0; 
32'd1265: dataIn2 = 32'd0; 
32'd1266: dataIn2 = 32'd1; 
32'd1267: dataIn2 = 32'd1; 
32'd1268: dataIn2 = 32'd1; 
32'd1269: dataIn2 = 32'd0; 
32'd1270: dataIn2 = 32'd0; 
32'd1271: dataIn2 = 32'd1; 
32'd1272: dataIn2 = 32'd0; 
32'd1273: dataIn2 = 32'd0; 
32'd1274: dataIn2 = 32'd1; 
32'd1275: dataIn2 = 32'd1; 
32'd1276: dataIn2 = 32'd1; 
32'd1277: dataIn2 = 32'd0; 
32'd1278: dataIn2 = 32'd0; 
32'd1279: dataIn2 = 32'd1; 
32'd1280: dataIn2 = 32'd1; 
32'd1281: dataIn2 = 32'd1; 
32'd1282: dataIn2 = 32'd0; 
32'd1283: dataIn2 = 32'd1; 
32'd1284: dataIn2 = 32'd1; 
32'd1285: dataIn2 = 32'd1; 
32'd1286: dataIn2 = 32'd0; 
32'd1287: dataIn2 = 32'd0; 
32'd1288: dataIn2 = 32'd1; 
32'd1289: dataIn2 = 32'd1; 
32'd1290: dataIn2 = 32'd1; 
32'd1291: dataIn2 = 32'd1; 
32'd1292: dataIn2 = 32'd0; 
32'd1293: dataIn2 = 32'd1; 
32'd1294: dataIn2 = 32'd0; 
32'd1295: dataIn2 = 32'd1; 
32'd1296: dataIn2 = 32'd0; 
32'd1297: dataIn2 = 32'd0; 
32'd1298: dataIn2 = 32'd1; 
32'd1299: dataIn2 = 32'd0; 
32'd1300: dataIn2 = 32'd1; 
32'd1301: dataIn2 = 32'd1; 
32'd1302: dataIn2 = 32'd0; 
32'd1303: dataIn2 = 32'd0; 
32'd1304: dataIn2 = 32'd1; 
32'd1305: dataIn2 = 32'd1; 
32'd1306: dataIn2 = 32'd0; 
32'd1307: dataIn2 = 32'd0; 
32'd1308: dataIn2 = 32'd1; 
32'd1309: dataIn2 = 32'd0; 
32'd1310: dataIn2 = 32'd1; 
32'd1311: dataIn2 = 32'd0; 
32'd1312: dataIn2 = 32'd0; 
32'd1313: dataIn2 = 32'd0; 
32'd1314: dataIn2 = 32'd0; 
32'd1315: dataIn2 = 32'd0; 
32'd1316: dataIn2 = 32'd1; 
32'd1317: dataIn2 = 32'd1; 
32'd1318: dataIn2 = 32'd0; 
32'd1319: dataIn2 = 32'd0; 
32'd1320: dataIn2 = 32'd0; 
32'd1321: dataIn2 = 32'd1; 
32'd1322: dataIn2 = 32'd1; 
32'd1323: dataIn2 = 32'd0; 
32'd1324: dataIn2 = 32'd1; 
32'd1325: dataIn2 = 32'd1; 
32'd1326: dataIn2 = 32'd0; 
32'd1327: dataIn2 = 32'd1; 
32'd1328: dataIn2 = 32'd1; 
32'd1329: dataIn2 = 32'd1; 
32'd1330: dataIn2 = 32'd1; 
32'd1331: dataIn2 = 32'd1; 
32'd1332: dataIn2 = 32'd1; 
32'd1333: dataIn2 = 32'd0; 
32'd1334: dataIn2 = 32'd0; 
32'd1335: dataIn2 = 32'd0; 
32'd1336: dataIn2 = 32'd1; 
32'd1337: dataIn2 = 32'd1; 
32'd1338: dataIn2 = 32'd1; 
32'd1339: dataIn2 = 32'd0; 
32'd1340: dataIn2 = 32'd1; 
32'd1341: dataIn2 = 32'd1; 
32'd1342: dataIn2 = 32'd0; 
32'd1343: dataIn2 = 32'd0; 
32'd1344: dataIn2 = 32'd0; 
32'd1345: dataIn2 = 32'd0; 
32'd1346: dataIn2 = 32'd0; 
32'd1347: dataIn2 = 32'd1; 
32'd1348: dataIn2 = 32'd1; 
32'd1349: dataIn2 = 32'd0; 
32'd1350: dataIn2 = 32'd1; 
32'd1351: dataIn2 = 32'd1; 
32'd1352: dataIn2 = 32'd0; 
32'd1353: dataIn2 = 32'd0; 
32'd1354: dataIn2 = 32'd1; 
32'd1355: dataIn2 = 32'd0; 
32'd1356: dataIn2 = 32'd0; 
32'd1357: dataIn2 = 32'd1; 
32'd1358: dataIn2 = 32'd0; 
32'd1359: dataIn2 = 32'd0; 
32'd1360: dataIn2 = 32'd0; 
32'd1361: dataIn2 = 32'd0; 
32'd1362: dataIn2 = 32'd0; 
32'd1363: dataIn2 = 32'd1; 
32'd1364: dataIn2 = 32'd1; 
32'd1365: dataIn2 = 32'd1; 
32'd1366: dataIn2 = 32'd1; 
32'd1367: dataIn2 = 32'd0; 
32'd1368: dataIn2 = 32'd1; 
32'd1369: dataIn2 = 32'd1; 
32'd1370: dataIn2 = 32'd0; 
32'd1371: dataIn2 = 32'd1; 
32'd1372: dataIn2 = 32'd1; 
32'd1373: dataIn2 = 32'd1; 
32'd1374: dataIn2 = 32'd1; 
32'd1375: dataIn2 = 32'd0; 
32'd1376: dataIn2 = 32'd1; 
32'd1377: dataIn2 = 32'd0; 
32'd1378: dataIn2 = 32'd0; 
32'd1379: dataIn2 = 32'd0; 
32'd1380: dataIn2 = 32'd0; 
32'd1381: dataIn2 = 32'd0; 
32'd1382: dataIn2 = 32'd0; 
32'd1383: dataIn2 = 32'd1; 
32'd1384: dataIn2 = 32'd1; 
32'd1385: dataIn2 = 32'd1; 
32'd1386: dataIn2 = 32'd1; 
32'd1387: dataIn2 = 32'd1; 
32'd1388: dataIn2 = 32'd0; 
32'd1389: dataIn2 = 32'd1; 
32'd1390: dataIn2 = 32'd0; 
32'd1391: dataIn2 = 32'd0; 
32'd1392: dataIn2 = 32'd0; 
32'd1393: dataIn2 = 32'd1; 
32'd1394: dataIn2 = 32'd1; 
32'd1395: dataIn2 = 32'd0; 
32'd1396: dataIn2 = 32'd0; 
32'd1397: dataIn2 = 32'd1; 
32'd1398: dataIn2 = 32'd1; 
32'd1399: dataIn2 = 32'd1; 
32'd1400: dataIn2 = 32'd0; 
32'd1401: dataIn2 = 32'd0; 
32'd1402: dataIn2 = 32'd1; 
32'd1403: dataIn2 = 32'd1; 
32'd1404: dataIn2 = 32'd0; 
32'd1405: dataIn2 = 32'd0; 
32'd1406: dataIn2 = 32'd1; 
32'd1407: dataIn2 = 32'd1; 
32'd1408: dataIn2 = 32'd0; 
32'd1409: dataIn2 = 32'd0; 
32'd1410: dataIn2 = 32'd1; 
32'd1411: dataIn2 = 32'd0; 
32'd1412: dataIn2 = 32'd0; 
32'd1413: dataIn2 = 32'd1; 
32'd1414: dataIn2 = 32'd0; 
32'd1415: dataIn2 = 32'd1; 
32'd1416: dataIn2 = 32'd0; 
32'd1417: dataIn2 = 32'd0; 
32'd1418: dataIn2 = 32'd1; 
32'd1419: dataIn2 = 32'd0; 
32'd1420: dataIn2 = 32'd0; 
32'd1421: dataIn2 = 32'd0; 
32'd1422: dataIn2 = 32'd1; 
32'd1423: dataIn2 = 32'd1; 
32'd1424: dataIn2 = 32'd1; 
32'd1425: dataIn2 = 32'd0; 
32'd1426: dataIn2 = 32'd1; 
32'd1427: dataIn2 = 32'd1; 
32'd1428: dataIn2 = 32'd1; 
32'd1429: dataIn2 = 32'd1; 
32'd1430: dataIn2 = 32'd1; 
32'd1431: dataIn2 = 32'd1; 
32'd1432: dataIn2 = 32'd1; 
32'd1433: dataIn2 = 32'd0; 
32'd1434: dataIn2 = 32'd1; 
32'd1435: dataIn2 = 32'd0; 
32'd1436: dataIn2 = 32'd1; 
32'd1437: dataIn2 = 32'd1; 
32'd1438: dataIn2 = 32'd0; 
32'd1439: dataIn2 = 32'd1; 
32'd1440: dataIn2 = 32'd1; 
32'd1441: dataIn2 = 32'd1; 
32'd1442: dataIn2 = 32'd1; 
32'd1443: dataIn2 = 32'd1; 
32'd1444: dataIn2 = 32'd0; 
32'd1445: dataIn2 = 32'd0; 
32'd1446: dataIn2 = 32'd0; 
32'd1447: dataIn2 = 32'd0; 
32'd1448: dataIn2 = 32'd0; 
32'd1449: dataIn2 = 32'd0; 
32'd1450: dataIn2 = 32'd1; 
32'd1451: dataIn2 = 32'd0; 
32'd1452: dataIn2 = 32'd1; 
32'd1453: dataIn2 = 32'd1; 
32'd1454: dataIn2 = 32'd0; 
32'd1455: dataIn2 = 32'd1; 
32'd1456: dataIn2 = 32'd0; 
32'd1457: dataIn2 = 32'd1; 
32'd1458: dataIn2 = 32'd0; 
32'd1459: dataIn2 = 32'd1; 
32'd1460: dataIn2 = 32'd1; 
32'd1461: dataIn2 = 32'd1; 
32'd1462: dataIn2 = 32'd0; 
32'd1463: dataIn2 = 32'd1; 
32'd1464: dataIn2 = 32'd0; 
32'd1465: dataIn2 = 32'd0; 
32'd1466: dataIn2 = 32'd0; 
32'd1467: dataIn2 = 32'd1; 
32'd1468: dataIn2 = 32'd0; 
32'd1469: dataIn2 = 32'd0; 
32'd1470: dataIn2 = 32'd0; 
32'd1471: dataIn2 = 32'd0; 
32'd1472: dataIn2 = 32'd1; 
32'd1473: dataIn2 = 32'd1; 
32'd1474: dataIn2 = 32'd0; 
32'd1475: dataIn2 = 32'd0; 
32'd1476: dataIn2 = 32'd0; 
32'd1477: dataIn2 = 32'd0; 
32'd1478: dataIn2 = 32'd0; 
32'd1479: dataIn2 = 32'd0; 
32'd1480: dataIn2 = 32'd0; 
32'd1481: dataIn2 = 32'd1; 
32'd1482: dataIn2 = 32'd1; 
32'd1483: dataIn2 = 32'd1; 
32'd1484: dataIn2 = 32'd1; 
32'd1485: dataIn2 = 32'd0; 
32'd1486: dataIn2 = 32'd1; 
32'd1487: dataIn2 = 32'd0; 
32'd1488: dataIn2 = 32'd1; 
32'd1489: dataIn2 = 32'd1; 
32'd1490: dataIn2 = 32'd0; 
32'd1491: dataIn2 = 32'd0; 
32'd1492: dataIn2 = 32'd1; 
32'd1493: dataIn2 = 32'd1; 
32'd1494: dataIn2 = 32'd0; 
32'd1495: dataIn2 = 32'd0; 
32'd1496: dataIn2 = 32'd1; 
32'd1497: dataIn2 = 32'd0; 
32'd1498: dataIn2 = 32'd1; 
32'd1499: dataIn2 = 32'd1; 
32'd1500: dataIn2 = 32'd0; 
32'd1501: dataIn2 = 32'd0; 
32'd1502: dataIn2 = 32'd0; 
32'd1503: dataIn2 = 32'd0; 
32'd1504: dataIn2 = 32'd0; 
32'd1505: dataIn2 = 32'd0; 
32'd1506: dataIn2 = 32'd0; 
32'd1507: dataIn2 = 32'd0; 
32'd1508: dataIn2 = 32'd0; 
32'd1509: dataIn2 = 32'd0; 
32'd1510: dataIn2 = 32'd1; 
32'd1511: dataIn2 = 32'd0; 
32'd1512: dataIn2 = 32'd1; 
32'd1513: dataIn2 = 32'd1; 
32'd1514: dataIn2 = 32'd0; 
32'd1515: dataIn2 = 32'd0; 
32'd1516: dataIn2 = 32'd0; 
32'd1517: dataIn2 = 32'd0; 
32'd1518: dataIn2 = 32'd0; 
32'd1519: dataIn2 = 32'd0; 
32'd1520: dataIn2 = 32'd1; 
32'd1521: dataIn2 = 32'd0; 
32'd1522: dataIn2 = 32'd0; 
32'd1523: dataIn2 = 32'd1; 
32'd1524: dataIn2 = 32'd1; 
32'd1525: dataIn2 = 32'd1; 
32'd1526: dataIn2 = 32'd0; 
32'd1527: dataIn2 = 32'd0; 
32'd1528: dataIn2 = 32'd0; 
32'd1529: dataIn2 = 32'd1; 
32'd1530: dataIn2 = 32'd0; 
32'd1531: dataIn2 = 32'd1; 
32'd1532: dataIn2 = 32'd1; 
32'd1533: dataIn2 = 32'd0; 
32'd1534: dataIn2 = 32'd0; 
32'd1535: dataIn2 = 32'd0; 
32'd1536: dataIn2 = 32'd1; 
32'd1537: dataIn2 = 32'd1; 
32'd1538: dataIn2 = 32'd1; 
32'd1539: dataIn2 = 32'd1; 
32'd1540: dataIn2 = 32'd0; 
32'd1541: dataIn2 = 32'd0; 
32'd1542: dataIn2 = 32'd0; 
32'd1543: dataIn2 = 32'd1; 
32'd1544: dataIn2 = 32'd0; 
32'd1545: dataIn2 = 32'd1; 
32'd1546: dataIn2 = 32'd1; 
32'd1547: dataIn2 = 32'd1; 
32'd1548: dataIn2 = 32'd1; 
32'd1549: dataIn2 = 32'd0; 
32'd1550: dataIn2 = 32'd1; 
32'd1551: dataIn2 = 32'd1; 
32'd1552: dataIn2 = 32'd1; 
32'd1553: dataIn2 = 32'd0; 
32'd1554: dataIn2 = 32'd0; 
32'd1555: dataIn2 = 32'd0; 
32'd1556: dataIn2 = 32'd0; 
32'd1557: dataIn2 = 32'd1; 
32'd1558: dataIn2 = 32'd1; 
32'd1559: dataIn2 = 32'd1; 
32'd1560: dataIn2 = 32'd0; 
32'd1561: dataIn2 = 32'd0; 
32'd1562: dataIn2 = 32'd1; 
32'd1563: dataIn2 = 32'd1; 
32'd1564: dataIn2 = 32'd1; 
32'd1565: dataIn2 = 32'd1; 
32'd1566: dataIn2 = 32'd0; 
32'd1567: dataIn2 = 32'd1; 
32'd1568: dataIn2 = 32'd0; 
32'd1569: dataIn2 = 32'd0; 
32'd1570: dataIn2 = 32'd0; 
32'd1571: dataIn2 = 32'd0; 
32'd1572: dataIn2 = 32'd1; 
32'd1573: dataIn2 = 32'd1; 
32'd1574: dataIn2 = 32'd0; 
32'd1575: dataIn2 = 32'd1; 
32'd1576: dataIn2 = 32'd1; 
32'd1577: dataIn2 = 32'd1; 
32'd1578: dataIn2 = 32'd1; 
32'd1579: dataIn2 = 32'd0; 
32'd1580: dataIn2 = 32'd0; 
32'd1581: dataIn2 = 32'd0; 
32'd1582: dataIn2 = 32'd0; 
32'd1583: dataIn2 = 32'd1; 
32'd1584: dataIn2 = 32'd0; 
32'd1585: dataIn2 = 32'd1; 
32'd1586: dataIn2 = 32'd0; 
32'd1587: dataIn2 = 32'd1; 
32'd1588: dataIn2 = 32'd1; 
32'd1589: dataIn2 = 32'd0; 
32'd1590: dataIn2 = 32'd0; 
32'd1591: dataIn2 = 32'd1; 
32'd1592: dataIn2 = 32'd1; 
32'd1593: dataIn2 = 32'd1; 
32'd1594: dataIn2 = 32'd0; 
32'd1595: dataIn2 = 32'd0; 
32'd1596: dataIn2 = 32'd1; 
32'd1597: dataIn2 = 32'd0; 
32'd1598: dataIn2 = 32'd0; 
32'd1599: dataIn2 = 32'd1; 
32'd1600: dataIn2 = 32'd1; 
32'd1601: dataIn2 = 32'd0; 
32'd1602: dataIn2 = 32'd1; 
32'd1603: dataIn2 = 32'd0; 
32'd1604: dataIn2 = 32'd1; 
32'd1605: dataIn2 = 32'd1; 
32'd1606: dataIn2 = 32'd0; 
32'd1607: dataIn2 = 32'd1; 
32'd1608: dataIn2 = 32'd0; 
32'd1609: dataIn2 = 32'd1; 
32'd1610: dataIn2 = 32'd0; 
32'd1611: dataIn2 = 32'd0; 
32'd1612: dataIn2 = 32'd1; 
32'd1613: dataIn2 = 32'd1; 
32'd1614: dataIn2 = 32'd1; 
32'd1615: dataIn2 = 32'd1; 
32'd1616: dataIn2 = 32'd0; 
32'd1617: dataIn2 = 32'd1; 
32'd1618: dataIn2 = 32'd1; 
32'd1619: dataIn2 = 32'd1; 
32'd1620: dataIn2 = 32'd1; 
32'd1621: dataIn2 = 32'd0; 
32'd1622: dataIn2 = 32'd0; 
32'd1623: dataIn2 = 32'd1; 
32'd1624: dataIn2 = 32'd1; 
32'd1625: dataIn2 = 32'd0; 
32'd1626: dataIn2 = 32'd0; 
32'd1627: dataIn2 = 32'd1; 
32'd1628: dataIn2 = 32'd0; 
32'd1629: dataIn2 = 32'd0; 
32'd1630: dataIn2 = 32'd0; 
32'd1631: dataIn2 = 32'd1; 
32'd1632: dataIn2 = 32'd1; 
32'd1633: dataIn2 = 32'd0; 
32'd1634: dataIn2 = 32'd1; 
32'd1635: dataIn2 = 32'd0; 
32'd1636: dataIn2 = 32'd0; 
32'd1637: dataIn2 = 32'd0; 
32'd1638: dataIn2 = 32'd0; 
32'd1639: dataIn2 = 32'd1; 
32'd1640: dataIn2 = 32'd0; 
32'd1641: dataIn2 = 32'd0; 
32'd1642: dataIn2 = 32'd1; 
32'd1643: dataIn2 = 32'd1; 
32'd1644: dataIn2 = 32'd0; 
32'd1645: dataIn2 = 32'd1; 
32'd1646: dataIn2 = 32'd0; 
32'd1647: dataIn2 = 32'd1; 
32'd1648: dataIn2 = 32'd1; 
32'd1649: dataIn2 = 32'd0; 
32'd1650: dataIn2 = 32'd0; 
32'd1651: dataIn2 = 32'd0; 
32'd1652: dataIn2 = 32'd0; 
32'd1653: dataIn2 = 32'd0; 
32'd1654: dataIn2 = 32'd0; 
32'd1655: dataIn2 = 32'd0; 
32'd1656: dataIn2 = 32'd1; 
32'd1657: dataIn2 = 32'd0; 
32'd1658: dataIn2 = 32'd0; 
32'd1659: dataIn2 = 32'd0; 
32'd1660: dataIn2 = 32'd1; 
32'd1661: dataIn2 = 32'd0; 
32'd1662: dataIn2 = 32'd1; 
32'd1663: dataIn2 = 32'd1; 
32'd1664: dataIn2 = 32'd1; 
32'd1665: dataIn2 = 32'd1; 
32'd1666: dataIn2 = 32'd1; 
32'd1667: dataIn2 = 32'd0; 
32'd1668: dataIn2 = 32'd0; 
32'd1669: dataIn2 = 32'd1; 
32'd1670: dataIn2 = 32'd0; 
32'd1671: dataIn2 = 32'd1; 
32'd1672: dataIn2 = 32'd0; 
32'd1673: dataIn2 = 32'd1; 
32'd1674: dataIn2 = 32'd0; 
32'd1675: dataIn2 = 32'd1; 
32'd1676: dataIn2 = 32'd0; 
32'd1677: dataIn2 = 32'd0; 
32'd1678: dataIn2 = 32'd0; 
32'd1679: dataIn2 = 32'd1; 
32'd1680: dataIn2 = 32'd0; 
32'd1681: dataIn2 = 32'd1; 
32'd1682: dataIn2 = 32'd1; 
32'd1683: dataIn2 = 32'd1; 
32'd1684: dataIn2 = 32'd1; 
32'd1685: dataIn2 = 32'd1; 
32'd1686: dataIn2 = 32'd1; 
32'd1687: dataIn2 = 32'd1; 
32'd1688: dataIn2 = 32'd0; 
32'd1689: dataIn2 = 32'd0; 
32'd1690: dataIn2 = 32'd0; 
32'd1691: dataIn2 = 32'd1; 
32'd1692: dataIn2 = 32'd1; 
32'd1693: dataIn2 = 32'd1; 
32'd1694: dataIn2 = 32'd0; 
32'd1695: dataIn2 = 32'd1; 
32'd1696: dataIn2 = 32'd0; 
32'd1697: dataIn2 = 32'd0; 
32'd1698: dataIn2 = 32'd1; 
32'd1699: dataIn2 = 32'd1; 
32'd1700: dataIn2 = 32'd1; 
32'd1701: dataIn2 = 32'd1; 
32'd1702: dataIn2 = 32'd1; 
32'd1703: dataIn2 = 32'd0; 
32'd1704: dataIn2 = 32'd1; 
32'd1705: dataIn2 = 32'd0; 
32'd1706: dataIn2 = 32'd1; 
32'd1707: dataIn2 = 32'd0; 
32'd1708: dataIn2 = 32'd0; 
32'd1709: dataIn2 = 32'd0; 
32'd1710: dataIn2 = 32'd0; 
32'd1711: dataIn2 = 32'd1; 
32'd1712: dataIn2 = 32'd1; 
32'd1713: dataIn2 = 32'd1; 
32'd1714: dataIn2 = 32'd0; 
32'd1715: dataIn2 = 32'd0; 
32'd1716: dataIn2 = 32'd0; 
32'd1717: dataIn2 = 32'd1; 
32'd1718: dataIn2 = 32'd0; 
32'd1719: dataIn2 = 32'd1; 
32'd1720: dataIn2 = 32'd1; 
32'd1721: dataIn2 = 32'd0; 
32'd1722: dataIn2 = 32'd0; 
32'd1723: dataIn2 = 32'd0; 
32'd1724: dataIn2 = 32'd0; 
32'd1725: dataIn2 = 32'd1; 
32'd1726: dataIn2 = 32'd0; 
32'd1727: dataIn2 = 32'd1; 
32'd1728: dataIn2 = 32'd0; 
32'd1729: dataIn2 = 32'd1; 
32'd1730: dataIn2 = 32'd0; 
32'd1731: dataIn2 = 32'd1; 
32'd1732: dataIn2 = 32'd0; 
32'd1733: dataIn2 = 32'd1; 
32'd1734: dataIn2 = 32'd0; 
32'd1735: dataIn2 = 32'd1; 
32'd1736: dataIn2 = 32'd1; 
32'd1737: dataIn2 = 32'd1; 
32'd1738: dataIn2 = 32'd0; 
32'd1739: dataIn2 = 32'd1; 
32'd1740: dataIn2 = 32'd1; 
32'd1741: dataIn2 = 32'd0; 
32'd1742: dataIn2 = 32'd0; 
32'd1743: dataIn2 = 32'd1; 
32'd1744: dataIn2 = 32'd1; 
32'd1745: dataIn2 = 32'd1; 
32'd1746: dataIn2 = 32'd1; 
32'd1747: dataIn2 = 32'd1; 
32'd1748: dataIn2 = 32'd0; 
32'd1749: dataIn2 = 32'd1; 
32'd1750: dataIn2 = 32'd0; 
32'd1751: dataIn2 = 32'd1; 
32'd1752: dataIn2 = 32'd1; 
32'd1753: dataIn2 = 32'd0; 
32'd1754: dataIn2 = 32'd0; 
32'd1755: dataIn2 = 32'd0; 
32'd1756: dataIn2 = 32'd0; 
32'd1757: dataIn2 = 32'd0; 
32'd1758: dataIn2 = 32'd1; 
32'd1759: dataIn2 = 32'd1; 
32'd1760: dataIn2 = 32'd1; 
32'd1761: dataIn2 = 32'd1; 
32'd1762: dataIn2 = 32'd1; 
32'd1763: dataIn2 = 32'd1; 
32'd1764: dataIn2 = 32'd1; 
32'd1765: dataIn2 = 32'd1; 
32'd1766: dataIn2 = 32'd0; 
32'd1767: dataIn2 = 32'd1; 
32'd1768: dataIn2 = 32'd0; 
32'd1769: dataIn2 = 32'd0; 
32'd1770: dataIn2 = 32'd0; 
32'd1771: dataIn2 = 32'd1; 
32'd1772: dataIn2 = 32'd0; 
32'd1773: dataIn2 = 32'd0; 
32'd1774: dataIn2 = 32'd0; 
32'd1775: dataIn2 = 32'd0; 
32'd1776: dataIn2 = 32'd0; 
32'd1777: dataIn2 = 32'd0; 
32'd1778: dataIn2 = 32'd0; 
32'd1779: dataIn2 = 32'd1; 
32'd1780: dataIn2 = 32'd1; 
32'd1781: dataIn2 = 32'd0; 
32'd1782: dataIn2 = 32'd1; 
32'd1783: dataIn2 = 32'd1; 
32'd1784: dataIn2 = 32'd0; 
32'd1785: dataIn2 = 32'd1; 
32'd1786: dataIn2 = 32'd0; 
32'd1787: dataIn2 = 32'd0; 
32'd1788: dataIn2 = 32'd0; 
32'd1789: dataIn2 = 32'd0; 
32'd1790: dataIn2 = 32'd0; 
32'd1791: dataIn2 = 32'd0; 
32'd1792: dataIn2 = 32'd1; 
32'd1793: dataIn2 = 32'd0; 
32'd1794: dataIn2 = 32'd1; 
32'd1795: dataIn2 = 32'd1; 
32'd1796: dataIn2 = 32'd0; 
32'd1797: dataIn2 = 32'd0; 
32'd1798: dataIn2 = 32'd1; 
32'd1799: dataIn2 = 32'd1; 
32'd1800: dataIn2 = 32'd1; 
32'd1801: dataIn2 = 32'd1; 
32'd1802: dataIn2 = 32'd0; 
32'd1803: dataIn2 = 32'd0; 
32'd1804: dataIn2 = 32'd1; 
32'd1805: dataIn2 = 32'd1; 
32'd1806: dataIn2 = 32'd1; 
32'd1807: dataIn2 = 32'd1; 
32'd1808: dataIn2 = 32'd1; 
32'd1809: dataIn2 = 32'd0; 
32'd1810: dataIn2 = 32'd1; 
32'd1811: dataIn2 = 32'd1; 
32'd1812: dataIn2 = 32'd1; 
32'd1813: dataIn2 = 32'd0; 
32'd1814: dataIn2 = 32'd0; 
32'd1815: dataIn2 = 32'd1; 
32'd1816: dataIn2 = 32'd1; 
32'd1817: dataIn2 = 32'd0; 
32'd1818: dataIn2 = 32'd1; 
32'd1819: dataIn2 = 32'd1; 
32'd1820: dataIn2 = 32'd1; 
32'd1821: dataIn2 = 32'd1; 
32'd1822: dataIn2 = 32'd0; 
32'd1823: dataIn2 = 32'd1; 
32'd1824: dataIn2 = 32'd1; 
32'd1825: dataIn2 = 32'd1; 
32'd1826: dataIn2 = 32'd1; 
32'd1827: dataIn2 = 32'd1; 
32'd1828: dataIn2 = 32'd1; 
32'd1829: dataIn2 = 32'd1; 
32'd1830: dataIn2 = 32'd1; 
32'd1831: dataIn2 = 32'd1; 
32'd1832: dataIn2 = 32'd1; 
32'd1833: dataIn2 = 32'd1; 
32'd1834: dataIn2 = 32'd1; 
32'd1835: dataIn2 = 32'd1; 
32'd1836: dataIn2 = 32'd0; 
32'd1837: dataIn2 = 32'd0; 
32'd1838: dataIn2 = 32'd1; 
32'd1839: dataIn2 = 32'd0; 
32'd1840: dataIn2 = 32'd0; 
32'd1841: dataIn2 = 32'd1; 
32'd1842: dataIn2 = 32'd0; 
32'd1843: dataIn2 = 32'd0; 
32'd1844: dataIn2 = 32'd0; 
32'd1845: dataIn2 = 32'd0; 
32'd1846: dataIn2 = 32'd0; 
32'd1847: dataIn2 = 32'd1; 
32'd1848: dataIn2 = 32'd1; 
32'd1849: dataIn2 = 32'd1; 
32'd1850: dataIn2 = 32'd0; 
32'd1851: dataIn2 = 32'd0; 
32'd1852: dataIn2 = 32'd1; 
32'd1853: dataIn2 = 32'd1; 
32'd1854: dataIn2 = 32'd0; 
32'd1855: dataIn2 = 32'd0; 
32'd1856: dataIn2 = 32'd0; 
32'd1857: dataIn2 = 32'd0; 
32'd1858: dataIn2 = 32'd1; 
32'd1859: dataIn2 = 32'd0; 
32'd1860: dataIn2 = 32'd1; 
32'd1861: dataIn2 = 32'd1; 
32'd1862: dataIn2 = 32'd0; 
32'd1863: dataIn2 = 32'd0; 
32'd1864: dataIn2 = 32'd1; 
32'd1865: dataIn2 = 32'd1; 
32'd1866: dataIn2 = 32'd0; 
32'd1867: dataIn2 = 32'd1; 
32'd1868: dataIn2 = 32'd1; 
32'd1869: dataIn2 = 32'd0; 
32'd1870: dataIn2 = 32'd1; 
32'd1871: dataIn2 = 32'd1; 
32'd1872: dataIn2 = 32'd1; 
32'd1873: dataIn2 = 32'd0; 
32'd1874: dataIn2 = 32'd1; 
32'd1875: dataIn2 = 32'd1; 
32'd1876: dataIn2 = 32'd1; 
32'd1877: dataIn2 = 32'd1; 
32'd1878: dataIn2 = 32'd1; 
32'd1879: dataIn2 = 32'd1; 
32'd1880: dataIn2 = 32'd1; 
32'd1881: dataIn2 = 32'd1; 
32'd1882: dataIn2 = 32'd1; 
32'd1883: dataIn2 = 32'd1; 
32'd1884: dataIn2 = 32'd1; 
32'd1885: dataIn2 = 32'd1; 
32'd1886: dataIn2 = 32'd1; 
32'd1887: dataIn2 = 32'd1; 
32'd1888: dataIn2 = 32'd1; 
32'd1889: dataIn2 = 32'd1; 
32'd1890: dataIn2 = 32'd0; 
32'd1891: dataIn2 = 32'd0; 
32'd1892: dataIn2 = 32'd1; 
32'd1893: dataIn2 = 32'd0; 
32'd1894: dataIn2 = 32'd0; 
32'd1895: dataIn2 = 32'd1; 
32'd1896: dataIn2 = 32'd1; 
32'd1897: dataIn2 = 32'd1; 
32'd1898: dataIn2 = 32'd0; 
32'd1899: dataIn2 = 32'd1; 
32'd1900: dataIn2 = 32'd1; 
32'd1901: dataIn2 = 32'd0; 
32'd1902: dataIn2 = 32'd0; 
32'd1903: dataIn2 = 32'd1; 
32'd1904: dataIn2 = 32'd1; 
32'd1905: dataIn2 = 32'd0; 
32'd1906: dataIn2 = 32'd1; 
32'd1907: dataIn2 = 32'd0; 
32'd1908: dataIn2 = 32'd1; 
32'd1909: dataIn2 = 32'd1; 
32'd1910: dataIn2 = 32'd0; 
32'd1911: dataIn2 = 32'd0; 
32'd1912: dataIn2 = 32'd1; 
32'd1913: dataIn2 = 32'd1; 
32'd1914: dataIn2 = 32'd1; 
32'd1915: dataIn2 = 32'd1; 
32'd1916: dataIn2 = 32'd1; 
32'd1917: dataIn2 = 32'd0; 
32'd1918: dataIn2 = 32'd1; 
32'd1919: dataIn2 = 32'd1; 
32'd1920: dataIn2 = 32'd1; 
32'd1921: dataIn2 = 32'd1; 
32'd1922: dataIn2 = 32'd0; 
32'd1923: dataIn2 = 32'd1; 
32'd1924: dataIn2 = 32'd0; 
32'd1925: dataIn2 = 32'd1; 
32'd1926: dataIn2 = 32'd0; 
32'd1927: dataIn2 = 32'd0; 
32'd1928: dataIn2 = 32'd0; 
32'd1929: dataIn2 = 32'd0; 
32'd1930: dataIn2 = 32'd0; 
32'd1931: dataIn2 = 32'd0; 
32'd1932: dataIn2 = 32'd1; 
32'd1933: dataIn2 = 32'd0; 
32'd1934: dataIn2 = 32'd0; 
32'd1935: dataIn2 = 32'd0; 
32'd1936: dataIn2 = 32'd1; 
32'd1937: dataIn2 = 32'd0; 
32'd1938: dataIn2 = 32'd1; 
32'd1939: dataIn2 = 32'd0; 
32'd1940: dataIn2 = 32'd1; 
32'd1941: dataIn2 = 32'd0; 
32'd1942: dataIn2 = 32'd0; 
32'd1943: dataIn2 = 32'd0; 
32'd1944: dataIn2 = 32'd1; 
32'd1945: dataIn2 = 32'd0; 
32'd1946: dataIn2 = 32'd0; 
32'd1947: dataIn2 = 32'd0; 
32'd1948: dataIn2 = 32'd0; 
32'd1949: dataIn2 = 32'd1; 
32'd1950: dataIn2 = 32'd1; 
32'd1951: dataIn2 = 32'd1; 
32'd1952: dataIn2 = 32'd0; 
32'd1953: dataIn2 = 32'd0; 
32'd1954: dataIn2 = 32'd0; 
32'd1955: dataIn2 = 32'd0; 
32'd1956: dataIn2 = 32'd0; 
32'd1957: dataIn2 = 32'd0; 
32'd1958: dataIn2 = 32'd1; 
32'd1959: dataIn2 = 32'd0; 
32'd1960: dataIn2 = 32'd0; 
32'd1961: dataIn2 = 32'd1; 
32'd1962: dataIn2 = 32'd0; 
32'd1963: dataIn2 = 32'd1; 
32'd1964: dataIn2 = 32'd0; 
32'd1965: dataIn2 = 32'd0; 
32'd1966: dataIn2 = 32'd0; 
32'd1967: dataIn2 = 32'd0; 
32'd1968: dataIn2 = 32'd0; 
32'd1969: dataIn2 = 32'd1; 
32'd1970: dataIn2 = 32'd0; 
32'd1971: dataIn2 = 32'd0; 
32'd1972: dataIn2 = 32'd0; 
32'd1973: dataIn2 = 32'd0; 
32'd1974: dataIn2 = 32'd1; 
32'd1975: dataIn2 = 32'd0; 
32'd1976: dataIn2 = 32'd0; 
32'd1977: dataIn2 = 32'd1; 
32'd1978: dataIn2 = 32'd1; 
32'd1979: dataIn2 = 32'd0; 
32'd1980: dataIn2 = 32'd0; 
32'd1981: dataIn2 = 32'd1; 
32'd1982: dataIn2 = 32'd1; 
32'd1983: dataIn2 = 32'd1; 
32'd1984: dataIn2 = 32'd0; 
32'd1985: dataIn2 = 32'd0; 
32'd1986: dataIn2 = 32'd1; 
32'd1987: dataIn2 = 32'd1; 
32'd1988: dataIn2 = 32'd0; 
32'd1989: dataIn2 = 32'd0; 
32'd1990: dataIn2 = 32'd1; 
32'd1991: dataIn2 = 32'd1; 
32'd1992: dataIn2 = 32'd1; 
32'd1993: dataIn2 = 32'd1; 
32'd1994: dataIn2 = 32'd1; 
32'd1995: dataIn2 = 32'd1; 
32'd1996: dataIn2 = 32'd0; 
32'd1997: dataIn2 = 32'd0; 
32'd1998: dataIn2 = 32'd1; 
32'd1999: dataIn2 = 32'd1; 
32'd2000: dataIn2 = 32'd0; 
32'd2001: dataIn2 = 32'd1; 
32'd2002: dataIn2 = 32'd1; 
32'd2003: dataIn2 = 32'd0; 
32'd2004: dataIn2 = 32'd1; 
32'd2005: dataIn2 = 32'd1; 
32'd2006: dataIn2 = 32'd0; 
32'd2007: dataIn2 = 32'd1; 
32'd2008: dataIn2 = 32'd0; 
32'd2009: dataIn2 = 32'd0; 
32'd2010: dataIn2 = 32'd0; 
32'd2011: dataIn2 = 32'd1; 
32'd2012: dataIn2 = 32'd1; 
32'd2013: dataIn2 = 32'd1; 
32'd2014: dataIn2 = 32'd1; 
32'd2015: dataIn2 = 32'd0; 
32'd2016: dataIn2 = 32'd0; 
32'd2017: dataIn2 = 32'd1; 
32'd2018: dataIn2 = 32'd1; 
32'd2019: dataIn2 = 32'd0; 
32'd2020: dataIn2 = 32'd0; 
32'd2021: dataIn2 = 32'd1; 
32'd2022: dataIn2 = 32'd0; 
32'd2023: dataIn2 = 32'd0; 
32'd2024: dataIn2 = 32'd1; 
32'd2025: dataIn2 = 32'd1; 
32'd2026: dataIn2 = 32'd1; 
32'd2027: dataIn2 = 32'd0; 
32'd2028: dataIn2 = 32'd0; 
32'd2029: dataIn2 = 32'd1; 
32'd2030: dataIn2 = 32'd1; 
32'd2031: dataIn2 = 32'd1; 
32'd2032: dataIn2 = 32'd1; 
32'd2033: dataIn2 = 32'd1; 
32'd2034: dataIn2 = 32'd0; 
32'd2035: dataIn2 = 32'd1; 
32'd2036: dataIn2 = 32'd0; 
32'd2037: dataIn2 = 32'd0; 
32'd2038: dataIn2 = 32'd0; 
32'd2039: dataIn2 = 32'd1; 
32'd2040: dataIn2 = 32'd1; 
32'd2041: dataIn2 = 32'd1; 
32'd2042: dataIn2 = 32'd1; 
32'd2043: dataIn2 = 32'd0; 
32'd2044: dataIn2 = 32'd0; 
32'd2045: dataIn2 = 32'd0; 
32'd2046: dataIn2 = 32'd0; 
32'd2047: dataIn2 = 32'd0; 
32'd2048: dataIn2 = 32'd1; 
32'd2049: dataIn2 = 32'd1; 
32'd2050: dataIn2 = 32'd0; 
32'd2051: dataIn2 = 32'd1; 
32'd2052: dataIn2 = 32'd0; 
32'd2053: dataIn2 = 32'd1; 
32'd2054: dataIn2 = 32'd0; 
32'd2055: dataIn2 = 32'd0; 
32'd2056: dataIn2 = 32'd1; 
32'd2057: dataIn2 = 32'd1; 
32'd2058: dataIn2 = 32'd1; 
32'd2059: dataIn2 = 32'd0; 
32'd2060: dataIn2 = 32'd0; 
32'd2061: dataIn2 = 32'd1; 
32'd2062: dataIn2 = 32'd0; 
32'd2063: dataIn2 = 32'd1; 
32'd2064: dataIn2 = 32'd1; 
32'd2065: dataIn2 = 32'd0; 
32'd2066: dataIn2 = 32'd0; 
32'd2067: dataIn2 = 32'd0; 
32'd2068: dataIn2 = 32'd1; 
32'd2069: dataIn2 = 32'd0; 
32'd2070: dataIn2 = 32'd0; 
32'd2071: dataIn2 = 32'd1; 
32'd2072: dataIn2 = 32'd1; 
32'd2073: dataIn2 = 32'd0; 
32'd2074: dataIn2 = 32'd1; 
32'd2075: dataIn2 = 32'd0; 
32'd2076: dataIn2 = 32'd0; 
32'd2077: dataIn2 = 32'd1; 
32'd2078: dataIn2 = 32'd0; 
32'd2079: dataIn2 = 32'd0; 
32'd2080: dataIn2 = 32'd1; 
32'd2081: dataIn2 = 32'd0; 
32'd2082: dataIn2 = 32'd1; 
32'd2083: dataIn2 = 32'd1; 
32'd2084: dataIn2 = 32'd1; 
32'd2085: dataIn2 = 32'd1; 
32'd2086: dataIn2 = 32'd0; 
32'd2087: dataIn2 = 32'd1; 
32'd2088: dataIn2 = 32'd0; 
32'd2089: dataIn2 = 32'd0; 
32'd2090: dataIn2 = 32'd1; 
32'd2091: dataIn2 = 32'd0; 
32'd2092: dataIn2 = 32'd0; 
32'd2093: dataIn2 = 32'd1; 
32'd2094: dataIn2 = 32'd0; 
32'd2095: dataIn2 = 32'd0; 
32'd2096: dataIn2 = 32'd1; 
32'd2097: dataIn2 = 32'd1; 
32'd2098: dataIn2 = 32'd1; 
32'd2099: dataIn2 = 32'd0; 
32'd2100: dataIn2 = 32'd1; 
32'd2101: dataIn2 = 32'd1; 
32'd2102: dataIn2 = 32'd1; 
32'd2103: dataIn2 = 32'd1; 
32'd2104: dataIn2 = 32'd1; 
32'd2105: dataIn2 = 32'd1; 
32'd2106: dataIn2 = 32'd0; 
32'd2107: dataIn2 = 32'd1; 
32'd2108: dataIn2 = 32'd1; 
32'd2109: dataIn2 = 32'd0; 
32'd2110: dataIn2 = 32'd0; 
32'd2111: dataIn2 = 32'd1; 
32'd2112: dataIn2 = 32'd0; 
32'd2113: dataIn2 = 32'd1; 
32'd2114: dataIn2 = 32'd0; 
32'd2115: dataIn2 = 32'd0; 
32'd2116: dataIn2 = 32'd1; 
32'd2117: dataIn2 = 32'd1; 
32'd2118: dataIn2 = 32'd1; 
32'd2119: dataIn2 = 32'd0; 
32'd2120: dataIn2 = 32'd0; 
32'd2121: dataIn2 = 32'd0; 
32'd2122: dataIn2 = 32'd0; 
32'd2123: dataIn2 = 32'd0; 
32'd2124: dataIn2 = 32'd1; 
32'd2125: dataIn2 = 32'd0; 
32'd2126: dataIn2 = 32'd0; 
32'd2127: dataIn2 = 32'd1; 
32'd2128: dataIn2 = 32'd1; 
32'd2129: dataIn2 = 32'd0; 
32'd2130: dataIn2 = 32'd0; 
32'd2131: dataIn2 = 32'd1; 
32'd2132: dataIn2 = 32'd1; 
32'd2133: dataIn2 = 32'd0; 
32'd2134: dataIn2 = 32'd1; 
32'd2135: dataIn2 = 32'd1; 
32'd2136: dataIn2 = 32'd1; 
32'd2137: dataIn2 = 32'd1; 
32'd2138: dataIn2 = 32'd0; 
32'd2139: dataIn2 = 32'd1; 
32'd2140: dataIn2 = 32'd0; 
32'd2141: dataIn2 = 32'd1; 
32'd2142: dataIn2 = 32'd0; 
32'd2143: dataIn2 = 32'd1; 
32'd2144: dataIn2 = 32'd1; 
32'd2145: dataIn2 = 32'd1; 
32'd2146: dataIn2 = 32'd1; 
32'd2147: dataIn2 = 32'd0; 
32'd2148: dataIn2 = 32'd1; 
32'd2149: dataIn2 = 32'd0; 
32'd2150: dataIn2 = 32'd1; 
32'd2151: dataIn2 = 32'd1; 
32'd2152: dataIn2 = 32'd0; 
32'd2153: dataIn2 = 32'd0; 
32'd2154: dataIn2 = 32'd1; 
32'd2155: dataIn2 = 32'd0; 
32'd2156: dataIn2 = 32'd0; 
32'd2157: dataIn2 = 32'd0; 
32'd2158: dataIn2 = 32'd0; 
32'd2159: dataIn2 = 32'd0; 
32'd2160: dataIn2 = 32'd1; 
32'd2161: dataIn2 = 32'd0; 
32'd2162: dataIn2 = 32'd0; 
32'd2163: dataIn2 = 32'd1; 
32'd2164: dataIn2 = 32'd1; 
32'd2165: dataIn2 = 32'd1; 
32'd2166: dataIn2 = 32'd0; 
32'd2167: dataIn2 = 32'd1; 
32'd2168: dataIn2 = 32'd1; 
32'd2169: dataIn2 = 32'd1; 
32'd2170: dataIn2 = 32'd1; 
32'd2171: dataIn2 = 32'd0; 
32'd2172: dataIn2 = 32'd0; 
32'd2173: dataIn2 = 32'd1; 
32'd2174: dataIn2 = 32'd0; 
32'd2175: dataIn2 = 32'd1; 
32'd2176: dataIn2 = 32'd0; 
32'd2177: dataIn2 = 32'd0; 
32'd2178: dataIn2 = 32'd1; 
32'd2179: dataIn2 = 32'd1; 
32'd2180: dataIn2 = 32'd0; 
32'd2181: dataIn2 = 32'd0; 
32'd2182: dataIn2 = 32'd1; 
32'd2183: dataIn2 = 32'd0; 
32'd2184: dataIn2 = 32'd1; 
32'd2185: dataIn2 = 32'd0; 
32'd2186: dataIn2 = 32'd0; 
32'd2187: dataIn2 = 32'd0; 
32'd2188: dataIn2 = 32'd0; 
32'd2189: dataIn2 = 32'd0; 
32'd2190: dataIn2 = 32'd0; 
32'd2191: dataIn2 = 32'd1; 
32'd2192: dataIn2 = 32'd1; 
32'd2193: dataIn2 = 32'd0; 
32'd2194: dataIn2 = 32'd1; 
32'd2195: dataIn2 = 32'd0; 
32'd2196: dataIn2 = 32'd1; 
32'd2197: dataIn2 = 32'd0; 
32'd2198: dataIn2 = 32'd1; 
32'd2199: dataIn2 = 32'd0; 
32'd2200: dataIn2 = 32'd0; 
32'd2201: dataIn2 = 32'd1; 
32'd2202: dataIn2 = 32'd0; 
32'd2203: dataIn2 = 32'd1; 
32'd2204: dataIn2 = 32'd0; 
32'd2205: dataIn2 = 32'd1; 
32'd2206: dataIn2 = 32'd1; 
32'd2207: dataIn2 = 32'd0; 
32'd2208: dataIn2 = 32'd1; 
32'd2209: dataIn2 = 32'd0; 
32'd2210: dataIn2 = 32'd0; 
32'd2211: dataIn2 = 32'd0; 
32'd2212: dataIn2 = 32'd0; 
32'd2213: dataIn2 = 32'd0; 
32'd2214: dataIn2 = 32'd0; 
32'd2215: dataIn2 = 32'd0; 
32'd2216: dataIn2 = 32'd0; 
32'd2217: dataIn2 = 32'd1; 
32'd2218: dataIn2 = 32'd1; 
32'd2219: dataIn2 = 32'd0; 
32'd2220: dataIn2 = 32'd1; 
32'd2221: dataIn2 = 32'd0; 
32'd2222: dataIn2 = 32'd1; 
32'd2223: dataIn2 = 32'd1; 
32'd2224: dataIn2 = 32'd0; 
32'd2225: dataIn2 = 32'd1; 
32'd2226: dataIn2 = 32'd1; 
32'd2227: dataIn2 = 32'd0; 
32'd2228: dataIn2 = 32'd0; 
32'd2229: dataIn2 = 32'd0; 
32'd2230: dataIn2 = 32'd0; 
32'd2231: dataIn2 = 32'd0; 
32'd2232: dataIn2 = 32'd0; 
32'd2233: dataIn2 = 32'd0; 
32'd2234: dataIn2 = 32'd1; 
32'd2235: dataIn2 = 32'd0; 
32'd2236: dataIn2 = 32'd0; 
32'd2237: dataIn2 = 32'd0; 
32'd2238: dataIn2 = 32'd0; 
32'd2239: dataIn2 = 32'd1; 
32'd2240: dataIn2 = 32'd1; 
32'd2241: dataIn2 = 32'd0; 
32'd2242: dataIn2 = 32'd1; 
32'd2243: dataIn2 = 32'd0; 
32'd2244: dataIn2 = 32'd1; 
32'd2245: dataIn2 = 32'd0; 
32'd2246: dataIn2 = 32'd0; 
32'd2247: dataIn2 = 32'd1; 
32'd2248: dataIn2 = 32'd1; 
32'd2249: dataIn2 = 32'd1; 
32'd2250: dataIn2 = 32'd0; 
32'd2251: dataIn2 = 32'd0; 
32'd2252: dataIn2 = 32'd0; 
32'd2253: dataIn2 = 32'd0; 
32'd2254: dataIn2 = 32'd1; 
32'd2255: dataIn2 = 32'd0; 
32'd2256: dataIn2 = 32'd1; 
32'd2257: dataIn2 = 32'd1; 
32'd2258: dataIn2 = 32'd0; 
32'd2259: dataIn2 = 32'd0; 
32'd2260: dataIn2 = 32'd0; 
32'd2261: dataIn2 = 32'd1; 
32'd2262: dataIn2 = 32'd1; 
32'd2263: dataIn2 = 32'd1; 
32'd2264: dataIn2 = 32'd0; 
32'd2265: dataIn2 = 32'd1; 
32'd2266: dataIn2 = 32'd1; 
32'd2267: dataIn2 = 32'd1; 
32'd2268: dataIn2 = 32'd0; 
32'd2269: dataIn2 = 32'd1; 
32'd2270: dataIn2 = 32'd0; 
32'd2271: dataIn2 = 32'd1; 
32'd2272: dataIn2 = 32'd1; 
32'd2273: dataIn2 = 32'd1; 
32'd2274: dataIn2 = 32'd0; 
32'd2275: dataIn2 = 32'd0; 
32'd2276: dataIn2 = 32'd1; 
32'd2277: dataIn2 = 32'd1; 
32'd2278: dataIn2 = 32'd1; 
32'd2279: dataIn2 = 32'd0; 
32'd2280: dataIn2 = 32'd1; 
32'd2281: dataIn2 = 32'd1; 
32'd2282: dataIn2 = 32'd1; 
32'd2283: dataIn2 = 32'd1; 
32'd2284: dataIn2 = 32'd0; 
32'd2285: dataIn2 = 32'd0; 
32'd2286: dataIn2 = 32'd0; 
32'd2287: dataIn2 = 32'd0; 
32'd2288: dataIn2 = 32'd1; 
32'd2289: dataIn2 = 32'd0; 
32'd2290: dataIn2 = 32'd1; 
32'd2291: dataIn2 = 32'd1; 
32'd2292: dataIn2 = 32'd0; 
32'd2293: dataIn2 = 32'd0; 
32'd2294: dataIn2 = 32'd1; 
32'd2295: dataIn2 = 32'd0; 
32'd2296: dataIn2 = 32'd1; 
32'd2297: dataIn2 = 32'd1; 
32'd2298: dataIn2 = 32'd1; 
32'd2299: dataIn2 = 32'd0; 
32'd2300: dataIn2 = 32'd1; 
32'd2301: dataIn2 = 32'd1; 
32'd2302: dataIn2 = 32'd1; 
32'd2303: dataIn2 = 32'd1; 
32'd2304: dataIn2 = 32'd1; 
32'd2305: dataIn2 = 32'd1; 
32'd2306: dataIn2 = 32'd1; 
32'd2307: dataIn2 = 32'd0; 
32'd2308: dataIn2 = 32'd1; 
32'd2309: dataIn2 = 32'd1; 
32'd2310: dataIn2 = 32'd1; 
32'd2311: dataIn2 = 32'd0; 
32'd2312: dataIn2 = 32'd0; 
32'd2313: dataIn2 = 32'd0; 
32'd2314: dataIn2 = 32'd0; 
32'd2315: dataIn2 = 32'd1; 
32'd2316: dataIn2 = 32'd1; 
32'd2317: dataIn2 = 32'd0; 
32'd2318: dataIn2 = 32'd1; 
32'd2319: dataIn2 = 32'd1; 
32'd2320: dataIn2 = 32'd1; 
32'd2321: dataIn2 = 32'd0; 
32'd2322: dataIn2 = 32'd0; 
32'd2323: dataIn2 = 32'd1; 
32'd2324: dataIn2 = 32'd1; 
32'd2325: dataIn2 = 32'd0; 
32'd2326: dataIn2 = 32'd1; 
32'd2327: dataIn2 = 32'd0; 
32'd2328: dataIn2 = 32'd0; 
32'd2329: dataIn2 = 32'd0; 
32'd2330: dataIn2 = 32'd0; 
32'd2331: dataIn2 = 32'd0; 
32'd2332: dataIn2 = 32'd1; 
32'd2333: dataIn2 = 32'd1; 
32'd2334: dataIn2 = 32'd0; 
32'd2335: dataIn2 = 32'd0; 
32'd2336: dataIn2 = 32'd1; 
32'd2337: dataIn2 = 32'd0; 
32'd2338: dataIn2 = 32'd0; 
32'd2339: dataIn2 = 32'd0; 
32'd2340: dataIn2 = 32'd0; 
32'd2341: dataIn2 = 32'd0; 
32'd2342: dataIn2 = 32'd0; 
32'd2343: dataIn2 = 32'd1; 
32'd2344: dataIn2 = 32'd1; 
32'd2345: dataIn2 = 32'd1; 
32'd2346: dataIn2 = 32'd1; 
32'd2347: dataIn2 = 32'd1; 
32'd2348: dataIn2 = 32'd0; 
32'd2349: dataIn2 = 32'd1; 
32'd2350: dataIn2 = 32'd1; 
32'd2351: dataIn2 = 32'd1; 
32'd2352: dataIn2 = 32'd0; 
32'd2353: dataIn2 = 32'd0; 
32'd2354: dataIn2 = 32'd1; 
32'd2355: dataIn2 = 32'd1; 
32'd2356: dataIn2 = 32'd1; 
32'd2357: dataIn2 = 32'd0; 
32'd2358: dataIn2 = 32'd0; 
32'd2359: dataIn2 = 32'd0; 
32'd2360: dataIn2 = 32'd1; 
32'd2361: dataIn2 = 32'd0; 
32'd2362: dataIn2 = 32'd0; 
32'd2363: dataIn2 = 32'd0; 
32'd2364: dataIn2 = 32'd0; 
32'd2365: dataIn2 = 32'd0; 
32'd2366: dataIn2 = 32'd0; 
32'd2367: dataIn2 = 32'd1; 
32'd2368: dataIn2 = 32'd0; 
32'd2369: dataIn2 = 32'd0; 
32'd2370: dataIn2 = 32'd0; 
32'd2371: dataIn2 = 32'd1; 
32'd2372: dataIn2 = 32'd0; 
32'd2373: dataIn2 = 32'd0; 
32'd2374: dataIn2 = 32'd0; 
32'd2375: dataIn2 = 32'd1; 
32'd2376: dataIn2 = 32'd1; 
32'd2377: dataIn2 = 32'd0; 
32'd2378: dataIn2 = 32'd0; 
32'd2379: dataIn2 = 32'd0; 
32'd2380: dataIn2 = 32'd0; 
32'd2381: dataIn2 = 32'd0; 
32'd2382: dataIn2 = 32'd1; 
32'd2383: dataIn2 = 32'd1; 
32'd2384: dataIn2 = 32'd1; 
32'd2385: dataIn2 = 32'd1; 
32'd2386: dataIn2 = 32'd0; 
32'd2387: dataIn2 = 32'd1; 
32'd2388: dataIn2 = 32'd1; 
32'd2389: dataIn2 = 32'd1; 
32'd2390: dataIn2 = 32'd0; 
32'd2391: dataIn2 = 32'd1; 
32'd2392: dataIn2 = 32'd0; 
32'd2393: dataIn2 = 32'd1; 
32'd2394: dataIn2 = 32'd0; 
32'd2395: dataIn2 = 32'd1; 
32'd2396: dataIn2 = 32'd0; 
32'd2397: dataIn2 = 32'd1; 
32'd2398: dataIn2 = 32'd0; 
32'd2399: dataIn2 = 32'd1; 
32'd2400: dataIn2 = 32'd1; 
32'd2401: dataIn2 = 32'd0; 
32'd2402: dataIn2 = 32'd1; 
32'd2403: dataIn2 = 32'd0; 
32'd2404: dataIn2 = 32'd0; 
32'd2405: dataIn2 = 32'd1; 
32'd2406: dataIn2 = 32'd0; 
32'd2407: dataIn2 = 32'd0; 
32'd2408: dataIn2 = 32'd1; 
32'd2409: dataIn2 = 32'd0; 
32'd2410: dataIn2 = 32'd0; 
32'd2411: dataIn2 = 32'd1; 
32'd2412: dataIn2 = 32'd0; 
32'd2413: dataIn2 = 32'd1; 
32'd2414: dataIn2 = 32'd1; 
32'd2415: dataIn2 = 32'd0; 
32'd2416: dataIn2 = 32'd1; 
32'd2417: dataIn2 = 32'd1; 
32'd2418: dataIn2 = 32'd1; 
32'd2419: dataIn2 = 32'd1; 
32'd2420: dataIn2 = 32'd0; 
32'd2421: dataIn2 = 32'd1; 
32'd2422: dataIn2 = 32'd0; 
32'd2423: dataIn2 = 32'd0; 
32'd2424: dataIn2 = 32'd1; 
32'd2425: dataIn2 = 32'd0; 
32'd2426: dataIn2 = 32'd0; 
32'd2427: dataIn2 = 32'd0; 
32'd2428: dataIn2 = 32'd1; 
32'd2429: dataIn2 = 32'd0; 
32'd2430: dataIn2 = 32'd0; 
32'd2431: dataIn2 = 32'd0; 
32'd2432: dataIn2 = 32'd1; 
32'd2433: dataIn2 = 32'd0; 
32'd2434: dataIn2 = 32'd1; 
32'd2435: dataIn2 = 32'd1; 
32'd2436: dataIn2 = 32'd1; 
32'd2437: dataIn2 = 32'd1; 
32'd2438: dataIn2 = 32'd1; 
32'd2439: dataIn2 = 32'd0; 
32'd2440: dataIn2 = 32'd0; 
32'd2441: dataIn2 = 32'd1; 
32'd2442: dataIn2 = 32'd0; 
32'd2443: dataIn2 = 32'd1; 
32'd2444: dataIn2 = 32'd1; 
32'd2445: dataIn2 = 32'd1; 
32'd2446: dataIn2 = 32'd1; 
32'd2447: dataIn2 = 32'd0; 
32'd2448: dataIn2 = 32'd1; 
32'd2449: dataIn2 = 32'd1; 
32'd2450: dataIn2 = 32'd0; 
32'd2451: dataIn2 = 32'd1; 
32'd2452: dataIn2 = 32'd1; 
32'd2453: dataIn2 = 32'd0; 
32'd2454: dataIn2 = 32'd0; 
32'd2455: dataIn2 = 32'd0; 
32'd2456: dataIn2 = 32'd0; 
32'd2457: dataIn2 = 32'd1; 
32'd2458: dataIn2 = 32'd0; 
32'd2459: dataIn2 = 32'd0; 
32'd2460: dataIn2 = 32'd1; 
32'd2461: dataIn2 = 32'd0; 
32'd2462: dataIn2 = 32'd1; 
32'd2463: dataIn2 = 32'd0; 
32'd2464: dataIn2 = 32'd0; 
32'd2465: dataIn2 = 32'd0; 
32'd2466: dataIn2 = 32'd1; 
32'd2467: dataIn2 = 32'd0; 
32'd2468: dataIn2 = 32'd0; 
32'd2469: dataIn2 = 32'd0; 
32'd2470: dataIn2 = 32'd0; 
32'd2471: dataIn2 = 32'd0; 
32'd2472: dataIn2 = 32'd1; 
32'd2473: dataIn2 = 32'd1; 
32'd2474: dataIn2 = 32'd0; 
32'd2475: dataIn2 = 32'd1; 
32'd2476: dataIn2 = 32'd1; 
32'd2477: dataIn2 = 32'd1; 
32'd2478: dataIn2 = 32'd0; 
32'd2479: dataIn2 = 32'd1; 
32'd2480: dataIn2 = 32'd0; 
32'd2481: dataIn2 = 32'd0; 
32'd2482: dataIn2 = 32'd0; 
32'd2483: dataIn2 = 32'd1; 
32'd2484: dataIn2 = 32'd0; 
32'd2485: dataIn2 = 32'd1; 
32'd2486: dataIn2 = 32'd0; 
32'd2487: dataIn2 = 32'd0; 
32'd2488: dataIn2 = 32'd1; 
32'd2489: dataIn2 = 32'd1; 
32'd2490: dataIn2 = 32'd1; 
32'd2491: dataIn2 = 32'd1; 
32'd2492: dataIn2 = 32'd1; 
32'd2493: dataIn2 = 32'd0; 
32'd2494: dataIn2 = 32'd0; 
32'd2495: dataIn2 = 32'd0; 
32'd2496: dataIn2 = 32'd1; 
32'd2497: dataIn2 = 32'd0; 
32'd2498: dataIn2 = 32'd1; 
32'd2499: dataIn2 = 32'd1; 
32'd2500: dataIn2 = 32'd0; 
32'd2501: dataIn2 = 32'd1; 
32'd2502: dataIn2 = 32'd1; 
32'd2503: dataIn2 = 32'd1; 
32'd2504: dataIn2 = 32'd1; 
32'd2505: dataIn2 = 32'd0; 
32'd2506: dataIn2 = 32'd0; 
32'd2507: dataIn2 = 32'd1; 
32'd2508: dataIn2 = 32'd1; 
32'd2509: dataIn2 = 32'd1; 
32'd2510: dataIn2 = 32'd1; 
32'd2511: dataIn2 = 32'd1; 
32'd2512: dataIn2 = 32'd1; 
32'd2513: dataIn2 = 32'd1; 
32'd2514: dataIn2 = 32'd1; 
32'd2515: dataIn2 = 32'd0; 
32'd2516: dataIn2 = 32'd0; 
32'd2517: dataIn2 = 32'd0; 
32'd2518: dataIn2 = 32'd0; 
32'd2519: dataIn2 = 32'd0; 
32'd2520: dataIn2 = 32'd1; 
32'd2521: dataIn2 = 32'd0; 
32'd2522: dataIn2 = 32'd1; 
32'd2523: dataIn2 = 32'd0; 
32'd2524: dataIn2 = 32'd0; 
32'd2525: dataIn2 = 32'd1; 
32'd2526: dataIn2 = 32'd1; 
32'd2527: dataIn2 = 32'd0; 
32'd2528: dataIn2 = 32'd0; 
32'd2529: dataIn2 = 32'd0; 
32'd2530: dataIn2 = 32'd1; 
32'd2531: dataIn2 = 32'd0; 
32'd2532: dataIn2 = 32'd0; 
32'd2533: dataIn2 = 32'd1; 
32'd2534: dataIn2 = 32'd0; 
32'd2535: dataIn2 = 32'd0; 
32'd2536: dataIn2 = 32'd1; 
32'd2537: dataIn2 = 32'd0; 
32'd2538: dataIn2 = 32'd1; 
32'd2539: dataIn2 = 32'd0; 
32'd2540: dataIn2 = 32'd0; 
32'd2541: dataIn2 = 32'd1; 
32'd2542: dataIn2 = 32'd1; 
32'd2543: dataIn2 = 32'd0; 
32'd2544: dataIn2 = 32'd1; 
32'd2545: dataIn2 = 32'd1; 
32'd2546: dataIn2 = 32'd0; 
32'd2547: dataIn2 = 32'd0; 
32'd2548: dataIn2 = 32'd0; 
32'd2549: dataIn2 = 32'd0; 
32'd2550: dataIn2 = 32'd0; 
32'd2551: dataIn2 = 32'd0; 
32'd2552: dataIn2 = 32'd0; 
32'd2553: dataIn2 = 32'd0; 
32'd2554: dataIn2 = 32'd1; 
32'd2555: dataIn2 = 32'd0; 
32'd2556: dataIn2 = 32'd0; 
32'd2557: dataIn2 = 32'd0; 
32'd2558: dataIn2 = 32'd0; 
32'd2559: dataIn2 = 32'd1; 
32'd2560: dataIn2 = 32'd0; 
32'd2561: dataIn2 = 32'd1; 
32'd2562: dataIn2 = 32'd1; 
32'd2563: dataIn2 = 32'd0; 
32'd2564: dataIn2 = 32'd0; 
32'd2565: dataIn2 = 32'd0; 
32'd2566: dataIn2 = 32'd1; 
32'd2567: dataIn2 = 32'd1; 
32'd2568: dataIn2 = 32'd0; 
32'd2569: dataIn2 = 32'd1; 
32'd2570: dataIn2 = 32'd1; 
32'd2571: dataIn2 = 32'd0; 
32'd2572: dataIn2 = 32'd0; 
32'd2573: dataIn2 = 32'd1; 
32'd2574: dataIn2 = 32'd0; 
32'd2575: dataIn2 = 32'd1; 
32'd2576: dataIn2 = 32'd1; 
32'd2577: dataIn2 = 32'd1; 
32'd2578: dataIn2 = 32'd1; 
32'd2579: dataIn2 = 32'd1; 
32'd2580: dataIn2 = 32'd0; 
32'd2581: dataIn2 = 32'd0; 
32'd2582: dataIn2 = 32'd0; 
32'd2583: dataIn2 = 32'd1; 
32'd2584: dataIn2 = 32'd1; 
32'd2585: dataIn2 = 32'd0; 
32'd2586: dataIn2 = 32'd0; 
32'd2587: dataIn2 = 32'd0; 
32'd2588: dataIn2 = 32'd1; 
32'd2589: dataIn2 = 32'd0; 
32'd2590: dataIn2 = 32'd0; 
32'd2591: dataIn2 = 32'd0; 
32'd2592: dataIn2 = 32'd1; 
32'd2593: dataIn2 = 32'd0; 
32'd2594: dataIn2 = 32'd0; 
32'd2595: dataIn2 = 32'd1; 
32'd2596: dataIn2 = 32'd0; 
32'd2597: dataIn2 = 32'd0; 
32'd2598: dataIn2 = 32'd0; 
32'd2599: dataIn2 = 32'd0; 
32'd2600: dataIn2 = 32'd0; 
32'd2601: dataIn2 = 32'd0; 
32'd2602: dataIn2 = 32'd1; 
32'd2603: dataIn2 = 32'd0; 
32'd2604: dataIn2 = 32'd1; 
32'd2605: dataIn2 = 32'd0; 
32'd2606: dataIn2 = 32'd0; 
32'd2607: dataIn2 = 32'd1; 
32'd2608: dataIn2 = 32'd1; 
32'd2609: dataIn2 = 32'd1; 
32'd2610: dataIn2 = 32'd1; 
32'd2611: dataIn2 = 32'd1; 
32'd2612: dataIn2 = 32'd0; 
32'd2613: dataIn2 = 32'd0; 
32'd2614: dataIn2 = 32'd0; 
32'd2615: dataIn2 = 32'd0; 
32'd2616: dataIn2 = 32'd0; 
32'd2617: dataIn2 = 32'd0; 
32'd2618: dataIn2 = 32'd0; 
32'd2619: dataIn2 = 32'd0; 
32'd2620: dataIn2 = 32'd0; 
32'd2621: dataIn2 = 32'd0; 
32'd2622: dataIn2 = 32'd0; 
32'd2623: dataIn2 = 32'd1; 
32'd2624: dataIn2 = 32'd0; 
32'd2625: dataIn2 = 32'd0; 
32'd2626: dataIn2 = 32'd0; 
32'd2627: dataIn2 = 32'd0; 
32'd2628: dataIn2 = 32'd0; 
32'd2629: dataIn2 = 32'd1; 
32'd2630: dataIn2 = 32'd1; 
32'd2631: dataIn2 = 32'd1; 
32'd2632: dataIn2 = 32'd0; 
32'd2633: dataIn2 = 32'd1; 
32'd2634: dataIn2 = 32'd0; 
32'd2635: dataIn2 = 32'd1; 
32'd2636: dataIn2 = 32'd0; 
32'd2637: dataIn2 = 32'd0; 
32'd2638: dataIn2 = 32'd0; 
32'd2639: dataIn2 = 32'd0; 
32'd2640: dataIn2 = 32'd1; 
32'd2641: dataIn2 = 32'd1; 
32'd2642: dataIn2 = 32'd0; 
32'd2643: dataIn2 = 32'd0; 
32'd2644: dataIn2 = 32'd0; 
32'd2645: dataIn2 = 32'd1; 
32'd2646: dataIn2 = 32'd0; 
32'd2647: dataIn2 = 32'd1; 
32'd2648: dataIn2 = 32'd1; 
32'd2649: dataIn2 = 32'd1; 
32'd2650: dataIn2 = 32'd0; 
32'd2651: dataIn2 = 32'd1; 
32'd2652: dataIn2 = 32'd1; 
32'd2653: dataIn2 = 32'd1; 
32'd2654: dataIn2 = 32'd1; 
32'd2655: dataIn2 = 32'd0; 
32'd2656: dataIn2 = 32'd1; 
32'd2657: dataIn2 = 32'd1; 
32'd2658: dataIn2 = 32'd1; 
32'd2659: dataIn2 = 32'd1; 
32'd2660: dataIn2 = 32'd1; 
32'd2661: dataIn2 = 32'd0; 
32'd2662: dataIn2 = 32'd0; 
32'd2663: dataIn2 = 32'd0; 
32'd2664: dataIn2 = 32'd1; 
32'd2665: dataIn2 = 32'd1; 
32'd2666: dataIn2 = 32'd0; 
32'd2667: dataIn2 = 32'd0; 
32'd2668: dataIn2 = 32'd1; 
32'd2669: dataIn2 = 32'd1; 
32'd2670: dataIn2 = 32'd0; 
32'd2671: dataIn2 = 32'd1; 
32'd2672: dataIn2 = 32'd1; 
32'd2673: dataIn2 = 32'd0; 
32'd2674: dataIn2 = 32'd1; 
32'd2675: dataIn2 = 32'd1; 
32'd2676: dataIn2 = 32'd0; 
32'd2677: dataIn2 = 32'd0; 
32'd2678: dataIn2 = 32'd1; 
32'd2679: dataIn2 = 32'd0; 
32'd2680: dataIn2 = 32'd1; 
32'd2681: dataIn2 = 32'd0; 
32'd2682: dataIn2 = 32'd0; 
32'd2683: dataIn2 = 32'd0; 
32'd2684: dataIn2 = 32'd0; 
32'd2685: dataIn2 = 32'd1; 
32'd2686: dataIn2 = 32'd1; 
32'd2687: dataIn2 = 32'd1; 
32'd2688: dataIn2 = 32'd1; 
32'd2689: dataIn2 = 32'd0; 
32'd2690: dataIn2 = 32'd0; 
32'd2691: dataIn2 = 32'd0; 
32'd2692: dataIn2 = 32'd1; 
32'd2693: dataIn2 = 32'd1; 
32'd2694: dataIn2 = 32'd1; 
32'd2695: dataIn2 = 32'd0; 
32'd2696: dataIn2 = 32'd0; 
32'd2697: dataIn2 = 32'd0; 
32'd2698: dataIn2 = 32'd1; 
32'd2699: dataIn2 = 32'd1; 
32'd2700: dataIn2 = 32'd0; 
32'd2701: dataIn2 = 32'd0; 
32'd2702: dataIn2 = 32'd0; 
32'd2703: dataIn2 = 32'd1; 
32'd2704: dataIn2 = 32'd1; 
32'd2705: dataIn2 = 32'd1; 
32'd2706: dataIn2 = 32'd1; 
32'd2707: dataIn2 = 32'd0; 
32'd2708: dataIn2 = 32'd0; 
32'd2709: dataIn2 = 32'd0; 
32'd2710: dataIn2 = 32'd1; 
32'd2711: dataIn2 = 32'd1; 
32'd2712: dataIn2 = 32'd1; 
32'd2713: dataIn2 = 32'd1; 
32'd2714: dataIn2 = 32'd0; 
32'd2715: dataIn2 = 32'd0; 
32'd2716: dataIn2 = 32'd1; 
32'd2717: dataIn2 = 32'd1; 
32'd2718: dataIn2 = 32'd1; 
32'd2719: dataIn2 = 32'd1; 
32'd2720: dataIn2 = 32'd1; 
32'd2721: dataIn2 = 32'd1; 
32'd2722: dataIn2 = 32'd0; 
32'd2723: dataIn2 = 32'd0; 
32'd2724: dataIn2 = 32'd1; 
32'd2725: dataIn2 = 32'd1; 
32'd2726: dataIn2 = 32'd0; 
32'd2727: dataIn2 = 32'd0; 
32'd2728: dataIn2 = 32'd0; 
32'd2729: dataIn2 = 32'd0; 
32'd2730: dataIn2 = 32'd1; 
32'd2731: dataIn2 = 32'd0; 
32'd2732: dataIn2 = 32'd0; 
32'd2733: dataIn2 = 32'd1; 
32'd2734: dataIn2 = 32'd1; 
32'd2735: dataIn2 = 32'd0; 
32'd2736: dataIn2 = 32'd0; 
32'd2737: dataIn2 = 32'd0; 
32'd2738: dataIn2 = 32'd1; 
32'd2739: dataIn2 = 32'd1; 
32'd2740: dataIn2 = 32'd1; 
32'd2741: dataIn2 = 32'd1; 
32'd2742: dataIn2 = 32'd0; 
32'd2743: dataIn2 = 32'd1; 
32'd2744: dataIn2 = 32'd0; 
32'd2745: dataIn2 = 32'd0; 
32'd2746: dataIn2 = 32'd1; 
32'd2747: dataIn2 = 32'd0; 
32'd2748: dataIn2 = 32'd0; 
32'd2749: dataIn2 = 32'd0; 
32'd2750: dataIn2 = 32'd0; 
32'd2751: dataIn2 = 32'd1; 
32'd2752: dataIn2 = 32'd1; 
32'd2753: dataIn2 = 32'd1; 
32'd2754: dataIn2 = 32'd1; 
32'd2755: dataIn2 = 32'd0; 
32'd2756: dataIn2 = 32'd0; 
32'd2757: dataIn2 = 32'd1; 
32'd2758: dataIn2 = 32'd1; 
32'd2759: dataIn2 = 32'd0; 
32'd2760: dataIn2 = 32'd0; 
32'd2761: dataIn2 = 32'd0; 
32'd2762: dataIn2 = 32'd1; 
32'd2763: dataIn2 = 32'd0; 
32'd2764: dataIn2 = 32'd1; 
32'd2765: dataIn2 = 32'd0; 
32'd2766: dataIn2 = 32'd0; 
32'd2767: dataIn2 = 32'd1; 
32'd2768: dataIn2 = 32'd0; 
32'd2769: dataIn2 = 32'd0; 
32'd2770: dataIn2 = 32'd1; 
32'd2771: dataIn2 = 32'd0; 
32'd2772: dataIn2 = 32'd0; 
32'd2773: dataIn2 = 32'd1; 
32'd2774: dataIn2 = 32'd1; 
32'd2775: dataIn2 = 32'd1; 
32'd2776: dataIn2 = 32'd1; 
32'd2777: dataIn2 = 32'd0; 
32'd2778: dataIn2 = 32'd0; 
32'd2779: dataIn2 = 32'd0; 
32'd2780: dataIn2 = 32'd1; 
32'd2781: dataIn2 = 32'd1; 
32'd2782: dataIn2 = 32'd1; 
32'd2783: dataIn2 = 32'd0; 
32'd2784: dataIn2 = 32'd0; 
32'd2785: dataIn2 = 32'd1; 
32'd2786: dataIn2 = 32'd1; 
32'd2787: dataIn2 = 32'd0; 
32'd2788: dataIn2 = 32'd0; 
32'd2789: dataIn2 = 32'd1; 
32'd2790: dataIn2 = 32'd1; 
32'd2791: dataIn2 = 32'd1; 
32'd2792: dataIn2 = 32'd1; 
32'd2793: dataIn2 = 32'd0; 
32'd2794: dataIn2 = 32'd1; 
32'd2795: dataIn2 = 32'd1; 
32'd2796: dataIn2 = 32'd1; 
32'd2797: dataIn2 = 32'd0; 
32'd2798: dataIn2 = 32'd0; 
32'd2799: dataIn2 = 32'd0; 
32'd2800: dataIn2 = 32'd1; 
32'd2801: dataIn2 = 32'd0; 
32'd2802: dataIn2 = 32'd0; 
32'd2803: dataIn2 = 32'd1; 
32'd2804: dataIn2 = 32'd0; 
32'd2805: dataIn2 = 32'd0; 
32'd2806: dataIn2 = 32'd0; 
32'd2807: dataIn2 = 32'd1; 
32'd2808: dataIn2 = 32'd0; 
32'd2809: dataIn2 = 32'd0; 
32'd2810: dataIn2 = 32'd0; 
32'd2811: dataIn2 = 32'd1; 
32'd2812: dataIn2 = 32'd0; 
32'd2813: dataIn2 = 32'd0; 
32'd2814: dataIn2 = 32'd1; 
32'd2815: dataIn2 = 32'd1; 
32'd2816: dataIn2 = 32'd1; 
32'd2817: dataIn2 = 32'd1; 
32'd2818: dataIn2 = 32'd1; 
32'd2819: dataIn2 = 32'd0; 
32'd2820: dataIn2 = 32'd0; 
32'd2821: dataIn2 = 32'd0; 
32'd2822: dataIn2 = 32'd1; 
32'd2823: dataIn2 = 32'd1; 
32'd2824: dataIn2 = 32'd1; 
32'd2825: dataIn2 = 32'd1; 
32'd2826: dataIn2 = 32'd1; 
32'd2827: dataIn2 = 32'd0; 
32'd2828: dataIn2 = 32'd0; 
32'd2829: dataIn2 = 32'd1; 
32'd2830: dataIn2 = 32'd0; 
32'd2831: dataIn2 = 32'd1; 
32'd2832: dataIn2 = 32'd0; 
32'd2833: dataIn2 = 32'd1; 
32'd2834: dataIn2 = 32'd0; 
32'd2835: dataIn2 = 32'd1; 
32'd2836: dataIn2 = 32'd1; 
32'd2837: dataIn2 = 32'd0; 
32'd2838: dataIn2 = 32'd0; 
32'd2839: dataIn2 = 32'd0; 
32'd2840: dataIn2 = 32'd0; 
32'd2841: dataIn2 = 32'd0; 
32'd2842: dataIn2 = 32'd0; 
32'd2843: dataIn2 = 32'd0; 
32'd2844: dataIn2 = 32'd0; 
32'd2845: dataIn2 = 32'd1; 
32'd2846: dataIn2 = 32'd0; 
32'd2847: dataIn2 = 32'd0; 
32'd2848: dataIn2 = 32'd1; 
32'd2849: dataIn2 = 32'd0; 
32'd2850: dataIn2 = 32'd1; 
32'd2851: dataIn2 = 32'd1; 
32'd2852: dataIn2 = 32'd0; 
32'd2853: dataIn2 = 32'd1; 
32'd2854: dataIn2 = 32'd0; 
32'd2855: dataIn2 = 32'd1; 
32'd2856: dataIn2 = 32'd0; 
32'd2857: dataIn2 = 32'd1; 
32'd2858: dataIn2 = 32'd0; 
32'd2859: dataIn2 = 32'd0; 
32'd2860: dataIn2 = 32'd1; 
32'd2861: dataIn2 = 32'd1; 
32'd2862: dataIn2 = 32'd1; 
32'd2863: dataIn2 = 32'd0; 
32'd2864: dataIn2 = 32'd0; 
32'd2865: dataIn2 = 32'd1; 
32'd2866: dataIn2 = 32'd1; 
32'd2867: dataIn2 = 32'd1; 
32'd2868: dataIn2 = 32'd1; 
32'd2869: dataIn2 = 32'd1; 
32'd2870: dataIn2 = 32'd0; 
32'd2871: dataIn2 = 32'd0; 
32'd2872: dataIn2 = 32'd0; 
32'd2873: dataIn2 = 32'd0; 
32'd2874: dataIn2 = 32'd1; 
32'd2875: dataIn2 = 32'd0; 
32'd2876: dataIn2 = 32'd0; 
32'd2877: dataIn2 = 32'd1; 
32'd2878: dataIn2 = 32'd1; 
32'd2879: dataIn2 = 32'd0; 
32'd2880: dataIn2 = 32'd0; 
32'd2881: dataIn2 = 32'd0; 
32'd2882: dataIn2 = 32'd0; 
32'd2883: dataIn2 = 32'd0; 
32'd2884: dataIn2 = 32'd0; 
32'd2885: dataIn2 = 32'd1; 
32'd2886: dataIn2 = 32'd1; 
32'd2887: dataIn2 = 32'd0; 
32'd2888: dataIn2 = 32'd0; 
32'd2889: dataIn2 = 32'd0; 
32'd2890: dataIn2 = 32'd0; 
32'd2891: dataIn2 = 32'd0; 
32'd2892: dataIn2 = 32'd1; 
32'd2893: dataIn2 = 32'd0; 
32'd2894: dataIn2 = 32'd0; 
32'd2895: dataIn2 = 32'd1; 
32'd2896: dataIn2 = 32'd1; 
32'd2897: dataIn2 = 32'd1; 
32'd2898: dataIn2 = 32'd1; 
32'd2899: dataIn2 = 32'd1; 
32'd2900: dataIn2 = 32'd1; 
32'd2901: dataIn2 = 32'd0; 
32'd2902: dataIn2 = 32'd0; 
32'd2903: dataIn2 = 32'd1; 
32'd2904: dataIn2 = 32'd1; 
32'd2905: dataIn2 = 32'd0; 
32'd2906: dataIn2 = 32'd0; 
32'd2907: dataIn2 = 32'd1; 
32'd2908: dataIn2 = 32'd1; 
32'd2909: dataIn2 = 32'd1; 
32'd2910: dataIn2 = 32'd0; 
32'd2911: dataIn2 = 32'd0; 
32'd2912: dataIn2 = 32'd0; 
32'd2913: dataIn2 = 32'd0; 
32'd2914: dataIn2 = 32'd1; 
32'd2915: dataIn2 = 32'd0; 
32'd2916: dataIn2 = 32'd0; 
32'd2917: dataIn2 = 32'd0; 
32'd2918: dataIn2 = 32'd0; 
32'd2919: dataIn2 = 32'd1; 
32'd2920: dataIn2 = 32'd0; 
32'd2921: dataIn2 = 32'd1; 
32'd2922: dataIn2 = 32'd0; 
32'd2923: dataIn2 = 32'd0; 
32'd2924: dataIn2 = 32'd1; 
32'd2925: dataIn2 = 32'd1; 
32'd2926: dataIn2 = 32'd1; 
32'd2927: dataIn2 = 32'd1; 
32'd2928: dataIn2 = 32'd0; 
32'd2929: dataIn2 = 32'd0; 
32'd2930: dataIn2 = 32'd1; 
32'd2931: dataIn2 = 32'd0; 
32'd2932: dataIn2 = 32'd0; 
32'd2933: dataIn2 = 32'd1; 
32'd2934: dataIn2 = 32'd1; 
32'd2935: dataIn2 = 32'd1; 
32'd2936: dataIn2 = 32'd1; 
32'd2937: dataIn2 = 32'd1; 
32'd2938: dataIn2 = 32'd0; 
32'd2939: dataIn2 = 32'd0; 
32'd2940: dataIn2 = 32'd0; 
32'd2941: dataIn2 = 32'd0; 
32'd2942: dataIn2 = 32'd1; 
32'd2943: dataIn2 = 32'd1; 
32'd2944: dataIn2 = 32'd1; 
32'd2945: dataIn2 = 32'd1; 
32'd2946: dataIn2 = 32'd1; 
32'd2947: dataIn2 = 32'd0; 
32'd2948: dataIn2 = 32'd1; 
32'd2949: dataIn2 = 32'd1; 
32'd2950: dataIn2 = 32'd1; 
32'd2951: dataIn2 = 32'd0; 
32'd2952: dataIn2 = 32'd1; 
32'd2953: dataIn2 = 32'd0; 
32'd2954: dataIn2 = 32'd1; 
32'd2955: dataIn2 = 32'd1; 
32'd2956: dataIn2 = 32'd0; 
32'd2957: dataIn2 = 32'd0; 
32'd2958: dataIn2 = 32'd0; 
32'd2959: dataIn2 = 32'd1; 
32'd2960: dataIn2 = 32'd0; 
32'd2961: dataIn2 = 32'd1; 
32'd2962: dataIn2 = 32'd1; 
32'd2963: dataIn2 = 32'd0; 
32'd2964: dataIn2 = 32'd0; 
32'd2965: dataIn2 = 32'd1; 
32'd2966: dataIn2 = 32'd0; 
32'd2967: dataIn2 = 32'd0; 
32'd2968: dataIn2 = 32'd1; 
32'd2969: dataIn2 = 32'd0; 
32'd2970: dataIn2 = 32'd1; 
32'd2971: dataIn2 = 32'd1; 
32'd2972: dataIn2 = 32'd1; 
32'd2973: dataIn2 = 32'd0; 
32'd2974: dataIn2 = 32'd0; 
32'd2975: dataIn2 = 32'd0; 
32'd2976: dataIn2 = 32'd1; 
32'd2977: dataIn2 = 32'd0; 
32'd2978: dataIn2 = 32'd0; 
32'd2979: dataIn2 = 32'd0; 
32'd2980: dataIn2 = 32'd0; 
32'd2981: dataIn2 = 32'd0; 
32'd2982: dataIn2 = 32'd1; 
32'd2983: dataIn2 = 32'd1; 
32'd2984: dataIn2 = 32'd0; 
32'd2985: dataIn2 = 32'd1; 
32'd2986: dataIn2 = 32'd0; 
32'd2987: dataIn2 = 32'd1; 
32'd2988: dataIn2 = 32'd1; 
32'd2989: dataIn2 = 32'd1; 
32'd2990: dataIn2 = 32'd1; 
32'd2991: dataIn2 = 32'd0; 
32'd2992: dataIn2 = 32'd1; 
32'd2993: dataIn2 = 32'd0; 
32'd2994: dataIn2 = 32'd0; 
32'd2995: dataIn2 = 32'd1; 
32'd2996: dataIn2 = 32'd1; 
32'd2997: dataIn2 = 32'd0; 
32'd2998: dataIn2 = 32'd1; 
32'd2999: dataIn2 = 32'd1; 
32'd3000: dataIn2 = 32'd0; 
32'd3001: dataIn2 = 32'd1; 
32'd3002: dataIn2 = 32'd0; 
32'd3003: dataIn2 = 32'd1; 
32'd3004: dataIn2 = 32'd0; 
32'd3005: dataIn2 = 32'd1; 
32'd3006: dataIn2 = 32'd1; 
32'd3007: dataIn2 = 32'd1; 
32'd3008: dataIn2 = 32'd1; 
32'd3009: dataIn2 = 32'd1; 
32'd3010: dataIn2 = 32'd0; 
32'd3011: dataIn2 = 32'd0; 
32'd3012: dataIn2 = 32'd0; 
32'd3013: dataIn2 = 32'd1; 
32'd3014: dataIn2 = 32'd0; 
32'd3015: dataIn2 = 32'd1; 
32'd3016: dataIn2 = 32'd0; 
32'd3017: dataIn2 = 32'd0; 
32'd3018: dataIn2 = 32'd0; 
32'd3019: dataIn2 = 32'd1; 
32'd3020: dataIn2 = 32'd1; 
32'd3021: dataIn2 = 32'd1; 
32'd3022: dataIn2 = 32'd0; 
32'd3023: dataIn2 = 32'd1; 
32'd3024: dataIn2 = 32'd1; 
32'd3025: dataIn2 = 32'd1; 
32'd3026: dataIn2 = 32'd1; 
32'd3027: dataIn2 = 32'd0; 
32'd3028: dataIn2 = 32'd0; 
32'd3029: dataIn2 = 32'd0; 
32'd3030: dataIn2 = 32'd0; 
32'd3031: dataIn2 = 32'd0; 
32'd3032: dataIn2 = 32'd1; 
32'd3033: dataIn2 = 32'd0; 
32'd3034: dataIn2 = 32'd1; 
32'd3035: dataIn2 = 32'd1; 
32'd3036: dataIn2 = 32'd0; 
32'd3037: dataIn2 = 32'd0; 
32'd3038: dataIn2 = 32'd1; 
32'd3039: dataIn2 = 32'd1; 
32'd3040: dataIn2 = 32'd0; 
32'd3041: dataIn2 = 32'd0; 
32'd3042: dataIn2 = 32'd1; 
32'd3043: dataIn2 = 32'd0; 
32'd3044: dataIn2 = 32'd1; 
32'd3045: dataIn2 = 32'd0; 
32'd3046: dataIn2 = 32'd0; 
32'd3047: dataIn2 = 32'd1; 
32'd3048: dataIn2 = 32'd0; 
32'd3049: dataIn2 = 32'd0; 
32'd3050: dataIn2 = 32'd0; 
32'd3051: dataIn2 = 32'd0; 
32'd3052: dataIn2 = 32'd1; 
32'd3053: dataIn2 = 32'd0; 
32'd3054: dataIn2 = 32'd0; 
32'd3055: dataIn2 = 32'd0; 
32'd3056: dataIn2 = 32'd1; 
32'd3057: dataIn2 = 32'd0; 
32'd3058: dataIn2 = 32'd1; 
32'd3059: dataIn2 = 32'd0; 
32'd3060: dataIn2 = 32'd0; 
32'd3061: dataIn2 = 32'd1; 
32'd3062: dataIn2 = 32'd0; 
32'd3063: dataIn2 = 32'd0; 
32'd3064: dataIn2 = 32'd1; 
32'd3065: dataIn2 = 32'd0; 
32'd3066: dataIn2 = 32'd0; 
32'd3067: dataIn2 = 32'd0; 
32'd3068: dataIn2 = 32'd1; 
32'd3069: dataIn2 = 32'd1; 
32'd3070: dataIn2 = 32'd0; 
32'd3071: dataIn2 = 32'd0; 
32'd3072: dataIn2 = 32'd1; 
32'd3073: dataIn2 = 32'd0; 
32'd3074: dataIn2 = 32'd1; 
32'd3075: dataIn2 = 32'd0; 
32'd3076: dataIn2 = 32'd1; 
32'd3077: dataIn2 = 32'd1; 
32'd3078: dataIn2 = 32'd1; 
32'd3079: dataIn2 = 32'd1; 
32'd3080: dataIn2 = 32'd0; 
32'd3081: dataIn2 = 32'd1; 
32'd3082: dataIn2 = 32'd1; 
32'd3083: dataIn2 = 32'd1; 
32'd3084: dataIn2 = 32'd1; 
32'd3085: dataIn2 = 32'd0; 
32'd3086: dataIn2 = 32'd0; 
32'd3087: dataIn2 = 32'd0; 
32'd3088: dataIn2 = 32'd0; 
32'd3089: dataIn2 = 32'd1; 
32'd3090: dataIn2 = 32'd0; 
32'd3091: dataIn2 = 32'd0; 
32'd3092: dataIn2 = 32'd0; 
32'd3093: dataIn2 = 32'd1; 
32'd3094: dataIn2 = 32'd0; 
32'd3095: dataIn2 = 32'd1; 
32'd3096: dataIn2 = 32'd1; 
32'd3097: dataIn2 = 32'd0; 
32'd3098: dataIn2 = 32'd1; 
32'd3099: dataIn2 = 32'd0; 
32'd3100: dataIn2 = 32'd0; 
32'd3101: dataIn2 = 32'd0; 
32'd3102: dataIn2 = 32'd1; 
32'd3103: dataIn2 = 32'd1; 
32'd3104: dataIn2 = 32'd0; 
32'd3105: dataIn2 = 32'd0; 
32'd3106: dataIn2 = 32'd0; 
32'd3107: dataIn2 = 32'd0; 
32'd3108: dataIn2 = 32'd1; 
32'd3109: dataIn2 = 32'd1; 
32'd3110: dataIn2 = 32'd1; 
32'd3111: dataIn2 = 32'd0; 
32'd3112: dataIn2 = 32'd0; 
32'd3113: dataIn2 = 32'd1; 
32'd3114: dataIn2 = 32'd0; 
32'd3115: dataIn2 = 32'd1; 
32'd3116: dataIn2 = 32'd0; 
32'd3117: dataIn2 = 32'd0; 
32'd3118: dataIn2 = 32'd1; 
32'd3119: dataIn2 = 32'd1; 
32'd3120: dataIn2 = 32'd0; 
32'd3121: dataIn2 = 32'd0; 
32'd3122: dataIn2 = 32'd0; 
32'd3123: dataIn2 = 32'd1; 
32'd3124: dataIn2 = 32'd0; 
32'd3125: dataIn2 = 32'd0; 
32'd3126: dataIn2 = 32'd0; 
32'd3127: dataIn2 = 32'd0; 
32'd3128: dataIn2 = 32'd0; 
32'd3129: dataIn2 = 32'd1; 
32'd3130: dataIn2 = 32'd0; 
32'd3131: dataIn2 = 32'd0; 
32'd3132: dataIn2 = 32'd1; 
32'd3133: dataIn2 = 32'd0; 
32'd3134: dataIn2 = 32'd1; 
32'd3135: dataIn2 = 32'd0; 
32'd3136: dataIn2 = 32'd1; 
32'd3137: dataIn2 = 32'd0; 
32'd3138: dataIn2 = 32'd1; 
32'd3139: dataIn2 = 32'd1; 
32'd3140: dataIn2 = 32'd0; 
32'd3141: dataIn2 = 32'd0; 
32'd3142: dataIn2 = 32'd0; 
32'd3143: dataIn2 = 32'd1; 
32'd3144: dataIn2 = 32'd1; 
32'd3145: dataIn2 = 32'd0; 
32'd3146: dataIn2 = 32'd0; 
32'd3147: dataIn2 = 32'd1; 
32'd3148: dataIn2 = 32'd0; 
32'd3149: dataIn2 = 32'd0; 
32'd3150: dataIn2 = 32'd1; 
32'd3151: dataIn2 = 32'd1; 
32'd3152: dataIn2 = 32'd1; 
32'd3153: dataIn2 = 32'd0; 
32'd3154: dataIn2 = 32'd1; 
32'd3155: dataIn2 = 32'd0; 
32'd3156: dataIn2 = 32'd1; 
32'd3157: dataIn2 = 32'd1; 
32'd3158: dataIn2 = 32'd0; 
32'd3159: dataIn2 = 32'd0; 
32'd3160: dataIn2 = 32'd1; 
32'd3161: dataIn2 = 32'd0; 
32'd3162: dataIn2 = 32'd1; 
32'd3163: dataIn2 = 32'd0; 
32'd3164: dataIn2 = 32'd1; 
32'd3165: dataIn2 = 32'd1; 
32'd3166: dataIn2 = 32'd0; 
32'd3167: dataIn2 = 32'd1; 
32'd3168: dataIn2 = 32'd1; 
32'd3169: dataIn2 = 32'd1; 
32'd3170: dataIn2 = 32'd1; 
32'd3171: dataIn2 = 32'd1; 
32'd3172: dataIn2 = 32'd0; 
32'd3173: dataIn2 = 32'd0; 
32'd3174: dataIn2 = 32'd1; 
32'd3175: dataIn2 = 32'd1; 
32'd3176: dataIn2 = 32'd1; 
32'd3177: dataIn2 = 32'd0; 
32'd3178: dataIn2 = 32'd0; 
32'd3179: dataIn2 = 32'd0; 
32'd3180: dataIn2 = 32'd0; 
32'd3181: dataIn2 = 32'd0; 
32'd3182: dataIn2 = 32'd0; 
32'd3183: dataIn2 = 32'd1; 
32'd3184: dataIn2 = 32'd1; 
32'd3185: dataIn2 = 32'd0; 
32'd3186: dataIn2 = 32'd1; 
32'd3187: dataIn2 = 32'd0; 
32'd3188: dataIn2 = 32'd0; 
32'd3189: dataIn2 = 32'd0; 
32'd3190: dataIn2 = 32'd0; 
32'd3191: dataIn2 = 32'd0; 
32'd3192: dataIn2 = 32'd0; 
32'd3193: dataIn2 = 32'd0; 
32'd3194: dataIn2 = 32'd0; 
32'd3195: dataIn2 = 32'd1; 
32'd3196: dataIn2 = 32'd1; 
32'd3197: dataIn2 = 32'd0; 
32'd3198: dataIn2 = 32'd0; 
32'd3199: dataIn2 = 32'd0; 
32'd3200: dataIn2 = 32'd0; 
32'd3201: dataIn2 = 32'd1; 
32'd3202: dataIn2 = 32'd1; 
32'd3203: dataIn2 = 32'd0; 
32'd3204: dataIn2 = 32'd0; 
32'd3205: dataIn2 = 32'd0; 
32'd3206: dataIn2 = 32'd1; 
32'd3207: dataIn2 = 32'd1; 
32'd3208: dataIn2 = 32'd0; 
32'd3209: dataIn2 = 32'd1; 
32'd3210: dataIn2 = 32'd1; 
32'd3211: dataIn2 = 32'd0; 
32'd3212: dataIn2 = 32'd0; 
32'd3213: dataIn2 = 32'd1; 
32'd3214: dataIn2 = 32'd0; 
32'd3215: dataIn2 = 32'd0; 
32'd3216: dataIn2 = 32'd1; 
32'd3217: dataIn2 = 32'd1; 
32'd3218: dataIn2 = 32'd0; 
32'd3219: dataIn2 = 32'd1; 
32'd3220: dataIn2 = 32'd1; 
32'd3221: dataIn2 = 32'd0; 
32'd3222: dataIn2 = 32'd1; 
32'd3223: dataIn2 = 32'd1; 
32'd3224: dataIn2 = 32'd1; 
32'd3225: dataIn2 = 32'd1; 
32'd3226: dataIn2 = 32'd0; 
32'd3227: dataIn2 = 32'd1; 
32'd3228: dataIn2 = 32'd0; 
32'd3229: dataIn2 = 32'd1; 
32'd3230: dataIn2 = 32'd0; 
32'd3231: dataIn2 = 32'd0; 
32'd3232: dataIn2 = 32'd1; 
32'd3233: dataIn2 = 32'd0; 
32'd3234: dataIn2 = 32'd1; 
32'd3235: dataIn2 = 32'd0; 
32'd3236: dataIn2 = 32'd1; 
32'd3237: dataIn2 = 32'd0; 
32'd3238: dataIn2 = 32'd0; 
32'd3239: dataIn2 = 32'd0; 
32'd3240: dataIn2 = 32'd0; 
32'd3241: dataIn2 = 32'd0; 
32'd3242: dataIn2 = 32'd1; 
32'd3243: dataIn2 = 32'd0; 
32'd3244: dataIn2 = 32'd0; 
32'd3245: dataIn2 = 32'd0; 
32'd3246: dataIn2 = 32'd1; 
32'd3247: dataIn2 = 32'd1; 
32'd3248: dataIn2 = 32'd1; 
32'd3249: dataIn2 = 32'd0; 
32'd3250: dataIn2 = 32'd1; 
32'd3251: dataIn2 = 32'd1; 
32'd3252: dataIn2 = 32'd1; 
32'd3253: dataIn2 = 32'd1; 
32'd3254: dataIn2 = 32'd0; 
32'd3255: dataIn2 = 32'd1; 
32'd3256: dataIn2 = 32'd0; 
32'd3257: dataIn2 = 32'd0; 
32'd3258: dataIn2 = 32'd1; 
32'd3259: dataIn2 = 32'd1; 
32'd3260: dataIn2 = 32'd1; 
32'd3261: dataIn2 = 32'd0; 
32'd3262: dataIn2 = 32'd0; 
32'd3263: dataIn2 = 32'd0; 
32'd3264: dataIn2 = 32'd0; 
32'd3265: dataIn2 = 32'd1; 
32'd3266: dataIn2 = 32'd0; 
32'd3267: dataIn2 = 32'd1; 
32'd3268: dataIn2 = 32'd1; 
32'd3269: dataIn2 = 32'd1; 
32'd3270: dataIn2 = 32'd0; 
32'd3271: dataIn2 = 32'd1; 
32'd3272: dataIn2 = 32'd0; 
32'd3273: dataIn2 = 32'd1; 
32'd3274: dataIn2 = 32'd1; 
32'd3275: dataIn2 = 32'd0; 
32'd3276: dataIn2 = 32'd0; 
32'd3277: dataIn2 = 32'd0; 
32'd3278: dataIn2 = 32'd1; 
32'd3279: dataIn2 = 32'd1; 
32'd3280: dataIn2 = 32'd0; 
32'd3281: dataIn2 = 32'd0; 
32'd3282: dataIn2 = 32'd0; 
32'd3283: dataIn2 = 32'd1; 
32'd3284: dataIn2 = 32'd1; 
32'd3285: dataIn2 = 32'd1; 
32'd3286: dataIn2 = 32'd0; 
32'd3287: dataIn2 = 32'd0; 
32'd3288: dataIn2 = 32'd1; 
32'd3289: dataIn2 = 32'd0; 
32'd3290: dataIn2 = 32'd1; 
32'd3291: dataIn2 = 32'd0; 
32'd3292: dataIn2 = 32'd0; 
32'd3293: dataIn2 = 32'd0; 
32'd3294: dataIn2 = 32'd0; 
32'd3295: dataIn2 = 32'd1; 
32'd3296: dataIn2 = 32'd0; 
32'd3297: dataIn2 = 32'd1; 
32'd3298: dataIn2 = 32'd1; 
32'd3299: dataIn2 = 32'd1; 
32'd3300: dataIn2 = 32'd0; 
32'd3301: dataIn2 = 32'd0; 
32'd3302: dataIn2 = 32'd1; 
32'd3303: dataIn2 = 32'd1; 
32'd3304: dataIn2 = 32'd1; 
32'd3305: dataIn2 = 32'd1; 
32'd3306: dataIn2 = 32'd1; 
32'd3307: dataIn2 = 32'd1; 
32'd3308: dataIn2 = 32'd1; 
32'd3309: dataIn2 = 32'd0; 
32'd3310: dataIn2 = 32'd1; 
32'd3311: dataIn2 = 32'd0; 
32'd3312: dataIn2 = 32'd0; 
32'd3313: dataIn2 = 32'd1; 
32'd3314: dataIn2 = 32'd0; 
32'd3315: dataIn2 = 32'd0; 
32'd3316: dataIn2 = 32'd1; 
32'd3317: dataIn2 = 32'd1; 
32'd3318: dataIn2 = 32'd1; 
32'd3319: dataIn2 = 32'd1; 
32'd3320: dataIn2 = 32'd1; 
32'd3321: dataIn2 = 32'd0; 
32'd3322: dataIn2 = 32'd0; 
32'd3323: dataIn2 = 32'd1; 
32'd3324: dataIn2 = 32'd1; 
32'd3325: dataIn2 = 32'd1; 
32'd3326: dataIn2 = 32'd0; 
32'd3327: dataIn2 = 32'd0; 
32'd3328: dataIn2 = 32'd0; 
32'd3329: dataIn2 = 32'd0; 
32'd3330: dataIn2 = 32'd1; 
32'd3331: dataIn2 = 32'd0; 
32'd3332: dataIn2 = 32'd0; 
32'd3333: dataIn2 = 32'd1; 
32'd3334: dataIn2 = 32'd1; 
32'd3335: dataIn2 = 32'd1; 
32'd3336: dataIn2 = 32'd1; 
32'd3337: dataIn2 = 32'd1; 
32'd3338: dataIn2 = 32'd1; 
32'd3339: dataIn2 = 32'd0; 
32'd3340: dataIn2 = 32'd1; 
32'd3341: dataIn2 = 32'd1; 
32'd3342: dataIn2 = 32'd1; 
32'd3343: dataIn2 = 32'd1; 
32'd3344: dataIn2 = 32'd0; 
32'd3345: dataIn2 = 32'd0; 
32'd3346: dataIn2 = 32'd0; 
32'd3347: dataIn2 = 32'd1; 
32'd3348: dataIn2 = 32'd1; 
32'd3349: dataIn2 = 32'd0; 
32'd3350: dataIn2 = 32'd1; 
32'd3351: dataIn2 = 32'd0; 
32'd3352: dataIn2 = 32'd1; 
32'd3353: dataIn2 = 32'd1; 
32'd3354: dataIn2 = 32'd0; 
32'd3355: dataIn2 = 32'd1; 
32'd3356: dataIn2 = 32'd1; 
32'd3357: dataIn2 = 32'd0; 
32'd3358: dataIn2 = 32'd0; 
32'd3359: dataIn2 = 32'd0; 
32'd3360: dataIn2 = 32'd0; 
32'd3361: dataIn2 = 32'd1; 
32'd3362: dataIn2 = 32'd0; 
32'd3363: dataIn2 = 32'd0; 
32'd3364: dataIn2 = 32'd0; 
32'd3365: dataIn2 = 32'd1; 
32'd3366: dataIn2 = 32'd0; 
32'd3367: dataIn2 = 32'd1; 
32'd3368: dataIn2 = 32'd1; 
32'd3369: dataIn2 = 32'd1; 
32'd3370: dataIn2 = 32'd0; 
32'd3371: dataIn2 = 32'd0; 
32'd3372: dataIn2 = 32'd0; 
32'd3373: dataIn2 = 32'd1; 
32'd3374: dataIn2 = 32'd0; 
32'd3375: dataIn2 = 32'd0; 
32'd3376: dataIn2 = 32'd1; 
32'd3377: dataIn2 = 32'd1; 
32'd3378: dataIn2 = 32'd1; 
32'd3379: dataIn2 = 32'd0; 
32'd3380: dataIn2 = 32'd1; 
32'd3381: dataIn2 = 32'd0; 
32'd3382: dataIn2 = 32'd0; 
32'd3383: dataIn2 = 32'd1; 
32'd3384: dataIn2 = 32'd0; 
32'd3385: dataIn2 = 32'd0; 
32'd3386: dataIn2 = 32'd1; 
32'd3387: dataIn2 = 32'd1; 
32'd3388: dataIn2 = 32'd1; 
32'd3389: dataIn2 = 32'd1; 
32'd3390: dataIn2 = 32'd0; 
32'd3391: dataIn2 = 32'd0; 
32'd3392: dataIn2 = 32'd0; 
32'd3393: dataIn2 = 32'd1; 
32'd3394: dataIn2 = 32'd1; 
32'd3395: dataIn2 = 32'd1; 
32'd3396: dataIn2 = 32'd0; 
32'd3397: dataIn2 = 32'd0; 
32'd3398: dataIn2 = 32'd0; 
32'd3399: dataIn2 = 32'd0; 
32'd3400: dataIn2 = 32'd1; 
32'd3401: dataIn2 = 32'd0; 
32'd3402: dataIn2 = 32'd0; 
32'd3403: dataIn2 = 32'd0; 
32'd3404: dataIn2 = 32'd0; 
32'd3405: dataIn2 = 32'd0; 
32'd3406: dataIn2 = 32'd1; 
32'd3407: dataIn2 = 32'd0; 
32'd3408: dataIn2 = 32'd1; 
32'd3409: dataIn2 = 32'd0; 
32'd3410: dataIn2 = 32'd0; 
32'd3411: dataIn2 = 32'd1; 
32'd3412: dataIn2 = 32'd0; 
32'd3413: dataIn2 = 32'd1; 
32'd3414: dataIn2 = 32'd0; 
32'd3415: dataIn2 = 32'd0; 
32'd3416: dataIn2 = 32'd1; 
32'd3417: dataIn2 = 32'd0; 
32'd3418: dataIn2 = 32'd1; 
32'd3419: dataIn2 = 32'd0; 
32'd3420: dataIn2 = 32'd1; 
32'd3421: dataIn2 = 32'd0; 
32'd3422: dataIn2 = 32'd1; 
32'd3423: dataIn2 = 32'd1; 
32'd3424: dataIn2 = 32'd0; 
32'd3425: dataIn2 = 32'd1; 
32'd3426: dataIn2 = 32'd1; 
32'd3427: dataIn2 = 32'd0; 
32'd3428: dataIn2 = 32'd0; 
32'd3429: dataIn2 = 32'd0; 
32'd3430: dataIn2 = 32'd0; 
32'd3431: dataIn2 = 32'd0; 
32'd3432: dataIn2 = 32'd1; 
32'd3433: dataIn2 = 32'd0; 
32'd3434: dataIn2 = 32'd0; 
32'd3435: dataIn2 = 32'd0; 
32'd3436: dataIn2 = 32'd1; 
32'd3437: dataIn2 = 32'd1; 
32'd3438: dataIn2 = 32'd0; 
32'd3439: dataIn2 = 32'd1; 
32'd3440: dataIn2 = 32'd0; 
32'd3441: dataIn2 = 32'd1; 
32'd3442: dataIn2 = 32'd0; 
32'd3443: dataIn2 = 32'd1; 
32'd3444: dataIn2 = 32'd1; 
32'd3445: dataIn2 = 32'd0; 
32'd3446: dataIn2 = 32'd0; 
32'd3447: dataIn2 = 32'd0; 
32'd3448: dataIn2 = 32'd1; 
32'd3449: dataIn2 = 32'd0; 
32'd3450: dataIn2 = 32'd0; 
32'd3451: dataIn2 = 32'd1; 
32'd3452: dataIn2 = 32'd1; 
32'd3453: dataIn2 = 32'd0; 
32'd3454: dataIn2 = 32'd0; 
32'd3455: dataIn2 = 32'd1; 
32'd3456: dataIn2 = 32'd1; 
32'd3457: dataIn2 = 32'd0; 
32'd3458: dataIn2 = 32'd1; 
32'd3459: dataIn2 = 32'd1; 
32'd3460: dataIn2 = 32'd1; 
32'd3461: dataIn2 = 32'd0; 
32'd3462: dataIn2 = 32'd0; 
32'd3463: dataIn2 = 32'd0; 
32'd3464: dataIn2 = 32'd0; 
32'd3465: dataIn2 = 32'd1; 
32'd3466: dataIn2 = 32'd1; 
32'd3467: dataIn2 = 32'd1; 
32'd3468: dataIn2 = 32'd1; 
32'd3469: dataIn2 = 32'd0; 
32'd3470: dataIn2 = 32'd1; 
32'd3471: dataIn2 = 32'd0; 
32'd3472: dataIn2 = 32'd0; 
32'd3473: dataIn2 = 32'd1; 
32'd3474: dataIn2 = 32'd0; 
32'd3475: dataIn2 = 32'd0; 
32'd3476: dataIn2 = 32'd1; 
32'd3477: dataIn2 = 32'd0; 
32'd3478: dataIn2 = 32'd0; 
32'd3479: dataIn2 = 32'd0; 
32'd3480: dataIn2 = 32'd1; 
32'd3481: dataIn2 = 32'd1; 
32'd3482: dataIn2 = 32'd0; 
32'd3483: dataIn2 = 32'd0; 
32'd3484: dataIn2 = 32'd0; 
32'd3485: dataIn2 = 32'd1; 
32'd3486: dataIn2 = 32'd1; 
32'd3487: dataIn2 = 32'd1; 
32'd3488: dataIn2 = 32'd1; 
32'd3489: dataIn2 = 32'd1; 
32'd3490: dataIn2 = 32'd0; 
32'd3491: dataIn2 = 32'd1; 
32'd3492: dataIn2 = 32'd1; 
32'd3493: dataIn2 = 32'd1; 
32'd3494: dataIn2 = 32'd1; 
32'd3495: dataIn2 = 32'd1; 
32'd3496: dataIn2 = 32'd0; 
32'd3497: dataIn2 = 32'd0; 
32'd3498: dataIn2 = 32'd1; 
32'd3499: dataIn2 = 32'd1; 
32'd3500: dataIn2 = 32'd0; 
32'd3501: dataIn2 = 32'd1; 
32'd3502: dataIn2 = 32'd0; 
32'd3503: dataIn2 = 32'd1; 
32'd3504: dataIn2 = 32'd1; 
32'd3505: dataIn2 = 32'd0; 
32'd3506: dataIn2 = 32'd0; 
32'd3507: dataIn2 = 32'd0; 
32'd3508: dataIn2 = 32'd1; 
32'd3509: dataIn2 = 32'd0; 
32'd3510: dataIn2 = 32'd0; 
32'd3511: dataIn2 = 32'd1; 
32'd3512: dataIn2 = 32'd0; 
32'd3513: dataIn2 = 32'd0; 
32'd3514: dataIn2 = 32'd0; 
32'd3515: dataIn2 = 32'd1; 
32'd3516: dataIn2 = 32'd0; 
32'd3517: dataIn2 = 32'd0; 
32'd3518: dataIn2 = 32'd1; 
32'd3519: dataIn2 = 32'd0; 
32'd3520: dataIn2 = 32'd1; 
32'd3521: dataIn2 = 32'd0; 
32'd3522: dataIn2 = 32'd0; 
32'd3523: dataIn2 = 32'd0; 
32'd3524: dataIn2 = 32'd0; 
32'd3525: dataIn2 = 32'd0; 
32'd3526: dataIn2 = 32'd1; 
32'd3527: dataIn2 = 32'd1; 
32'd3528: dataIn2 = 32'd0; 
32'd3529: dataIn2 = 32'd1; 
32'd3530: dataIn2 = 32'd1; 
32'd3531: dataIn2 = 32'd1; 
32'd3532: dataIn2 = 32'd1; 
32'd3533: dataIn2 = 32'd0; 
32'd3534: dataIn2 = 32'd1; 
32'd3535: dataIn2 = 32'd0; 
32'd3536: dataIn2 = 32'd0; 
32'd3537: dataIn2 = 32'd0; 
32'd3538: dataIn2 = 32'd0; 
32'd3539: dataIn2 = 32'd0; 
32'd3540: dataIn2 = 32'd1; 
32'd3541: dataIn2 = 32'd0; 
32'd3542: dataIn2 = 32'd1; 
32'd3543: dataIn2 = 32'd1; 
32'd3544: dataIn2 = 32'd1; 
32'd3545: dataIn2 = 32'd1; 
32'd3546: dataIn2 = 32'd1; 
32'd3547: dataIn2 = 32'd1; 
32'd3548: dataIn2 = 32'd0; 
32'd3549: dataIn2 = 32'd0; 
32'd3550: dataIn2 = 32'd1; 
32'd3551: dataIn2 = 32'd0; 
32'd3552: dataIn2 = 32'd1; 
32'd3553: dataIn2 = 32'd0; 
32'd3554: dataIn2 = 32'd0; 
32'd3555: dataIn2 = 32'd0; 
32'd3556: dataIn2 = 32'd1; 
32'd3557: dataIn2 = 32'd0; 
32'd3558: dataIn2 = 32'd1; 
32'd3559: dataIn2 = 32'd1; 
32'd3560: dataIn2 = 32'd0; 
32'd3561: dataIn2 = 32'd1; 
32'd3562: dataIn2 = 32'd0; 
32'd3563: dataIn2 = 32'd0; 
32'd3564: dataIn2 = 32'd1; 
32'd3565: dataIn2 = 32'd1; 
32'd3566: dataIn2 = 32'd0; 
32'd3567: dataIn2 = 32'd1; 
32'd3568: dataIn2 = 32'd0; 
32'd3569: dataIn2 = 32'd0; 
32'd3570: dataIn2 = 32'd0; 
32'd3571: dataIn2 = 32'd1; 
32'd3572: dataIn2 = 32'd0; 
32'd3573: dataIn2 = 32'd1; 
32'd3574: dataIn2 = 32'd1; 
32'd3575: dataIn2 = 32'd0; 
32'd3576: dataIn2 = 32'd1; 
32'd3577: dataIn2 = 32'd1; 
32'd3578: dataIn2 = 32'd1; 
32'd3579: dataIn2 = 32'd1; 
32'd3580: dataIn2 = 32'd0; 
32'd3581: dataIn2 = 32'd0; 
32'd3582: dataIn2 = 32'd0; 
32'd3583: dataIn2 = 32'd0; 
32'd3584: dataIn2 = 32'd1; 
32'd3585: dataIn2 = 32'd1; 
32'd3586: dataIn2 = 32'd1; 
32'd3587: dataIn2 = 32'd0; 
32'd3588: dataIn2 = 32'd0; 
32'd3589: dataIn2 = 32'd0; 
32'd3590: dataIn2 = 32'd0; 
32'd3591: dataIn2 = 32'd0; 
32'd3592: dataIn2 = 32'd1; 
32'd3593: dataIn2 = 32'd0; 
32'd3594: dataIn2 = 32'd0; 
32'd3595: dataIn2 = 32'd1; 
32'd3596: dataIn2 = 32'd1; 
32'd3597: dataIn2 = 32'd1; 
32'd3598: dataIn2 = 32'd0; 
32'd3599: dataIn2 = 32'd0; 
32'd3600: dataIn2 = 32'd1; 
32'd3601: dataIn2 = 32'd0; 
32'd3602: dataIn2 = 32'd0; 
32'd3603: dataIn2 = 32'd0; 
32'd3604: dataIn2 = 32'd0; 
32'd3605: dataIn2 = 32'd0; 
32'd3606: dataIn2 = 32'd0; 
32'd3607: dataIn2 = 32'd0; 
32'd3608: dataIn2 = 32'd1; 
32'd3609: dataIn2 = 32'd1; 
32'd3610: dataIn2 = 32'd1; 
32'd3611: dataIn2 = 32'd1; 
32'd3612: dataIn2 = 32'd1; 
32'd3613: dataIn2 = 32'd1; 
32'd3614: dataIn2 = 32'd1; 
32'd3615: dataIn2 = 32'd0; 
32'd3616: dataIn2 = 32'd0; 
32'd3617: dataIn2 = 32'd0; 
32'd3618: dataIn2 = 32'd1; 
32'd3619: dataIn2 = 32'd1; 
32'd3620: dataIn2 = 32'd0; 
32'd3621: dataIn2 = 32'd1; 
32'd3622: dataIn2 = 32'd1; 
32'd3623: dataIn2 = 32'd1; 
32'd3624: dataIn2 = 32'd0; 
32'd3625: dataIn2 = 32'd1; 
32'd3626: dataIn2 = 32'd1; 
32'd3627: dataIn2 = 32'd0; 
32'd3628: dataIn2 = 32'd1; 
32'd3629: dataIn2 = 32'd1; 
32'd3630: dataIn2 = 32'd1; 
32'd3631: dataIn2 = 32'd1; 
32'd3632: dataIn2 = 32'd0; 
32'd3633: dataIn2 = 32'd0; 
32'd3634: dataIn2 = 32'd0; 
32'd3635: dataIn2 = 32'd0; 
32'd3636: dataIn2 = 32'd0; 
32'd3637: dataIn2 = 32'd1; 
32'd3638: dataIn2 = 32'd0; 
32'd3639: dataIn2 = 32'd1; 
32'd3640: dataIn2 = 32'd1; 
32'd3641: dataIn2 = 32'd0; 
32'd3642: dataIn2 = 32'd1; 
32'd3643: dataIn2 = 32'd0; 
32'd3644: dataIn2 = 32'd1; 
32'd3645: dataIn2 = 32'd1; 
32'd3646: dataIn2 = 32'd1; 
32'd3647: dataIn2 = 32'd0; 
32'd3648: dataIn2 = 32'd0; 
32'd3649: dataIn2 = 32'd1; 
32'd3650: dataIn2 = 32'd1; 
32'd3651: dataIn2 = 32'd1; 
32'd3652: dataIn2 = 32'd0; 
32'd3653: dataIn2 = 32'd0; 
32'd3654: dataIn2 = 32'd0; 
32'd3655: dataIn2 = 32'd1; 
32'd3656: dataIn2 = 32'd1; 
32'd3657: dataIn2 = 32'd0; 
32'd3658: dataIn2 = 32'd0; 
32'd3659: dataIn2 = 32'd0; 
32'd3660: dataIn2 = 32'd1; 
32'd3661: dataIn2 = 32'd1; 
32'd3662: dataIn2 = 32'd1; 
32'd3663: dataIn2 = 32'd0; 
32'd3664: dataIn2 = 32'd0; 
32'd3665: dataIn2 = 32'd0; 
32'd3666: dataIn2 = 32'd1; 
32'd3667: dataIn2 = 32'd1; 
32'd3668: dataIn2 = 32'd0; 
32'd3669: dataIn2 = 32'd1; 
32'd3670: dataIn2 = 32'd0; 
32'd3671: dataIn2 = 32'd1; 
32'd3672: dataIn2 = 32'd1; 
32'd3673: dataIn2 = 32'd0; 
32'd3674: dataIn2 = 32'd1; 
32'd3675: dataIn2 = 32'd1; 
32'd3676: dataIn2 = 32'd1; 
32'd3677: dataIn2 = 32'd0; 
32'd3678: dataIn2 = 32'd0; 
32'd3679: dataIn2 = 32'd0; 
32'd3680: dataIn2 = 32'd1; 
32'd3681: dataIn2 = 32'd1; 
32'd3682: dataIn2 = 32'd1; 
32'd3683: dataIn2 = 32'd0; 
32'd3684: dataIn2 = 32'd0; 
32'd3685: dataIn2 = 32'd0; 
32'd3686: dataIn2 = 32'd1; 
32'd3687: dataIn2 = 32'd0; 
32'd3688: dataIn2 = 32'd0; 
32'd3689: dataIn2 = 32'd1; 
32'd3690: dataIn2 = 32'd1; 
32'd3691: dataIn2 = 32'd0; 
32'd3692: dataIn2 = 32'd1; 
32'd3693: dataIn2 = 32'd1; 
32'd3694: dataIn2 = 32'd0; 
32'd3695: dataIn2 = 32'd1; 
32'd3696: dataIn2 = 32'd0; 
32'd3697: dataIn2 = 32'd1; 
32'd3698: dataIn2 = 32'd0; 
32'd3699: dataIn2 = 32'd0; 
32'd3700: dataIn2 = 32'd1; 
32'd3701: dataIn2 = 32'd0; 
32'd3702: dataIn2 = 32'd1; 
32'd3703: dataIn2 = 32'd0; 
32'd3704: dataIn2 = 32'd1; 
32'd3705: dataIn2 = 32'd1; 
32'd3706: dataIn2 = 32'd0; 
32'd3707: dataIn2 = 32'd0; 
32'd3708: dataIn2 = 32'd0; 
32'd3709: dataIn2 = 32'd1; 
32'd3710: dataIn2 = 32'd1; 
32'd3711: dataIn2 = 32'd1; 
32'd3712: dataIn2 = 32'd0; 
32'd3713: dataIn2 = 32'd0; 
32'd3714: dataIn2 = 32'd0; 
32'd3715: dataIn2 = 32'd1; 
32'd3716: dataIn2 = 32'd0; 
32'd3717: dataIn2 = 32'd0; 
32'd3718: dataIn2 = 32'd0; 
32'd3719: dataIn2 = 32'd1; 
32'd3720: dataIn2 = 32'd1; 
32'd3721: dataIn2 = 32'd1; 
32'd3722: dataIn2 = 32'd1; 
32'd3723: dataIn2 = 32'd1; 
32'd3724: dataIn2 = 32'd1; 
32'd3725: dataIn2 = 32'd0; 
32'd3726: dataIn2 = 32'd0; 
32'd3727: dataIn2 = 32'd1; 
32'd3728: dataIn2 = 32'd1; 
32'd3729: dataIn2 = 32'd1; 
32'd3730: dataIn2 = 32'd0; 
32'd3731: dataIn2 = 32'd0; 
32'd3732: dataIn2 = 32'd1; 
32'd3733: dataIn2 = 32'd1; 
32'd3734: dataIn2 = 32'd1; 
32'd3735: dataIn2 = 32'd1; 
32'd3736: dataIn2 = 32'd0; 
32'd3737: dataIn2 = 32'd0; 
32'd3738: dataIn2 = 32'd1; 
32'd3739: dataIn2 = 32'd0; 
32'd3740: dataIn2 = 32'd1; 
32'd3741: dataIn2 = 32'd0; 
32'd3742: dataIn2 = 32'd1; 
32'd3743: dataIn2 = 32'd1; 
32'd3744: dataIn2 = 32'd1; 
32'd3745: dataIn2 = 32'd0; 
32'd3746: dataIn2 = 32'd0; 
32'd3747: dataIn2 = 32'd1; 
32'd3748: dataIn2 = 32'd1; 
32'd3749: dataIn2 = 32'd1; 
32'd3750: dataIn2 = 32'd1; 
32'd3751: dataIn2 = 32'd1; 
32'd3752: dataIn2 = 32'd1; 
32'd3753: dataIn2 = 32'd1; 
32'd3754: dataIn2 = 32'd1; 
32'd3755: dataIn2 = 32'd0; 
32'd3756: dataIn2 = 32'd0; 
32'd3757: dataIn2 = 32'd0; 
32'd3758: dataIn2 = 32'd1; 
32'd3759: dataIn2 = 32'd0; 
32'd3760: dataIn2 = 32'd1; 
32'd3761: dataIn2 = 32'd1; 
32'd3762: dataIn2 = 32'd1; 
32'd3763: dataIn2 = 32'd0; 
32'd3764: dataIn2 = 32'd1; 
32'd3765: dataIn2 = 32'd0; 
32'd3766: dataIn2 = 32'd1; 
32'd3767: dataIn2 = 32'd1; 
32'd3768: dataIn2 = 32'd0; 
32'd3769: dataIn2 = 32'd0; 
32'd3770: dataIn2 = 32'd1; 
32'd3771: dataIn2 = 32'd0; 
32'd3772: dataIn2 = 32'd0; 
32'd3773: dataIn2 = 32'd1; 
32'd3774: dataIn2 = 32'd1; 
32'd3775: dataIn2 = 32'd0; 
32'd3776: dataIn2 = 32'd0; 
32'd3777: dataIn2 = 32'd0; 
32'd3778: dataIn2 = 32'd1; 
32'd3779: dataIn2 = 32'd0; 
32'd3780: dataIn2 = 32'd1; 
32'd3781: dataIn2 = 32'd1; 
32'd3782: dataIn2 = 32'd0; 
32'd3783: dataIn2 = 32'd1; 
32'd3784: dataIn2 = 32'd1; 
32'd3785: dataIn2 = 32'd0; 
32'd3786: dataIn2 = 32'd1; 
32'd3787: dataIn2 = 32'd0; 
32'd3788: dataIn2 = 32'd1; 
32'd3789: dataIn2 = 32'd1; 
32'd3790: dataIn2 = 32'd1; 
32'd3791: dataIn2 = 32'd1; 
32'd3792: dataIn2 = 32'd1; 
32'd3793: dataIn2 = 32'd0; 
32'd3794: dataIn2 = 32'd1; 
32'd3795: dataIn2 = 32'd1; 
32'd3796: dataIn2 = 32'd0; 
32'd3797: dataIn2 = 32'd1; 
32'd3798: dataIn2 = 32'd1; 
32'd3799: dataIn2 = 32'd0; 
32'd3800: dataIn2 = 32'd1; 
32'd3801: dataIn2 = 32'd0; 
32'd3802: dataIn2 = 32'd1; 
32'd3803: dataIn2 = 32'd1; 
32'd3804: dataIn2 = 32'd1; 
32'd3805: dataIn2 = 32'd1; 
32'd3806: dataIn2 = 32'd1; 
32'd3807: dataIn2 = 32'd0; 
32'd3808: dataIn2 = 32'd0; 
32'd3809: dataIn2 = 32'd0; 
32'd3810: dataIn2 = 32'd1; 
32'd3811: dataIn2 = 32'd1; 
32'd3812: dataIn2 = 32'd0; 
32'd3813: dataIn2 = 32'd0; 
32'd3814: dataIn2 = 32'd0; 
32'd3815: dataIn2 = 32'd0; 
32'd3816: dataIn2 = 32'd0; 
32'd3817: dataIn2 = 32'd0; 
32'd3818: dataIn2 = 32'd0; 
32'd3819: dataIn2 = 32'd0; 
32'd3820: dataIn2 = 32'd1; 
32'd3821: dataIn2 = 32'd1; 
32'd3822: dataIn2 = 32'd0; 
32'd3823: dataIn2 = 32'd1; 
32'd3824: dataIn2 = 32'd1; 
32'd3825: dataIn2 = 32'd1; 
32'd3826: dataIn2 = 32'd1; 
32'd3827: dataIn2 = 32'd1; 
32'd3828: dataIn2 = 32'd1; 
32'd3829: dataIn2 = 32'd0; 
32'd3830: dataIn2 = 32'd1; 
32'd3831: dataIn2 = 32'd1; 
32'd3832: dataIn2 = 32'd1; 
32'd3833: dataIn2 = 32'd1; 
32'd3834: dataIn2 = 32'd1; 
32'd3835: dataIn2 = 32'd0; 
32'd3836: dataIn2 = 32'd0; 
32'd3837: dataIn2 = 32'd1; 
32'd3838: dataIn2 = 32'd0; 
32'd3839: dataIn2 = 32'd1; 
32'd3840: dataIn2 = 32'd0; 
32'd3841: dataIn2 = 32'd1; 
32'd3842: dataIn2 = 32'd1; 
32'd3843: dataIn2 = 32'd1; 
32'd3844: dataIn2 = 32'd0; 
32'd3845: dataIn2 = 32'd0; 
32'd3846: dataIn2 = 32'd0; 
32'd3847: dataIn2 = 32'd0; 
32'd3848: dataIn2 = 32'd0; 
32'd3849: dataIn2 = 32'd1; 
32'd3850: dataIn2 = 32'd0; 
32'd3851: dataIn2 = 32'd1; 
32'd3852: dataIn2 = 32'd1; 
32'd3853: dataIn2 = 32'd0; 
32'd3854: dataIn2 = 32'd0; 
32'd3855: dataIn2 = 32'd1; 
32'd3856: dataIn2 = 32'd1; 
32'd3857: dataIn2 = 32'd1; 
32'd3858: dataIn2 = 32'd1; 
32'd3859: dataIn2 = 32'd1; 
32'd3860: dataIn2 = 32'd0; 
32'd3861: dataIn2 = 32'd0; 
32'd3862: dataIn2 = 32'd1; 
32'd3863: dataIn2 = 32'd1; 
32'd3864: dataIn2 = 32'd1; 
32'd3865: dataIn2 = 32'd1; 
32'd3866: dataIn2 = 32'd1; 
32'd3867: dataIn2 = 32'd1; 
32'd3868: dataIn2 = 32'd1; 
32'd3869: dataIn2 = 32'd1; 
32'd3870: dataIn2 = 32'd0; 
32'd3871: dataIn2 = 32'd1; 
32'd3872: dataIn2 = 32'd0; 
32'd3873: dataIn2 = 32'd1; 
32'd3874: dataIn2 = 32'd0; 
32'd3875: dataIn2 = 32'd1; 
32'd3876: dataIn2 = 32'd1; 
32'd3877: dataIn2 = 32'd1; 
32'd3878: dataIn2 = 32'd0; 
32'd3879: dataIn2 = 32'd1; 
32'd3880: dataIn2 = 32'd1; 
32'd3881: dataIn2 = 32'd0; 
32'd3882: dataIn2 = 32'd0; 
32'd3883: dataIn2 = 32'd1; 
32'd3884: dataIn2 = 32'd0; 
32'd3885: dataIn2 = 32'd1; 
32'd3886: dataIn2 = 32'd1; 
32'd3887: dataIn2 = 32'd0; 
32'd3888: dataIn2 = 32'd1; 
32'd3889: dataIn2 = 32'd0; 
32'd3890: dataIn2 = 32'd1; 
32'd3891: dataIn2 = 32'd1; 
32'd3892: dataIn2 = 32'd1; 
32'd3893: dataIn2 = 32'd0; 
32'd3894: dataIn2 = 32'd0; 
32'd3895: dataIn2 = 32'd1; 
32'd3896: dataIn2 = 32'd1; 
32'd3897: dataIn2 = 32'd1; 
32'd3898: dataIn2 = 32'd1; 
32'd3899: dataIn2 = 32'd0; 
32'd3900: dataIn2 = 32'd0; 
32'd3901: dataIn2 = 32'd1; 
32'd3902: dataIn2 = 32'd1; 
32'd3903: dataIn2 = 32'd1; 
32'd3904: dataIn2 = 32'd0; 
32'd3905: dataIn2 = 32'd1; 
32'd3906: dataIn2 = 32'd1; 
32'd3907: dataIn2 = 32'd1; 
32'd3908: dataIn2 = 32'd0; 
32'd3909: dataIn2 = 32'd1; 
32'd3910: dataIn2 = 32'd0; 
32'd3911: dataIn2 = 32'd1; 
32'd3912: dataIn2 = 32'd0; 
32'd3913: dataIn2 = 32'd1; 
32'd3914: dataIn2 = 32'd0; 
32'd3915: dataIn2 = 32'd1; 
32'd3916: dataIn2 = 32'd0; 
32'd3917: dataIn2 = 32'd0; 
32'd3918: dataIn2 = 32'd0; 
32'd3919: dataIn2 = 32'd1; 
32'd3920: dataIn2 = 32'd1; 
32'd3921: dataIn2 = 32'd0; 
32'd3922: dataIn2 = 32'd0; 
32'd3923: dataIn2 = 32'd0; 
32'd3924: dataIn2 = 32'd0; 
32'd3925: dataIn2 = 32'd1; 
32'd3926: dataIn2 = 32'd0; 
32'd3927: dataIn2 = 32'd1; 
32'd3928: dataIn2 = 32'd0; 
32'd3929: dataIn2 = 32'd0; 
32'd3930: dataIn2 = 32'd0; 
32'd3931: dataIn2 = 32'd1; 
32'd3932: dataIn2 = 32'd1; 
32'd3933: dataIn2 = 32'd0; 
32'd3934: dataIn2 = 32'd0; 
32'd3935: dataIn2 = 32'd0; 
32'd3936: dataIn2 = 32'd0; 
32'd3937: dataIn2 = 32'd1; 
32'd3938: dataIn2 = 32'd1; 
32'd3939: dataIn2 = 32'd0; 
32'd3940: dataIn2 = 32'd0; 
32'd3941: dataIn2 = 32'd1; 
32'd3942: dataIn2 = 32'd1; 
32'd3943: dataIn2 = 32'd0; 
32'd3944: dataIn2 = 32'd1; 
32'd3945: dataIn2 = 32'd1; 
32'd3946: dataIn2 = 32'd1; 
32'd3947: dataIn2 = 32'd0; 
32'd3948: dataIn2 = 32'd1; 
32'd3949: dataIn2 = 32'd1; 
32'd3950: dataIn2 = 32'd0; 
32'd3951: dataIn2 = 32'd0; 
32'd3952: dataIn2 = 32'd0; 
32'd3953: dataIn2 = 32'd1; 
32'd3954: dataIn2 = 32'd1; 
32'd3955: dataIn2 = 32'd0; 
32'd3956: dataIn2 = 32'd0; 
32'd3957: dataIn2 = 32'd0; 
32'd3958: dataIn2 = 32'd1; 
32'd3959: dataIn2 = 32'd0; 
32'd3960: dataIn2 = 32'd0; 
32'd3961: dataIn2 = 32'd0; 
32'd3962: dataIn2 = 32'd1; 
32'd3963: dataIn2 = 32'd0; 
32'd3964: dataIn2 = 32'd0; 
32'd3965: dataIn2 = 32'd1; 
32'd3966: dataIn2 = 32'd0; 
32'd3967: dataIn2 = 32'd1; 
32'd3968: dataIn2 = 32'd1; 
32'd3969: dataIn2 = 32'd1; 
32'd3970: dataIn2 = 32'd1; 
32'd3971: dataIn2 = 32'd1; 
32'd3972: dataIn2 = 32'd0; 
32'd3973: dataIn2 = 32'd0; 
32'd3974: dataIn2 = 32'd0; 
32'd3975: dataIn2 = 32'd1; 
32'd3976: dataIn2 = 32'd0; 
32'd3977: dataIn2 = 32'd1; 
32'd3978: dataIn2 = 32'd0; 
32'd3979: dataIn2 = 32'd0; 
32'd3980: dataIn2 = 32'd0; 
32'd3981: dataIn2 = 32'd1; 
32'd3982: dataIn2 = 32'd0; 
32'd3983: dataIn2 = 32'd1; 
32'd3984: dataIn2 = 32'd1; 
32'd3985: dataIn2 = 32'd0; 
32'd3986: dataIn2 = 32'd1; 
32'd3987: dataIn2 = 32'd1; 
32'd3988: dataIn2 = 32'd1; 
32'd3989: dataIn2 = 32'd0; 
32'd3990: dataIn2 = 32'd0; 
32'd3991: dataIn2 = 32'd1; 
32'd3992: dataIn2 = 32'd1; 
32'd3993: dataIn2 = 32'd0; 
32'd3994: dataIn2 = 32'd1; 
32'd3995: dataIn2 = 32'd1; 
32'd3996: dataIn2 = 32'd0; 
32'd3997: dataIn2 = 32'd1; 
32'd3998: dataIn2 = 32'd1; 
32'd3999: dataIn2 = 32'd1; 
32'd4000: dataIn2 = 32'd0; 
32'd4001: dataIn2 = 32'd1; 
32'd4002: dataIn2 = 32'd0; 
32'd4003: dataIn2 = 32'd1; 
32'd4004: dataIn2 = 32'd0; 
32'd4005: dataIn2 = 32'd0; 
32'd4006: dataIn2 = 32'd0; 
32'd4007: dataIn2 = 32'd1; 
32'd4008: dataIn2 = 32'd1; 
32'd4009: dataIn2 = 32'd0; 
32'd4010: dataIn2 = 32'd1; 
32'd4011: dataIn2 = 32'd0; 
32'd4012: dataIn2 = 32'd0; 
32'd4013: dataIn2 = 32'd1; 
32'd4014: dataIn2 = 32'd0; 
32'd4015: dataIn2 = 32'd1; 
32'd4016: dataIn2 = 32'd1; 
32'd4017: dataIn2 = 32'd0; 
32'd4018: dataIn2 = 32'd1; 
32'd4019: dataIn2 = 32'd1; 
32'd4020: dataIn2 = 32'd0; 
32'd4021: dataIn2 = 32'd0; 
32'd4022: dataIn2 = 32'd1; 
32'd4023: dataIn2 = 32'd1; 
32'd4024: dataIn2 = 32'd1; 
32'd4025: dataIn2 = 32'd1; 
32'd4026: dataIn2 = 32'd1; 
32'd4027: dataIn2 = 32'd1; 
32'd4028: dataIn2 = 32'd0; 
32'd4029: dataIn2 = 32'd1; 
32'd4030: dataIn2 = 32'd0; 
32'd4031: dataIn2 = 32'd1; 
32'd4032: dataIn2 = 32'd0; 
32'd4033: dataIn2 = 32'd0; 
32'd4034: dataIn2 = 32'd0; 
32'd4035: dataIn2 = 32'd1; 
32'd4036: dataIn2 = 32'd1; 
32'd4037: dataIn2 = 32'd1; 
32'd4038: dataIn2 = 32'd0; 
32'd4039: dataIn2 = 32'd0; 
32'd4040: dataIn2 = 32'd0; 
32'd4041: dataIn2 = 32'd0; 
32'd4042: dataIn2 = 32'd0; 
32'd4043: dataIn2 = 32'd1; 
32'd4044: dataIn2 = 32'd1; 
32'd4045: dataIn2 = 32'd0; 
32'd4046: dataIn2 = 32'd1; 
32'd4047: dataIn2 = 32'd1; 
32'd4048: dataIn2 = 32'd1; 
32'd4049: dataIn2 = 32'd0; 
32'd4050: dataIn2 = 32'd0; 
32'd4051: dataIn2 = 32'd1; 
32'd4052: dataIn2 = 32'd0; 
32'd4053: dataIn2 = 32'd1; 
32'd4054: dataIn2 = 32'd0; 
32'd4055: dataIn2 = 32'd1; 
32'd4056: dataIn2 = 32'd1; 
32'd4057: dataIn2 = 32'd1; 
32'd4058: dataIn2 = 32'd1; 
32'd4059: dataIn2 = 32'd0; 
32'd4060: dataIn2 = 32'd1; 
32'd4061: dataIn2 = 32'd1; 
32'd4062: dataIn2 = 32'd1; 
32'd4063: dataIn2 = 32'd0; 
32'd4064: dataIn2 = 32'd0; 
32'd4065: dataIn2 = 32'd1; 
32'd4066: dataIn2 = 32'd1; 
32'd4067: dataIn2 = 32'd0; 
32'd4068: dataIn2 = 32'd0; 
32'd4069: dataIn2 = 32'd0; 
32'd4070: dataIn2 = 32'd0; 
32'd4071: dataIn2 = 32'd1; 
32'd4072: dataIn2 = 32'd1; 
32'd4073: dataIn2 = 32'd1; 
32'd4074: dataIn2 = 32'd0; 
32'd4075: dataIn2 = 32'd1; 
32'd4076: dataIn2 = 32'd1; 
32'd4077: dataIn2 = 32'd1; 
32'd4078: dataIn2 = 32'd0; 
32'd4079: dataIn2 = 32'd0; 
32'd4080: dataIn2 = 32'd1; 
32'd4081: dataIn2 = 32'd1; 
32'd4082: dataIn2 = 32'd1; 
32'd4083: dataIn2 = 32'd1; 
32'd4084: dataIn2 = 32'd1; 
32'd4085: dataIn2 = 32'd1; 
32'd4086: dataIn2 = 32'd0; 
32'd4087: dataIn2 = 32'd1; 
32'd4088: dataIn2 = 32'd1; 
32'd4089: dataIn2 = 32'd1; 
32'd4090: dataIn2 = 32'd0; 
32'd4091: dataIn2 = 32'd1; 
32'd4092: dataIn2 = 32'd1; 
32'd4093: dataIn2 = 32'd0; 
32'd4094: dataIn2 = 32'd0; 
32'd4095: dataIn2 = 32'd1; 
32'd4096: dataIn2 = 32'd0; 
32'd4097: dataIn2 = 32'd0; 
32'd4098: dataIn2 = 32'd0; 
32'd4099: dataIn2 = 32'd1; 
32'd4100: dataIn2 = 32'd1; 
32'd4101: dataIn2 = 32'd0; 
32'd4102: dataIn2 = 32'd1; 
32'd4103: dataIn2 = 32'd0; 
32'd4104: dataIn2 = 32'd0; 
32'd4105: dataIn2 = 32'd0; 
32'd4106: dataIn2 = 32'd1; 
32'd4107: dataIn2 = 32'd1; 
32'd4108: dataIn2 = 32'd0; 
32'd4109: dataIn2 = 32'd0; 
32'd4110: dataIn2 = 32'd1; 
32'd4111: dataIn2 = 32'd1; 
32'd4112: dataIn2 = 32'd0; 
32'd4113: dataIn2 = 32'd0; 
32'd4114: dataIn2 = 32'd0; 
32'd4115: dataIn2 = 32'd0; 
32'd4116: dataIn2 = 32'd1; 
32'd4117: dataIn2 = 32'd1; 
32'd4118: dataIn2 = 32'd0; 
32'd4119: dataIn2 = 32'd0; 
32'd4120: dataIn2 = 32'd1; 
32'd4121: dataIn2 = 32'd0; 
32'd4122: dataIn2 = 32'd0; 
32'd4123: dataIn2 = 32'd1; 
32'd4124: dataIn2 = 32'd1; 
32'd4125: dataIn2 = 32'd1; 
32'd4126: dataIn2 = 32'd0; 
32'd4127: dataIn2 = 32'd0; 
32'd4128: dataIn2 = 32'd0; 
32'd4129: dataIn2 = 32'd1; 
32'd4130: dataIn2 = 32'd0; 
32'd4131: dataIn2 = 32'd1; 
32'd4132: dataIn2 = 32'd1; 
32'd4133: dataIn2 = 32'd0; 
32'd4134: dataIn2 = 32'd1; 
32'd4135: dataIn2 = 32'd0; 
32'd4136: dataIn2 = 32'd0; 
32'd4137: dataIn2 = 32'd1; 
32'd4138: dataIn2 = 32'd0; 
32'd4139: dataIn2 = 32'd1; 
32'd4140: dataIn2 = 32'd1; 
32'd4141: dataIn2 = 32'd0; 
32'd4142: dataIn2 = 32'd1; 
32'd4143: dataIn2 = 32'd0; 
32'd4144: dataIn2 = 32'd1; 
32'd4145: dataIn2 = 32'd1; 
32'd4146: dataIn2 = 32'd0; 
32'd4147: dataIn2 = 32'd0; 
32'd4148: dataIn2 = 32'd0; 
32'd4149: dataIn2 = 32'd1; 
32'd4150: dataIn2 = 32'd1; 
32'd4151: dataIn2 = 32'd0; 
32'd4152: dataIn2 = 32'd0; 
32'd4153: dataIn2 = 32'd1; 
32'd4154: dataIn2 = 32'd0; 
32'd4155: dataIn2 = 32'd0; 
32'd4156: dataIn2 = 32'd0; 
32'd4157: dataIn2 = 32'd0; 
32'd4158: dataIn2 = 32'd1; 
32'd4159: dataIn2 = 32'd0; 
32'd4160: dataIn2 = 32'd1; 
32'd4161: dataIn2 = 32'd1; 
32'd4162: dataIn2 = 32'd0; 
32'd4163: dataIn2 = 32'd1; 
32'd4164: dataIn2 = 32'd0; 
32'd4165: dataIn2 = 32'd0; 
32'd4166: dataIn2 = 32'd1; 
32'd4167: dataIn2 = 32'd0; 
32'd4168: dataIn2 = 32'd1; 
32'd4169: dataIn2 = 32'd0; 
32'd4170: dataIn2 = 32'd0; 
32'd4171: dataIn2 = 32'd0; 
32'd4172: dataIn2 = 32'd0; 
32'd4173: dataIn2 = 32'd0; 
32'd4174: dataIn2 = 32'd1; 
32'd4175: dataIn2 = 32'd1; 
32'd4176: dataIn2 = 32'd0; 
32'd4177: dataIn2 = 32'd1; 
32'd4178: dataIn2 = 32'd1; 
32'd4179: dataIn2 = 32'd0; 
32'd4180: dataIn2 = 32'd1; 
32'd4181: dataIn2 = 32'd0; 
32'd4182: dataIn2 = 32'd0; 
32'd4183: dataIn2 = 32'd0; 
32'd4184: dataIn2 = 32'd0; 
32'd4185: dataIn2 = 32'd1; 
32'd4186: dataIn2 = 32'd1; 
32'd4187: dataIn2 = 32'd1; 
32'd4188: dataIn2 = 32'd1; 
32'd4189: dataIn2 = 32'd1; 
32'd4190: dataIn2 = 32'd0; 
32'd4191: dataIn2 = 32'd0; 
32'd4192: dataIn2 = 32'd0; 
32'd4193: dataIn2 = 32'd0; 
32'd4194: dataIn2 = 32'd0; 
32'd4195: dataIn2 = 32'd1; 
32'd4196: dataIn2 = 32'd0; 
32'd4197: dataIn2 = 32'd0; 
32'd4198: dataIn2 = 32'd1; 
32'd4199: dataIn2 = 32'd0; 
32'd4200: dataIn2 = 32'd0; 
32'd4201: dataIn2 = 32'd0; 
32'd4202: dataIn2 = 32'd1; 
32'd4203: dataIn2 = 32'd0; 
32'd4204: dataIn2 = 32'd0; 
32'd4205: dataIn2 = 32'd1; 
32'd4206: dataIn2 = 32'd1; 
32'd4207: dataIn2 = 32'd0; 
32'd4208: dataIn2 = 32'd1; 
32'd4209: dataIn2 = 32'd1; 
32'd4210: dataIn2 = 32'd0; 
32'd4211: dataIn2 = 32'd1; 
32'd4212: dataIn2 = 32'd0; 
32'd4213: dataIn2 = 32'd1; 
32'd4214: dataIn2 = 32'd0; 
32'd4215: dataIn2 = 32'd1; 
32'd4216: dataIn2 = 32'd0; 
32'd4217: dataIn2 = 32'd0; 
32'd4218: dataIn2 = 32'd1; 
32'd4219: dataIn2 = 32'd1; 
32'd4220: dataIn2 = 32'd1; 
32'd4221: dataIn2 = 32'd1; 
32'd4222: dataIn2 = 32'd1; 
32'd4223: dataIn2 = 32'd1; 
32'd4224: dataIn2 = 32'd0; 
32'd4225: dataIn2 = 32'd0; 
32'd4226: dataIn2 = 32'd1; 
32'd4227: dataIn2 = 32'd1; 
32'd4228: dataIn2 = 32'd0; 
32'd4229: dataIn2 = 32'd0; 
32'd4230: dataIn2 = 32'd1; 
32'd4231: dataIn2 = 32'd1; 
32'd4232: dataIn2 = 32'd0; 
32'd4233: dataIn2 = 32'd1; 
32'd4234: dataIn2 = 32'd0; 
32'd4235: dataIn2 = 32'd0; 
32'd4236: dataIn2 = 32'd0; 
32'd4237: dataIn2 = 32'd1; 
32'd4238: dataIn2 = 32'd1; 
32'd4239: dataIn2 = 32'd0; 
32'd4240: dataIn2 = 32'd0; 
32'd4241: dataIn2 = 32'd1; 
32'd4242: dataIn2 = 32'd0; 
32'd4243: dataIn2 = 32'd1; 
32'd4244: dataIn2 = 32'd1; 
32'd4245: dataIn2 = 32'd1; 
32'd4246: dataIn2 = 32'd0; 
32'd4247: dataIn2 = 32'd1; 
32'd4248: dataIn2 = 32'd1; 
32'd4249: dataIn2 = 32'd0; 
32'd4250: dataIn2 = 32'd1; 
32'd4251: dataIn2 = 32'd1; 
32'd4252: dataIn2 = 32'd1; 
32'd4253: dataIn2 = 32'd0; 
32'd4254: dataIn2 = 32'd0; 
32'd4255: dataIn2 = 32'd0; 
32'd4256: dataIn2 = 32'd0; 
32'd4257: dataIn2 = 32'd1; 
32'd4258: dataIn2 = 32'd0; 
32'd4259: dataIn2 = 32'd1; 
32'd4260: dataIn2 = 32'd0; 
32'd4261: dataIn2 = 32'd1; 
32'd4262: dataIn2 = 32'd0; 
32'd4263: dataIn2 = 32'd0; 
32'd4264: dataIn2 = 32'd0; 
32'd4265: dataIn2 = 32'd0; 
32'd4266: dataIn2 = 32'd1; 
32'd4267: dataIn2 = 32'd1; 
32'd4268: dataIn2 = 32'd1; 
32'd4269: dataIn2 = 32'd1; 
32'd4270: dataIn2 = 32'd0; 
32'd4271: dataIn2 = 32'd0; 
32'd4272: dataIn2 = 32'd1; 
32'd4273: dataIn2 = 32'd1; 
32'd4274: dataIn2 = 32'd1; 
32'd4275: dataIn2 = 32'd1; 
32'd4276: dataIn2 = 32'd0; 
32'd4277: dataIn2 = 32'd0; 
32'd4278: dataIn2 = 32'd1; 
32'd4279: dataIn2 = 32'd1; 
32'd4280: dataIn2 = 32'd0; 
32'd4281: dataIn2 = 32'd0; 
32'd4282: dataIn2 = 32'd1; 
32'd4283: dataIn2 = 32'd0; 
32'd4284: dataIn2 = 32'd1; 
32'd4285: dataIn2 = 32'd0; 
32'd4286: dataIn2 = 32'd0; 
32'd4287: dataIn2 = 32'd1; 
32'd4288: dataIn2 = 32'd1; 
32'd4289: dataIn2 = 32'd1; 
32'd4290: dataIn2 = 32'd1; 
32'd4291: dataIn2 = 32'd1; 
32'd4292: dataIn2 = 32'd0; 
32'd4293: dataIn2 = 32'd1; 
32'd4294: dataIn2 = 32'd0; 
32'd4295: dataIn2 = 32'd1; 
32'd4296: dataIn2 = 32'd1; 
32'd4297: dataIn2 = 32'd1; 
32'd4298: dataIn2 = 32'd0; 
32'd4299: dataIn2 = 32'd0; 
32'd4300: dataIn2 = 32'd0; 
32'd4301: dataIn2 = 32'd0; 
32'd4302: dataIn2 = 32'd1; 
32'd4303: dataIn2 = 32'd0; 
32'd4304: dataIn2 = 32'd0; 
32'd4305: dataIn2 = 32'd1; 
32'd4306: dataIn2 = 32'd0; 
32'd4307: dataIn2 = 32'd1; 
32'd4308: dataIn2 = 32'd0; 
32'd4309: dataIn2 = 32'd0; 
32'd4310: dataIn2 = 32'd1; 
32'd4311: dataIn2 = 32'd1; 
32'd4312: dataIn2 = 32'd1; 
32'd4313: dataIn2 = 32'd0; 
32'd4314: dataIn2 = 32'd1; 
32'd4315: dataIn2 = 32'd1; 
32'd4316: dataIn2 = 32'd0; 
32'd4317: dataIn2 = 32'd1; 
32'd4318: dataIn2 = 32'd0; 
32'd4319: dataIn2 = 32'd0; 
32'd4320: dataIn2 = 32'd1; 
32'd4321: dataIn2 = 32'd0; 
32'd4322: dataIn2 = 32'd1; 
32'd4323: dataIn2 = 32'd0; 
32'd4324: dataIn2 = 32'd0; 
32'd4325: dataIn2 = 32'd1; 
32'd4326: dataIn2 = 32'd1; 
32'd4327: dataIn2 = 32'd0; 
32'd4328: dataIn2 = 32'd0; 
32'd4329: dataIn2 = 32'd0; 
32'd4330: dataIn2 = 32'd0; 
32'd4331: dataIn2 = 32'd1; 
32'd4332: dataIn2 = 32'd0; 
32'd4333: dataIn2 = 32'd1; 
32'd4334: dataIn2 = 32'd1; 
32'd4335: dataIn2 = 32'd0; 
32'd4336: dataIn2 = 32'd0; 
32'd4337: dataIn2 = 32'd0; 
32'd4338: dataIn2 = 32'd1; 
32'd4339: dataIn2 = 32'd0; 
32'd4340: dataIn2 = 32'd0; 
32'd4341: dataIn2 = 32'd1; 
32'd4342: dataIn2 = 32'd1; 
32'd4343: dataIn2 = 32'd0; 
32'd4344: dataIn2 = 32'd0; 
32'd4345: dataIn2 = 32'd1; 
32'd4346: dataIn2 = 32'd1; 
32'd4347: dataIn2 = 32'd1; 
32'd4348: dataIn2 = 32'd0; 
32'd4349: dataIn2 = 32'd0; 
32'd4350: dataIn2 = 32'd0; 
32'd4351: dataIn2 = 32'd0; 
32'd4352: dataIn2 = 32'd1; 
32'd4353: dataIn2 = 32'd0; 
32'd4354: dataIn2 = 32'd1; 
32'd4355: dataIn2 = 32'd1; 
32'd4356: dataIn2 = 32'd1; 
32'd4357: dataIn2 = 32'd0; 
32'd4358: dataIn2 = 32'd1; 
32'd4359: dataIn2 = 32'd1; 
32'd4360: dataIn2 = 32'd1; 
32'd4361: dataIn2 = 32'd1; 
32'd4362: dataIn2 = 32'd0; 
32'd4363: dataIn2 = 32'd1; 
32'd4364: dataIn2 = 32'd0; 
32'd4365: dataIn2 = 32'd0; 
32'd4366: dataIn2 = 32'd1; 
32'd4367: dataIn2 = 32'd1; 
32'd4368: dataIn2 = 32'd0; 
32'd4369: dataIn2 = 32'd1; 
32'd4370: dataIn2 = 32'd1; 
32'd4371: dataIn2 = 32'd1; 
32'd4372: dataIn2 = 32'd0; 
32'd4373: dataIn2 = 32'd0; 
32'd4374: dataIn2 = 32'd1; 
32'd4375: dataIn2 = 32'd0; 
32'd4376: dataIn2 = 32'd1; 
32'd4377: dataIn2 = 32'd0; 
32'd4378: dataIn2 = 32'd1; 
32'd4379: dataIn2 = 32'd0; 
32'd4380: dataIn2 = 32'd1; 
32'd4381: dataIn2 = 32'd0; 
32'd4382: dataIn2 = 32'd1; 
32'd4383: dataIn2 = 32'd0; 
32'd4384: dataIn2 = 32'd0; 
32'd4385: dataIn2 = 32'd1; 
32'd4386: dataIn2 = 32'd0; 
32'd4387: dataIn2 = 32'd1; 
32'd4388: dataIn2 = 32'd1; 
32'd4389: dataIn2 = 32'd1; 
32'd4390: dataIn2 = 32'd1; 
32'd4391: dataIn2 = 32'd0; 
32'd4392: dataIn2 = 32'd0; 
32'd4393: dataIn2 = 32'd1; 
32'd4394: dataIn2 = 32'd0; 
32'd4395: dataIn2 = 32'd0; 
32'd4396: dataIn2 = 32'd1; 
32'd4397: dataIn2 = 32'd0; 
32'd4398: dataIn2 = 32'd1; 
32'd4399: dataIn2 = 32'd1; 
32'd4400: dataIn2 = 32'd0; 
32'd4401: dataIn2 = 32'd1; 
32'd4402: dataIn2 = 32'd1; 
32'd4403: dataIn2 = 32'd1; 
32'd4404: dataIn2 = 32'd0; 
32'd4405: dataIn2 = 32'd0; 
32'd4406: dataIn2 = 32'd0; 
32'd4407: dataIn2 = 32'd1; 
32'd4408: dataIn2 = 32'd0; 
32'd4409: dataIn2 = 32'd0; 
32'd4410: dataIn2 = 32'd1; 
32'd4411: dataIn2 = 32'd0; 
32'd4412: dataIn2 = 32'd1; 
32'd4413: dataIn2 = 32'd1; 
32'd4414: dataIn2 = 32'd1; 
32'd4415: dataIn2 = 32'd0; 
32'd4416: dataIn2 = 32'd0; 
32'd4417: dataIn2 = 32'd1; 
32'd4418: dataIn2 = 32'd0; 
32'd4419: dataIn2 = 32'd0; 
32'd4420: dataIn2 = 32'd1; 
32'd4421: dataIn2 = 32'd1; 
32'd4422: dataIn2 = 32'd0; 
32'd4423: dataIn2 = 32'd0; 
32'd4424: dataIn2 = 32'd1; 
32'd4425: dataIn2 = 32'd0; 
32'd4426: dataIn2 = 32'd1; 
32'd4427: dataIn2 = 32'd0; 
32'd4428: dataIn2 = 32'd1; 
32'd4429: dataIn2 = 32'd0; 
32'd4430: dataIn2 = 32'd1; 
32'd4431: dataIn2 = 32'd1; 
32'd4432: dataIn2 = 32'd1; 
32'd4433: dataIn2 = 32'd1; 
32'd4434: dataIn2 = 32'd1; 
32'd4435: dataIn2 = 32'd0; 
32'd4436: dataIn2 = 32'd0; 
32'd4437: dataIn2 = 32'd1; 
32'd4438: dataIn2 = 32'd0; 
32'd4439: dataIn2 = 32'd1; 
32'd4440: dataIn2 = 32'd1; 
32'd4441: dataIn2 = 32'd1; 
32'd4442: dataIn2 = 32'd1; 
32'd4443: dataIn2 = 32'd0; 
32'd4444: dataIn2 = 32'd0; 
32'd4445: dataIn2 = 32'd1; 
32'd4446: dataIn2 = 32'd1; 
32'd4447: dataIn2 = 32'd0; 
32'd4448: dataIn2 = 32'd0; 
32'd4449: dataIn2 = 32'd1; 
32'd4450: dataIn2 = 32'd1; 
32'd4451: dataIn2 = 32'd0; 
32'd4452: dataIn2 = 32'd1; 
32'd4453: dataIn2 = 32'd1; 
32'd4454: dataIn2 = 32'd0; 
32'd4455: dataIn2 = 32'd1; 
32'd4456: dataIn2 = 32'd1; 
32'd4457: dataIn2 = 32'd1; 
32'd4458: dataIn2 = 32'd1; 
32'd4459: dataIn2 = 32'd0; 
32'd4460: dataIn2 = 32'd1; 
32'd4461: dataIn2 = 32'd0; 
32'd4462: dataIn2 = 32'd0; 
32'd4463: dataIn2 = 32'd1; 
32'd4464: dataIn2 = 32'd1; 
32'd4465: dataIn2 = 32'd1; 
32'd4466: dataIn2 = 32'd0; 
32'd4467: dataIn2 = 32'd1; 
32'd4468: dataIn2 = 32'd1; 
32'd4469: dataIn2 = 32'd1; 
32'd4470: dataIn2 = 32'd0; 
32'd4471: dataIn2 = 32'd1; 
32'd4472: dataIn2 = 32'd1; 
32'd4473: dataIn2 = 32'd0; 
32'd4474: dataIn2 = 32'd1; 
32'd4475: dataIn2 = 32'd1; 
32'd4476: dataIn2 = 32'd0; 
32'd4477: dataIn2 = 32'd0; 
32'd4478: dataIn2 = 32'd1; 
32'd4479: dataIn2 = 32'd0; 
32'd4480: dataIn2 = 32'd1; 
32'd4481: dataIn2 = 32'd0; 
32'd4482: dataIn2 = 32'd1; 
32'd4483: dataIn2 = 32'd0; 
32'd4484: dataIn2 = 32'd0; 
32'd4485: dataIn2 = 32'd1; 
32'd4486: dataIn2 = 32'd0; 
32'd4487: dataIn2 = 32'd1; 
32'd4488: dataIn2 = 32'd1; 
32'd4489: dataIn2 = 32'd1; 
32'd4490: dataIn2 = 32'd1; 
32'd4491: dataIn2 = 32'd1; 
32'd4492: dataIn2 = 32'd1; 
32'd4493: dataIn2 = 32'd1; 
32'd4494: dataIn2 = 32'd0; 
32'd4495: dataIn2 = 32'd0; 
32'd4496: dataIn2 = 32'd1; 
32'd4497: dataIn2 = 32'd0; 
32'd4498: dataIn2 = 32'd1; 
32'd4499: dataIn2 = 32'd1; 
32'd4500: dataIn2 = 32'd0; 
32'd4501: dataIn2 = 32'd1; 
32'd4502: dataIn2 = 32'd1; 
32'd4503: dataIn2 = 32'd0; 
32'd4504: dataIn2 = 32'd0; 
32'd4505: dataIn2 = 32'd1; 
32'd4506: dataIn2 = 32'd1; 
32'd4507: dataIn2 = 32'd0; 
32'd4508: dataIn2 = 32'd1; 
32'd4509: dataIn2 = 32'd0; 
32'd4510: dataIn2 = 32'd1; 
32'd4511: dataIn2 = 32'd1; 
32'd4512: dataIn2 = 32'd1; 
32'd4513: dataIn2 = 32'd0; 
32'd4514: dataIn2 = 32'd0; 
32'd4515: dataIn2 = 32'd1; 
32'd4516: dataIn2 = 32'd0; 
32'd4517: dataIn2 = 32'd1; 
32'd4518: dataIn2 = 32'd0; 
32'd4519: dataIn2 = 32'd0; 
32'd4520: dataIn2 = 32'd1; 
32'd4521: dataIn2 = 32'd0; 
32'd4522: dataIn2 = 32'd1; 
32'd4523: dataIn2 = 32'd0; 
32'd4524: dataIn2 = 32'd0; 
32'd4525: dataIn2 = 32'd1; 
32'd4526: dataIn2 = 32'd1; 
32'd4527: dataIn2 = 32'd0; 
32'd4528: dataIn2 = 32'd0; 
32'd4529: dataIn2 = 32'd0; 
32'd4530: dataIn2 = 32'd0; 
32'd4531: dataIn2 = 32'd0; 
32'd4532: dataIn2 = 32'd1; 
32'd4533: dataIn2 = 32'd0; 
32'd4534: dataIn2 = 32'd0; 
32'd4535: dataIn2 = 32'd1; 
32'd4536: dataIn2 = 32'd1; 
32'd4537: dataIn2 = 32'd1; 
32'd4538: dataIn2 = 32'd0; 
32'd4539: dataIn2 = 32'd0; 
32'd4540: dataIn2 = 32'd0; 
32'd4541: dataIn2 = 32'd1; 
32'd4542: dataIn2 = 32'd0; 
32'd4543: dataIn2 = 32'd0; 
32'd4544: dataIn2 = 32'd0; 
32'd4545: dataIn2 = 32'd1; 
32'd4546: dataIn2 = 32'd0; 
32'd4547: dataIn2 = 32'd1; 
32'd4548: dataIn2 = 32'd0; 
32'd4549: dataIn2 = 32'd0; 
32'd4550: dataIn2 = 32'd1; 
32'd4551: dataIn2 = 32'd1; 
32'd4552: dataIn2 = 32'd1; 
32'd4553: dataIn2 = 32'd0; 
32'd4554: dataIn2 = 32'd0; 
32'd4555: dataIn2 = 32'd1; 
32'd4556: dataIn2 = 32'd1; 
32'd4557: dataIn2 = 32'd0; 
32'd4558: dataIn2 = 32'd0; 
32'd4559: dataIn2 = 32'd0; 
32'd4560: dataIn2 = 32'd0; 
32'd4561: dataIn2 = 32'd0; 
32'd4562: dataIn2 = 32'd0; 
32'd4563: dataIn2 = 32'd0; 
32'd4564: dataIn2 = 32'd0; 
32'd4565: dataIn2 = 32'd0; 
32'd4566: dataIn2 = 32'd0; 
32'd4567: dataIn2 = 32'd1; 
32'd4568: dataIn2 = 32'd1; 
32'd4569: dataIn2 = 32'd0; 
32'd4570: dataIn2 = 32'd1; 
32'd4571: dataIn2 = 32'd0; 
32'd4572: dataIn2 = 32'd1; 
32'd4573: dataIn2 = 32'd1; 
32'd4574: dataIn2 = 32'd1; 
32'd4575: dataIn2 = 32'd1; 
32'd4576: dataIn2 = 32'd0; 
32'd4577: dataIn2 = 32'd1; 
32'd4578: dataIn2 = 32'd0; 
32'd4579: dataIn2 = 32'd0; 
32'd4580: dataIn2 = 32'd0; 
32'd4581: dataIn2 = 32'd0; 
32'd4582: dataIn2 = 32'd1; 
32'd4583: dataIn2 = 32'd0; 
32'd4584: dataIn2 = 32'd1; 
32'd4585: dataIn2 = 32'd0; 
32'd4586: dataIn2 = 32'd1; 
32'd4587: dataIn2 = 32'd1; 
32'd4588: dataIn2 = 32'd1; 
32'd4589: dataIn2 = 32'd1; 
32'd4590: dataIn2 = 32'd1; 
32'd4591: dataIn2 = 32'd1; 
32'd4592: dataIn2 = 32'd1; 
32'd4593: dataIn2 = 32'd0; 
32'd4594: dataIn2 = 32'd0; 
32'd4595: dataIn2 = 32'd1; 
32'd4596: dataIn2 = 32'd1; 
32'd4597: dataIn2 = 32'd0; 
32'd4598: dataIn2 = 32'd1; 
32'd4599: dataIn2 = 32'd0; 
32'd4600: dataIn2 = 32'd0; 
32'd4601: dataIn2 = 32'd1; 
32'd4602: dataIn2 = 32'd0; 
32'd4603: dataIn2 = 32'd0; 
32'd4604: dataIn2 = 32'd0; 
32'd4605: dataIn2 = 32'd0; 
32'd4606: dataIn2 = 32'd1; 
32'd4607: dataIn2 = 32'd0; 
32'd4608: dataIn2 = 32'd0; 
32'd4609: dataIn2 = 32'd1; 
32'd4610: dataIn2 = 32'd1; 
32'd4611: dataIn2 = 32'd1; 
32'd4612: dataIn2 = 32'd1; 
32'd4613: dataIn2 = 32'd1; 
32'd4614: dataIn2 = 32'd0; 
32'd4615: dataIn2 = 32'd0; 
32'd4616: dataIn2 = 32'd0; 
32'd4617: dataIn2 = 32'd0; 
32'd4618: dataIn2 = 32'd0; 
32'd4619: dataIn2 = 32'd1; 
32'd4620: dataIn2 = 32'd1; 
32'd4621: dataIn2 = 32'd1; 
32'd4622: dataIn2 = 32'd0; 
32'd4623: dataIn2 = 32'd0; 
32'd4624: dataIn2 = 32'd1; 
32'd4625: dataIn2 = 32'd1; 
32'd4626: dataIn2 = 32'd0; 
32'd4627: dataIn2 = 32'd0; 
32'd4628: dataIn2 = 32'd1; 
32'd4629: dataIn2 = 32'd1; 
32'd4630: dataIn2 = 32'd1; 
32'd4631: dataIn2 = 32'd0; 
32'd4632: dataIn2 = 32'd1; 
32'd4633: dataIn2 = 32'd0; 
32'd4634: dataIn2 = 32'd1; 
32'd4635: dataIn2 = 32'd1; 
32'd4636: dataIn2 = 32'd1; 
32'd4637: dataIn2 = 32'd1; 
32'd4638: dataIn2 = 32'd0; 
32'd4639: dataIn2 = 32'd1; 
32'd4640: dataIn2 = 32'd0; 
32'd4641: dataIn2 = 32'd1; 
32'd4642: dataIn2 = 32'd0; 
32'd4643: dataIn2 = 32'd0; 
32'd4644: dataIn2 = 32'd0; 
32'd4645: dataIn2 = 32'd1; 
32'd4646: dataIn2 = 32'd0; 
32'd4647: dataIn2 = 32'd0; 
32'd4648: dataIn2 = 32'd0; 
32'd4649: dataIn2 = 32'd0; 
32'd4650: dataIn2 = 32'd1; 
32'd4651: dataIn2 = 32'd0; 
32'd4652: dataIn2 = 32'd1; 
32'd4653: dataIn2 = 32'd1; 
32'd4654: dataIn2 = 32'd1; 
32'd4655: dataIn2 = 32'd0; 
32'd4656: dataIn2 = 32'd1; 
32'd4657: dataIn2 = 32'd0; 
32'd4658: dataIn2 = 32'd0; 
32'd4659: dataIn2 = 32'd1; 
32'd4660: dataIn2 = 32'd0; 
32'd4661: dataIn2 = 32'd0; 
32'd4662: dataIn2 = 32'd1; 
32'd4663: dataIn2 = 32'd1; 
32'd4664: dataIn2 = 32'd1; 
32'd4665: dataIn2 = 32'd1; 
32'd4666: dataIn2 = 32'd0; 
32'd4667: dataIn2 = 32'd1; 
32'd4668: dataIn2 = 32'd1; 
32'd4669: dataIn2 = 32'd0; 
32'd4670: dataIn2 = 32'd0; 
32'd4671: dataIn2 = 32'd0; 
32'd4672: dataIn2 = 32'd0; 
32'd4673: dataIn2 = 32'd0; 
32'd4674: dataIn2 = 32'd1; 
32'd4675: dataIn2 = 32'd0; 
32'd4676: dataIn2 = 32'd1; 
32'd4677: dataIn2 = 32'd0; 
32'd4678: dataIn2 = 32'd0; 
32'd4679: dataIn2 = 32'd1; 
32'd4680: dataIn2 = 32'd1; 
32'd4681: dataIn2 = 32'd0; 
32'd4682: dataIn2 = 32'd1; 
32'd4683: dataIn2 = 32'd0; 
32'd4684: dataIn2 = 32'd0; 
32'd4685: dataIn2 = 32'd1; 
32'd4686: dataIn2 = 32'd0; 
32'd4687: dataIn2 = 32'd1; 
32'd4688: dataIn2 = 32'd0; 
32'd4689: dataIn2 = 32'd0; 
32'd4690: dataIn2 = 32'd1; 
32'd4691: dataIn2 = 32'd1; 
32'd4692: dataIn2 = 32'd1; 
32'd4693: dataIn2 = 32'd0; 
32'd4694: dataIn2 = 32'd0; 
32'd4695: dataIn2 = 32'd1; 
32'd4696: dataIn2 = 32'd1; 
32'd4697: dataIn2 = 32'd1; 
32'd4698: dataIn2 = 32'd1; 
32'd4699: dataIn2 = 32'd1; 
32'd4700: dataIn2 = 32'd0; 
32'd4701: dataIn2 = 32'd1; 
32'd4702: dataIn2 = 32'd0; 
32'd4703: dataIn2 = 32'd1; 
32'd4704: dataIn2 = 32'd1; 
32'd4705: dataIn2 = 32'd1; 
32'd4706: dataIn2 = 32'd1; 
32'd4707: dataIn2 = 32'd0; 
32'd4708: dataIn2 = 32'd0; 
32'd4709: dataIn2 = 32'd1; 
32'd4710: dataIn2 = 32'd1; 
32'd4711: dataIn2 = 32'd1; 
32'd4712: dataIn2 = 32'd1; 
32'd4713: dataIn2 = 32'd1; 
32'd4714: dataIn2 = 32'd1; 
32'd4715: dataIn2 = 32'd1; 
32'd4716: dataIn2 = 32'd0; 
32'd4717: dataIn2 = 32'd1; 
32'd4718: dataIn2 = 32'd1; 
32'd4719: dataIn2 = 32'd0; 
32'd4720: dataIn2 = 32'd1; 
32'd4721: dataIn2 = 32'd1; 
32'd4722: dataIn2 = 32'd0; 
32'd4723: dataIn2 = 32'd1; 
32'd4724: dataIn2 = 32'd1; 
32'd4725: dataIn2 = 32'd1; 
32'd4726: dataIn2 = 32'd1; 
32'd4727: dataIn2 = 32'd1; 
32'd4728: dataIn2 = 32'd0; 
32'd4729: dataIn2 = 32'd0; 
32'd4730: dataIn2 = 32'd1; 
32'd4731: dataIn2 = 32'd0; 
32'd4732: dataIn2 = 32'd0; 
32'd4733: dataIn2 = 32'd1; 
32'd4734: dataIn2 = 32'd0; 
32'd4735: dataIn2 = 32'd1; 
32'd4736: dataIn2 = 32'd1; 
32'd4737: dataIn2 = 32'd0; 
32'd4738: dataIn2 = 32'd1; 
32'd4739: dataIn2 = 32'd0; 
32'd4740: dataIn2 = 32'd1; 
32'd4741: dataIn2 = 32'd1; 
32'd4742: dataIn2 = 32'd1; 
32'd4743: dataIn2 = 32'd1; 
32'd4744: dataIn2 = 32'd1; 
32'd4745: dataIn2 = 32'd0; 
32'd4746: dataIn2 = 32'd0; 
32'd4747: dataIn2 = 32'd0; 
32'd4748: dataIn2 = 32'd1; 
32'd4749: dataIn2 = 32'd0; 
32'd4750: dataIn2 = 32'd1; 
32'd4751: dataIn2 = 32'd0; 
32'd4752: dataIn2 = 32'd1; 
32'd4753: dataIn2 = 32'd0; 
32'd4754: dataIn2 = 32'd0; 
32'd4755: dataIn2 = 32'd1; 
32'd4756: dataIn2 = 32'd1; 
32'd4757: dataIn2 = 32'd0; 
32'd4758: dataIn2 = 32'd0; 
32'd4759: dataIn2 = 32'd1; 
32'd4760: dataIn2 = 32'd0; 
32'd4761: dataIn2 = 32'd1; 
32'd4762: dataIn2 = 32'd0; 
32'd4763: dataIn2 = 32'd1; 
32'd4764: dataIn2 = 32'd1; 
32'd4765: dataIn2 = 32'd0; 
32'd4766: dataIn2 = 32'd0; 
32'd4767: dataIn2 = 32'd0; 
32'd4768: dataIn2 = 32'd1; 
32'd4769: dataIn2 = 32'd0; 
32'd4770: dataIn2 = 32'd0; 
32'd4771: dataIn2 = 32'd1; 
32'd4772: dataIn2 = 32'd0; 
32'd4773: dataIn2 = 32'd0; 
32'd4774: dataIn2 = 32'd0; 
32'd4775: dataIn2 = 32'd1; 
32'd4776: dataIn2 = 32'd1; 
32'd4777: dataIn2 = 32'd0; 
32'd4778: dataIn2 = 32'd1; 
32'd4779: dataIn2 = 32'd1; 
32'd4780: dataIn2 = 32'd0; 
32'd4781: dataIn2 = 32'd1; 
32'd4782: dataIn2 = 32'd1; 
32'd4783: dataIn2 = 32'd0; 
32'd4784: dataIn2 = 32'd1; 
32'd4785: dataIn2 = 32'd1; 
32'd4786: dataIn2 = 32'd1; 
32'd4787: dataIn2 = 32'd0; 
32'd4788: dataIn2 = 32'd1; 
32'd4789: dataIn2 = 32'd1; 
32'd4790: dataIn2 = 32'd1; 
32'd4791: dataIn2 = 32'd0; 
32'd4792: dataIn2 = 32'd1; 
32'd4793: dataIn2 = 32'd0; 
32'd4794: dataIn2 = 32'd0; 
32'd4795: dataIn2 = 32'd0; 
32'd4796: dataIn2 = 32'd0; 
32'd4797: dataIn2 = 32'd1; 
32'd4798: dataIn2 = 32'd1; 
32'd4799: dataIn2 = 32'd1; 
32'd4800: dataIn2 = 32'd0; 
32'd4801: dataIn2 = 32'd0; 
32'd4802: dataIn2 = 32'd1; 
32'd4803: dataIn2 = 32'd0; 
32'd4804: dataIn2 = 32'd1; 
32'd4805: dataIn2 = 32'd1; 
32'd4806: dataIn2 = 32'd0; 
32'd4807: dataIn2 = 32'd0; 
32'd4808: dataIn2 = 32'd0; 
32'd4809: dataIn2 = 32'd1; 
32'd4810: dataIn2 = 32'd1; 
32'd4811: dataIn2 = 32'd0; 
32'd4812: dataIn2 = 32'd1; 
32'd4813: dataIn2 = 32'd0; 
32'd4814: dataIn2 = 32'd0; 
32'd4815: dataIn2 = 32'd1; 
32'd4816: dataIn2 = 32'd1; 
32'd4817: dataIn2 = 32'd0; 
32'd4818: dataIn2 = 32'd1; 
32'd4819: dataIn2 = 32'd0; 
32'd4820: dataIn2 = 32'd0; 
32'd4821: dataIn2 = 32'd1; 
32'd4822: dataIn2 = 32'd0; 
32'd4823: dataIn2 = 32'd0; 
32'd4824: dataIn2 = 32'd1; 
32'd4825: dataIn2 = 32'd1; 
32'd4826: dataIn2 = 32'd0; 
32'd4827: dataIn2 = 32'd0; 
32'd4828: dataIn2 = 32'd1; 
32'd4829: dataIn2 = 32'd1; 
32'd4830: dataIn2 = 32'd1; 
32'd4831: dataIn2 = 32'd0; 
32'd4832: dataIn2 = 32'd1; 
32'd4833: dataIn2 = 32'd0; 
32'd4834: dataIn2 = 32'd0; 
32'd4835: dataIn2 = 32'd0; 
32'd4836: dataIn2 = 32'd0; 
32'd4837: dataIn2 = 32'd1; 
32'd4838: dataIn2 = 32'd0; 
32'd4839: dataIn2 = 32'd0; 
32'd4840: dataIn2 = 32'd0; 
32'd4841: dataIn2 = 32'd0; 
32'd4842: dataIn2 = 32'd1; 
32'd4843: dataIn2 = 32'd1; 
32'd4844: dataIn2 = 32'd0; 
32'd4845: dataIn2 = 32'd1; 
32'd4846: dataIn2 = 32'd1; 
32'd4847: dataIn2 = 32'd1; 
32'd4848: dataIn2 = 32'd1; 
32'd4849: dataIn2 = 32'd0; 
32'd4850: dataIn2 = 32'd0; 
32'd4851: dataIn2 = 32'd0; 
32'd4852: dataIn2 = 32'd1; 
32'd4853: dataIn2 = 32'd1; 
32'd4854: dataIn2 = 32'd0; 
32'd4855: dataIn2 = 32'd1; 
32'd4856: dataIn2 = 32'd1; 
32'd4857: dataIn2 = 32'd0; 
32'd4858: dataIn2 = 32'd0; 
32'd4859: dataIn2 = 32'd0; 
32'd4860: dataIn2 = 32'd1; 
32'd4861: dataIn2 = 32'd1; 
32'd4862: dataIn2 = 32'd1; 
32'd4863: dataIn2 = 32'd1; 
32'd4864: dataIn2 = 32'd0; 
32'd4865: dataIn2 = 32'd1; 
32'd4866: dataIn2 = 32'd0; 
32'd4867: dataIn2 = 32'd0; 
32'd4868: dataIn2 = 32'd0; 
32'd4869: dataIn2 = 32'd0; 
32'd4870: dataIn2 = 32'd1; 
32'd4871: dataIn2 = 32'd0; 
32'd4872: dataIn2 = 32'd1; 
32'd4873: dataIn2 = 32'd1; 
32'd4874: dataIn2 = 32'd0; 
32'd4875: dataIn2 = 32'd1; 
32'd4876: dataIn2 = 32'd0; 
32'd4877: dataIn2 = 32'd1; 
32'd4878: dataIn2 = 32'd0; 
32'd4879: dataIn2 = 32'd0; 
32'd4880: dataIn2 = 32'd0; 
32'd4881: dataIn2 = 32'd1; 
32'd4882: dataIn2 = 32'd1; 
32'd4883: dataIn2 = 32'd1; 
32'd4884: dataIn2 = 32'd1; 
32'd4885: dataIn2 = 32'd0; 
32'd4886: dataIn2 = 32'd1; 
32'd4887: dataIn2 = 32'd0; 
32'd4888: dataIn2 = 32'd0; 
32'd4889: dataIn2 = 32'd0; 
32'd4890: dataIn2 = 32'd1; 
32'd4891: dataIn2 = 32'd0; 
32'd4892: dataIn2 = 32'd1; 
32'd4893: dataIn2 = 32'd1; 
32'd4894: dataIn2 = 32'd0; 
32'd4895: dataIn2 = 32'd0; 
32'd4896: dataIn2 = 32'd0; 
32'd4897: dataIn2 = 32'd0; 
32'd4898: dataIn2 = 32'd1; 
32'd4899: dataIn2 = 32'd1; 
32'd4900: dataIn2 = 32'd1; 
32'd4901: dataIn2 = 32'd1; 
32'd4902: dataIn2 = 32'd1; 
32'd4903: dataIn2 = 32'd1; 
32'd4904: dataIn2 = 32'd0; 
32'd4905: dataIn2 = 32'd1; 
32'd4906: dataIn2 = 32'd0; 
32'd4907: dataIn2 = 32'd0; 
32'd4908: dataIn2 = 32'd0; 
32'd4909: dataIn2 = 32'd1; 
32'd4910: dataIn2 = 32'd1; 
32'd4911: dataIn2 = 32'd0; 
32'd4912: dataIn2 = 32'd0; 
32'd4913: dataIn2 = 32'd0; 
32'd4914: dataIn2 = 32'd1; 
32'd4915: dataIn2 = 32'd0; 
32'd4916: dataIn2 = 32'd1; 
32'd4917: dataIn2 = 32'd0; 
32'd4918: dataIn2 = 32'd0; 
32'd4919: dataIn2 = 32'd0; 
32'd4920: dataIn2 = 32'd1; 
32'd4921: dataIn2 = 32'd0; 
32'd4922: dataIn2 = 32'd0; 
32'd4923: dataIn2 = 32'd0; 
32'd4924: dataIn2 = 32'd1; 
32'd4925: dataIn2 = 32'd0; 
32'd4926: dataIn2 = 32'd0; 
32'd4927: dataIn2 = 32'd1; 
32'd4928: dataIn2 = 32'd0; 
32'd4929: dataIn2 = 32'd0; 
32'd4930: dataIn2 = 32'd0; 
32'd4931: dataIn2 = 32'd1; 
32'd4932: dataIn2 = 32'd1; 
32'd4933: dataIn2 = 32'd0; 
32'd4934: dataIn2 = 32'd0; 
32'd4935: dataIn2 = 32'd0; 
32'd4936: dataIn2 = 32'd0; 
32'd4937: dataIn2 = 32'd1; 
32'd4938: dataIn2 = 32'd1; 
32'd4939: dataIn2 = 32'd1; 
32'd4940: dataIn2 = 32'd0; 
32'd4941: dataIn2 = 32'd1; 
32'd4942: dataIn2 = 32'd0; 
32'd4943: dataIn2 = 32'd0; 
32'd4944: dataIn2 = 32'd1; 
32'd4945: dataIn2 = 32'd0; 
32'd4946: dataIn2 = 32'd0; 
32'd4947: dataIn2 = 32'd0; 
32'd4948: dataIn2 = 32'd0; 
32'd4949: dataIn2 = 32'd1; 
32'd4950: dataIn2 = 32'd1; 
32'd4951: dataIn2 = 32'd1; 
32'd4952: dataIn2 = 32'd0; 
32'd4953: dataIn2 = 32'd1; 
32'd4954: dataIn2 = 32'd0; 
32'd4955: dataIn2 = 32'd0; 
32'd4956: dataIn2 = 32'd1; 
32'd4957: dataIn2 = 32'd1; 
32'd4958: dataIn2 = 32'd0; 
32'd4959: dataIn2 = 32'd1; 
32'd4960: dataIn2 = 32'd1; 
32'd4961: dataIn2 = 32'd0; 
32'd4962: dataIn2 = 32'd0; 
32'd4963: dataIn2 = 32'd1; 
32'd4964: dataIn2 = 32'd0; 
32'd4965: dataIn2 = 32'd0; 
32'd4966: dataIn2 = 32'd0; 
32'd4967: dataIn2 = 32'd0; 
32'd4968: dataIn2 = 32'd1; 
32'd4969: dataIn2 = 32'd0; 
32'd4970: dataIn2 = 32'd0; 
32'd4971: dataIn2 = 32'd0; 
32'd4972: dataIn2 = 32'd1; 
32'd4973: dataIn2 = 32'd0; 
32'd4974: dataIn2 = 32'd1; 
32'd4975: dataIn2 = 32'd1; 
32'd4976: dataIn2 = 32'd0; 
32'd4977: dataIn2 = 32'd1; 
32'd4978: dataIn2 = 32'd0; 
32'd4979: dataIn2 = 32'd1; 
32'd4980: dataIn2 = 32'd1; 
32'd4981: dataIn2 = 32'd0; 
32'd4982: dataIn2 = 32'd1; 
32'd4983: dataIn2 = 32'd0; 
32'd4984: dataIn2 = 32'd0; 
32'd4985: dataIn2 = 32'd0; 
32'd4986: dataIn2 = 32'd0; 
32'd4987: dataIn2 = 32'd0; 
32'd4988: dataIn2 = 32'd1; 
32'd4989: dataIn2 = 32'd1; 
32'd4990: dataIn2 = 32'd0; 
32'd4991: dataIn2 = 32'd1; 
32'd4992: dataIn2 = 32'd0; 
32'd4993: dataIn2 = 32'd1; 
32'd4994: dataIn2 = 32'd1; 
32'd4995: dataIn2 = 32'd1; 
32'd4996: dataIn2 = 32'd0; 
32'd4997: dataIn2 = 32'd1; 
32'd4998: dataIn2 = 32'd0; 
32'd4999: dataIn2 = 32'd1; 
32'd5000: dataIn2 = 32'd0; 
32'd5001: dataIn2 = 32'd0; 
32'd5002: dataIn2 = 32'd0; 
32'd5003: dataIn2 = 32'd0; 
32'd5004: dataIn2 = 32'd1; 
32'd5005: dataIn2 = 32'd0; 
32'd5006: dataIn2 = 32'd1; 
32'd5007: dataIn2 = 32'd0; 
32'd5008: dataIn2 = 32'd0; 
32'd5009: dataIn2 = 32'd0; 
32'd5010: dataIn2 = 32'd1; 
32'd5011: dataIn2 = 32'd1; 
32'd5012: dataIn2 = 32'd0; 
32'd5013: dataIn2 = 32'd0; 
32'd5014: dataIn2 = 32'd0; 
32'd5015: dataIn2 = 32'd0; 
32'd5016: dataIn2 = 32'd1; 
32'd5017: dataIn2 = 32'd0; 
32'd5018: dataIn2 = 32'd1; 
32'd5019: dataIn2 = 32'd0; 
32'd5020: dataIn2 = 32'd0; 
32'd5021: dataIn2 = 32'd1; 
32'd5022: dataIn2 = 32'd1; 
32'd5023: dataIn2 = 32'd0; 
32'd5024: dataIn2 = 32'd1; 
32'd5025: dataIn2 = 32'd1; 
32'd5026: dataIn2 = 32'd1; 
32'd5027: dataIn2 = 32'd1; 
32'd5028: dataIn2 = 32'd1; 
32'd5029: dataIn2 = 32'd0; 
32'd5030: dataIn2 = 32'd1; 
32'd5031: dataIn2 = 32'd1; 
32'd5032: dataIn2 = 32'd0; 
32'd5033: dataIn2 = 32'd1; 
32'd5034: dataIn2 = 32'd0; 
32'd5035: dataIn2 = 32'd1; 
32'd5036: dataIn2 = 32'd1; 
32'd5037: dataIn2 = 32'd0; 
32'd5038: dataIn2 = 32'd1; 
32'd5039: dataIn2 = 32'd1; 
32'd5040: dataIn2 = 32'd0; 
32'd5041: dataIn2 = 32'd0; 
32'd5042: dataIn2 = 32'd0; 
32'd5043: dataIn2 = 32'd1; 
32'd5044: dataIn2 = 32'd0; 
32'd5045: dataIn2 = 32'd0; 
32'd5046: dataIn2 = 32'd0; 
32'd5047: dataIn2 = 32'd0; 
32'd5048: dataIn2 = 32'd0; 
32'd5049: dataIn2 = 32'd0; 
32'd5050: dataIn2 = 32'd1; 
32'd5051: dataIn2 = 32'd1; 
32'd5052: dataIn2 = 32'd1; 
32'd5053: dataIn2 = 32'd0; 
32'd5054: dataIn2 = 32'd1; 
32'd5055: dataIn2 = 32'd1; 
32'd5056: dataIn2 = 32'd0; 
32'd5057: dataIn2 = 32'd1; 
32'd5058: dataIn2 = 32'd1; 
32'd5059: dataIn2 = 32'd0; 
32'd5060: dataIn2 = 32'd0; 
32'd5061: dataIn2 = 32'd0; 
32'd5062: dataIn2 = 32'd1; 
32'd5063: dataIn2 = 32'd0; 
32'd5064: dataIn2 = 32'd0; 
32'd5065: dataIn2 = 32'd1; 
32'd5066: dataIn2 = 32'd1; 
32'd5067: dataIn2 = 32'd0; 
32'd5068: dataIn2 = 32'd0; 
32'd5069: dataIn2 = 32'd0; 
32'd5070: dataIn2 = 32'd1; 
32'd5071: dataIn2 = 32'd1; 
32'd5072: dataIn2 = 32'd0; 
32'd5073: dataIn2 = 32'd1; 
32'd5074: dataIn2 = 32'd0; 
32'd5075: dataIn2 = 32'd0; 
32'd5076: dataIn2 = 32'd1; 
32'd5077: dataIn2 = 32'd0; 
32'd5078: dataIn2 = 32'd1; 
32'd5079: dataIn2 = 32'd1; 
32'd5080: dataIn2 = 32'd0; 
32'd5081: dataIn2 = 32'd0; 
32'd5082: dataIn2 = 32'd0; 
32'd5083: dataIn2 = 32'd0; 
32'd5084: dataIn2 = 32'd1; 
32'd5085: dataIn2 = 32'd0; 
32'd5086: dataIn2 = 32'd1; 
32'd5087: dataIn2 = 32'd1; 
32'd5088: dataIn2 = 32'd1; 
32'd5089: dataIn2 = 32'd1; 
32'd5090: dataIn2 = 32'd1; 
32'd5091: dataIn2 = 32'd1; 
32'd5092: dataIn2 = 32'd1; 
32'd5093: dataIn2 = 32'd1; 
32'd5094: dataIn2 = 32'd1; 
32'd5095: dataIn2 = 32'd0; 
32'd5096: dataIn2 = 32'd0; 
32'd5097: dataIn2 = 32'd0; 
32'd5098: dataIn2 = 32'd0; 
32'd5099: dataIn2 = 32'd0; 
32'd5100: dataIn2 = 32'd1; 
32'd5101: dataIn2 = 32'd1; 
32'd5102: dataIn2 = 32'd1; 
32'd5103: dataIn2 = 32'd0; 
32'd5104: dataIn2 = 32'd0; 
32'd5105: dataIn2 = 32'd1; 
32'd5106: dataIn2 = 32'd0; 
32'd5107: dataIn2 = 32'd0; 
32'd5108: dataIn2 = 32'd0; 
32'd5109: dataIn2 = 32'd1; 
32'd5110: dataIn2 = 32'd0; 
32'd5111: dataIn2 = 32'd0; 
32'd5112: dataIn2 = 32'd0; 
32'd5113: dataIn2 = 32'd0; 
32'd5114: dataIn2 = 32'd0; 
32'd5115: dataIn2 = 32'd0; 
32'd5116: dataIn2 = 32'd1; 
32'd5117: dataIn2 = 32'd0; 
32'd5118: dataIn2 = 32'd1; 
32'd5119: dataIn2 = 32'd0; 
32'd5120: dataIn2 = 32'd0; 
32'd5121: dataIn2 = 32'd1; 
32'd5122: dataIn2 = 32'd0; 
32'd5123: dataIn2 = 32'd0; 
32'd5124: dataIn2 = 32'd0; 
32'd5125: dataIn2 = 32'd0; 
32'd5126: dataIn2 = 32'd0; 
32'd5127: dataIn2 = 32'd0; 
32'd5128: dataIn2 = 32'd0; 
32'd5129: dataIn2 = 32'd1; 
32'd5130: dataIn2 = 32'd1; 
32'd5131: dataIn2 = 32'd1; 
32'd5132: dataIn2 = 32'd1; 
32'd5133: dataIn2 = 32'd1; 
32'd5134: dataIn2 = 32'd0; 
32'd5135: dataIn2 = 32'd0; 
32'd5136: dataIn2 = 32'd0; 
32'd5137: dataIn2 = 32'd0; 
32'd5138: dataIn2 = 32'd1; 
32'd5139: dataIn2 = 32'd0; 
32'd5140: dataIn2 = 32'd1; 
32'd5141: dataIn2 = 32'd1; 
32'd5142: dataIn2 = 32'd0; 
32'd5143: dataIn2 = 32'd0; 
32'd5144: dataIn2 = 32'd0; 
32'd5145: dataIn2 = 32'd1; 
32'd5146: dataIn2 = 32'd1; 
32'd5147: dataIn2 = 32'd0; 
32'd5148: dataIn2 = 32'd1; 
32'd5149: dataIn2 = 32'd1; 
32'd5150: dataIn2 = 32'd0; 
32'd5151: dataIn2 = 32'd0; 
32'd5152: dataIn2 = 32'd0; 
32'd5153: dataIn2 = 32'd1; 
32'd5154: dataIn2 = 32'd1; 
32'd5155: dataIn2 = 32'd1; 
32'd5156: dataIn2 = 32'd1; 
32'd5157: dataIn2 = 32'd0; 
32'd5158: dataIn2 = 32'd1; 
32'd5159: dataIn2 = 32'd1; 
32'd5160: dataIn2 = 32'd1; 
32'd5161: dataIn2 = 32'd1; 
32'd5162: dataIn2 = 32'd0; 
32'd5163: dataIn2 = 32'd0; 
32'd5164: dataIn2 = 32'd1; 
32'd5165: dataIn2 = 32'd1; 
32'd5166: dataIn2 = 32'd0; 
32'd5167: dataIn2 = 32'd1; 
32'd5168: dataIn2 = 32'd0; 
32'd5169: dataIn2 = 32'd1; 
32'd5170: dataIn2 = 32'd0; 
32'd5171: dataIn2 = 32'd1; 
32'd5172: dataIn2 = 32'd0; 
32'd5173: dataIn2 = 32'd0; 
32'd5174: dataIn2 = 32'd1; 
32'd5175: dataIn2 = 32'd0; 
32'd5176: dataIn2 = 32'd1; 
32'd5177: dataIn2 = 32'd1; 
32'd5178: dataIn2 = 32'd1; 
32'd5179: dataIn2 = 32'd0; 
32'd5180: dataIn2 = 32'd0; 
32'd5181: dataIn2 = 32'd0; 
32'd5182: dataIn2 = 32'd1; 
32'd5183: dataIn2 = 32'd0; 
32'd5184: dataIn2 = 32'd1; 
32'd5185: dataIn2 = 32'd0; 
32'd5186: dataIn2 = 32'd1; 
32'd5187: dataIn2 = 32'd0; 
32'd5188: dataIn2 = 32'd1; 
32'd5189: dataIn2 = 32'd0; 
32'd5190: dataIn2 = 32'd0; 
32'd5191: dataIn2 = 32'd0; 
32'd5192: dataIn2 = 32'd1; 
32'd5193: dataIn2 = 32'd1; 
32'd5194: dataIn2 = 32'd1; 
32'd5195: dataIn2 = 32'd1; 
32'd5196: dataIn2 = 32'd0; 
32'd5197: dataIn2 = 32'd1; 
32'd5198: dataIn2 = 32'd0; 
32'd5199: dataIn2 = 32'd1; 
32'd5200: dataIn2 = 32'd0; 
32'd5201: dataIn2 = 32'd1; 
32'd5202: dataIn2 = 32'd0; 
32'd5203: dataIn2 = 32'd1; 
32'd5204: dataIn2 = 32'd0; 
32'd5205: dataIn2 = 32'd1; 
32'd5206: dataIn2 = 32'd1; 
32'd5207: dataIn2 = 32'd0; 
32'd5208: dataIn2 = 32'd0; 
32'd5209: dataIn2 = 32'd1; 
32'd5210: dataIn2 = 32'd0; 
32'd5211: dataIn2 = 32'd0; 
32'd5212: dataIn2 = 32'd1; 
32'd5213: dataIn2 = 32'd0; 
32'd5214: dataIn2 = 32'd1; 
32'd5215: dataIn2 = 32'd0; 
32'd5216: dataIn2 = 32'd0; 
32'd5217: dataIn2 = 32'd0; 
32'd5218: dataIn2 = 32'd0; 
32'd5219: dataIn2 = 32'd1; 
32'd5220: dataIn2 = 32'd1; 
32'd5221: dataIn2 = 32'd1; 
32'd5222: dataIn2 = 32'd1; 
32'd5223: dataIn2 = 32'd0; 
32'd5224: dataIn2 = 32'd0; 
32'd5225: dataIn2 = 32'd0; 
32'd5226: dataIn2 = 32'd1; 
32'd5227: dataIn2 = 32'd1; 
32'd5228: dataIn2 = 32'd1; 
32'd5229: dataIn2 = 32'd1; 
32'd5230: dataIn2 = 32'd0; 
32'd5231: dataIn2 = 32'd1; 
32'd5232: dataIn2 = 32'd1; 
32'd5233: dataIn2 = 32'd0; 
32'd5234: dataIn2 = 32'd1; 
32'd5235: dataIn2 = 32'd1; 
32'd5236: dataIn2 = 32'd0; 
32'd5237: dataIn2 = 32'd0; 
32'd5238: dataIn2 = 32'd1; 
32'd5239: dataIn2 = 32'd1; 
32'd5240: dataIn2 = 32'd0; 
32'd5241: dataIn2 = 32'd1; 
32'd5242: dataIn2 = 32'd0; 
32'd5243: dataIn2 = 32'd0; 
32'd5244: dataIn2 = 32'd0; 
32'd5245: dataIn2 = 32'd0; 
32'd5246: dataIn2 = 32'd1; 
32'd5247: dataIn2 = 32'd1; 
32'd5248: dataIn2 = 32'd1; 
32'd5249: dataIn2 = 32'd0; 
32'd5250: dataIn2 = 32'd1; 
32'd5251: dataIn2 = 32'd0; 
32'd5252: dataIn2 = 32'd0; 
32'd5253: dataIn2 = 32'd0; 
32'd5254: dataIn2 = 32'd0; 
32'd5255: dataIn2 = 32'd0; 
32'd5256: dataIn2 = 32'd1; 
32'd5257: dataIn2 = 32'd0; 
32'd5258: dataIn2 = 32'd1; 
32'd5259: dataIn2 = 32'd1; 
32'd5260: dataIn2 = 32'd1; 
32'd5261: dataIn2 = 32'd1; 
32'd5262: dataIn2 = 32'd0; 
32'd5263: dataIn2 = 32'd1; 
32'd5264: dataIn2 = 32'd0; 
32'd5265: dataIn2 = 32'd0; 
32'd5266: dataIn2 = 32'd0; 
32'd5267: dataIn2 = 32'd0; 
32'd5268: dataIn2 = 32'd0; 
32'd5269: dataIn2 = 32'd1; 
32'd5270: dataIn2 = 32'd1; 
32'd5271: dataIn2 = 32'd1; 
32'd5272: dataIn2 = 32'd0; 
32'd5273: dataIn2 = 32'd1; 
32'd5274: dataIn2 = 32'd0; 
32'd5275: dataIn2 = 32'd1; 
32'd5276: dataIn2 = 32'd1; 
32'd5277: dataIn2 = 32'd1; 
32'd5278: dataIn2 = 32'd1; 
32'd5279: dataIn2 = 32'd0; 
32'd5280: dataIn2 = 32'd0; 
32'd5281: dataIn2 = 32'd0; 
32'd5282: dataIn2 = 32'd0; 
32'd5283: dataIn2 = 32'd1; 
32'd5284: dataIn2 = 32'd0; 
32'd5285: dataIn2 = 32'd0; 
32'd5286: dataIn2 = 32'd0; 
32'd5287: dataIn2 = 32'd0; 
32'd5288: dataIn2 = 32'd1; 
32'd5289: dataIn2 = 32'd1; 
32'd5290: dataIn2 = 32'd0; 
32'd5291: dataIn2 = 32'd0; 
32'd5292: dataIn2 = 32'd1; 
32'd5293: dataIn2 = 32'd0; 
32'd5294: dataIn2 = 32'd1; 
32'd5295: dataIn2 = 32'd0; 
32'd5296: dataIn2 = 32'd1; 
32'd5297: dataIn2 = 32'd1; 
32'd5298: dataIn2 = 32'd1; 
32'd5299: dataIn2 = 32'd0; 
32'd5300: dataIn2 = 32'd1; 
32'd5301: dataIn2 = 32'd0; 
32'd5302: dataIn2 = 32'd1; 
32'd5303: dataIn2 = 32'd0; 
32'd5304: dataIn2 = 32'd0; 
32'd5305: dataIn2 = 32'd1; 
32'd5306: dataIn2 = 32'd1; 
32'd5307: dataIn2 = 32'd0; 
32'd5308: dataIn2 = 32'd1; 
32'd5309: dataIn2 = 32'd1; 
32'd5310: dataIn2 = 32'd1; 
32'd5311: dataIn2 = 32'd0; 
32'd5312: dataIn2 = 32'd1; 
32'd5313: dataIn2 = 32'd0; 
32'd5314: dataIn2 = 32'd0; 
32'd5315: dataIn2 = 32'd0; 
32'd5316: dataIn2 = 32'd1; 
32'd5317: dataIn2 = 32'd1; 
32'd5318: dataIn2 = 32'd1; 
32'd5319: dataIn2 = 32'd1; 
32'd5320: dataIn2 = 32'd1; 
32'd5321: dataIn2 = 32'd0; 
32'd5322: dataIn2 = 32'd1; 
32'd5323: dataIn2 = 32'd1; 
32'd5324: dataIn2 = 32'd1; 
32'd5325: dataIn2 = 32'd1; 
32'd5326: dataIn2 = 32'd1; 
32'd5327: dataIn2 = 32'd0; 
32'd5328: dataIn2 = 32'd1; 
32'd5329: dataIn2 = 32'd1; 
32'd5330: dataIn2 = 32'd0; 
32'd5331: dataIn2 = 32'd1; 
32'd5332: dataIn2 = 32'd0; 
32'd5333: dataIn2 = 32'd0; 
32'd5334: dataIn2 = 32'd0; 
32'd5335: dataIn2 = 32'd1; 
32'd5336: dataIn2 = 32'd1; 
32'd5337: dataIn2 = 32'd1; 
32'd5338: dataIn2 = 32'd1; 
32'd5339: dataIn2 = 32'd0; 
32'd5340: dataIn2 = 32'd0; 
32'd5341: dataIn2 = 32'd0; 
32'd5342: dataIn2 = 32'd0; 
32'd5343: dataIn2 = 32'd1; 
32'd5344: dataIn2 = 32'd1; 
32'd5345: dataIn2 = 32'd1; 
32'd5346: dataIn2 = 32'd1; 
32'd5347: dataIn2 = 32'd0; 
32'd5348: dataIn2 = 32'd0; 
32'd5349: dataIn2 = 32'd0; 
32'd5350: dataIn2 = 32'd1; 
32'd5351: dataIn2 = 32'd1; 
32'd5352: dataIn2 = 32'd0; 
32'd5353: dataIn2 = 32'd0; 
32'd5354: dataIn2 = 32'd0; 
32'd5355: dataIn2 = 32'd0; 
32'd5356: dataIn2 = 32'd0; 
32'd5357: dataIn2 = 32'd1; 
32'd5358: dataIn2 = 32'd0; 
32'd5359: dataIn2 = 32'd1; 
32'd5360: dataIn2 = 32'd0; 
32'd5361: dataIn2 = 32'd1; 
32'd5362: dataIn2 = 32'd1; 
32'd5363: dataIn2 = 32'd0; 
32'd5364: dataIn2 = 32'd0; 
32'd5365: dataIn2 = 32'd0; 
32'd5366: dataIn2 = 32'd1; 
32'd5367: dataIn2 = 32'd0; 
32'd5368: dataIn2 = 32'd0; 
32'd5369: dataIn2 = 32'd1; 
32'd5370: dataIn2 = 32'd0; 
32'd5371: dataIn2 = 32'd1; 
32'd5372: dataIn2 = 32'd0; 
32'd5373: dataIn2 = 32'd1; 
32'd5374: dataIn2 = 32'd1; 
32'd5375: dataIn2 = 32'd1; 
32'd5376: dataIn2 = 32'd1; 
32'd5377: dataIn2 = 32'd0; 
32'd5378: dataIn2 = 32'd0; 
32'd5379: dataIn2 = 32'd0; 
32'd5380: dataIn2 = 32'd0; 
32'd5381: dataIn2 = 32'd0; 
32'd5382: dataIn2 = 32'd0; 
32'd5383: dataIn2 = 32'd0; 
32'd5384: dataIn2 = 32'd1; 
32'd5385: dataIn2 = 32'd0; 
32'd5386: dataIn2 = 32'd1; 
32'd5387: dataIn2 = 32'd0; 
32'd5388: dataIn2 = 32'd1; 
32'd5389: dataIn2 = 32'd0; 
32'd5390: dataIn2 = 32'd1; 
32'd5391: dataIn2 = 32'd1; 
32'd5392: dataIn2 = 32'd1; 
32'd5393: dataIn2 = 32'd0; 
32'd5394: dataIn2 = 32'd1; 
32'd5395: dataIn2 = 32'd0; 
32'd5396: dataIn2 = 32'd0; 
32'd5397: dataIn2 = 32'd1; 
32'd5398: dataIn2 = 32'd1; 
32'd5399: dataIn2 = 32'd1; 
32'd5400: dataIn2 = 32'd0; 
32'd5401: dataIn2 = 32'd0; 
32'd5402: dataIn2 = 32'd1; 
32'd5403: dataIn2 = 32'd1; 
32'd5404: dataIn2 = 32'd1; 
32'd5405: dataIn2 = 32'd1; 
32'd5406: dataIn2 = 32'd1; 
32'd5407: dataIn2 = 32'd0; 
32'd5408: dataIn2 = 32'd1; 
32'd5409: dataIn2 = 32'd0; 
32'd5410: dataIn2 = 32'd0; 
32'd5411: dataIn2 = 32'd0; 
32'd5412: dataIn2 = 32'd1; 
32'd5413: dataIn2 = 32'd1; 
32'd5414: dataIn2 = 32'd1; 
32'd5415: dataIn2 = 32'd1; 
32'd5416: dataIn2 = 32'd0; 
32'd5417: dataIn2 = 32'd0; 
32'd5418: dataIn2 = 32'd0; 
32'd5419: dataIn2 = 32'd0; 
32'd5420: dataIn2 = 32'd1; 
32'd5421: dataIn2 = 32'd0; 
32'd5422: dataIn2 = 32'd1; 
32'd5423: dataIn2 = 32'd1; 
32'd5424: dataIn2 = 32'd1; 
32'd5425: dataIn2 = 32'd1; 
32'd5426: dataIn2 = 32'd1; 
32'd5427: dataIn2 = 32'd1; 
32'd5428: dataIn2 = 32'd0; 
32'd5429: dataIn2 = 32'd0; 
32'd5430: dataIn2 = 32'd0; 
32'd5431: dataIn2 = 32'd1; 
32'd5432: dataIn2 = 32'd1; 
32'd5433: dataIn2 = 32'd0; 
32'd5434: dataIn2 = 32'd1; 
32'd5435: dataIn2 = 32'd0; 
32'd5436: dataIn2 = 32'd0; 
32'd5437: dataIn2 = 32'd1; 
32'd5438: dataIn2 = 32'd1; 
32'd5439: dataIn2 = 32'd0; 
32'd5440: dataIn2 = 32'd1; 
32'd5441: dataIn2 = 32'd1; 
32'd5442: dataIn2 = 32'd1; 
32'd5443: dataIn2 = 32'd0; 
32'd5444: dataIn2 = 32'd0; 
32'd5445: dataIn2 = 32'd1; 
32'd5446: dataIn2 = 32'd1; 
32'd5447: dataIn2 = 32'd0; 
32'd5448: dataIn2 = 32'd0; 
32'd5449: dataIn2 = 32'd0; 
32'd5450: dataIn2 = 32'd0; 
32'd5451: dataIn2 = 32'd0; 
32'd5452: dataIn2 = 32'd0; 
32'd5453: dataIn2 = 32'd0; 
32'd5454: dataIn2 = 32'd1; 
32'd5455: dataIn2 = 32'd1; 
32'd5456: dataIn2 = 32'd1; 
32'd5457: dataIn2 = 32'd1; 
32'd5458: dataIn2 = 32'd1; 
32'd5459: dataIn2 = 32'd1; 
32'd5460: dataIn2 = 32'd0; 
32'd5461: dataIn2 = 32'd0; 
32'd5462: dataIn2 = 32'd0; 
32'd5463: dataIn2 = 32'd0; 
32'd5464: dataIn2 = 32'd0; 
32'd5465: dataIn2 = 32'd1; 
32'd5466: dataIn2 = 32'd0; 
32'd5467: dataIn2 = 32'd1; 
32'd5468: dataIn2 = 32'd0; 
32'd5469: dataIn2 = 32'd0; 
32'd5470: dataIn2 = 32'd0; 
32'd5471: dataIn2 = 32'd0; 
32'd5472: dataIn2 = 32'd0; 
32'd5473: dataIn2 = 32'd1; 
32'd5474: dataIn2 = 32'd1; 
32'd5475: dataIn2 = 32'd0; 
32'd5476: dataIn2 = 32'd0; 
32'd5477: dataIn2 = 32'd1; 
32'd5478: dataIn2 = 32'd0; 
32'd5479: dataIn2 = 32'd1; 
32'd5480: dataIn2 = 32'd1; 
32'd5481: dataIn2 = 32'd0; 
32'd5482: dataIn2 = 32'd1; 
32'd5483: dataIn2 = 32'd0; 
32'd5484: dataIn2 = 32'd1; 
32'd5485: dataIn2 = 32'd1; 
32'd5486: dataIn2 = 32'd0; 
32'd5487: dataIn2 = 32'd0; 
32'd5488: dataIn2 = 32'd1; 
32'd5489: dataIn2 = 32'd0; 
32'd5490: dataIn2 = 32'd1; 
32'd5491: dataIn2 = 32'd0; 
32'd5492: dataIn2 = 32'd0; 
32'd5493: dataIn2 = 32'd0; 
32'd5494: dataIn2 = 32'd0; 
32'd5495: dataIn2 = 32'd1; 
32'd5496: dataIn2 = 32'd1; 
32'd5497: dataIn2 = 32'd0; 
32'd5498: dataIn2 = 32'd1; 
32'd5499: dataIn2 = 32'd0; 
32'd5500: dataIn2 = 32'd0; 
32'd5501: dataIn2 = 32'd0; 
32'd5502: dataIn2 = 32'd1; 
32'd5503: dataIn2 = 32'd1; 
32'd5504: dataIn2 = 32'd1; 
32'd5505: dataIn2 = 32'd0; 
32'd5506: dataIn2 = 32'd0; 
32'd5507: dataIn2 = 32'd0; 
32'd5508: dataIn2 = 32'd1; 
32'd5509: dataIn2 = 32'd1; 
32'd5510: dataIn2 = 32'd0; 
32'd5511: dataIn2 = 32'd1; 
32'd5512: dataIn2 = 32'd0; 
32'd5513: dataIn2 = 32'd1; 
32'd5514: dataIn2 = 32'd1; 
32'd5515: dataIn2 = 32'd0; 
32'd5516: dataIn2 = 32'd0; 
32'd5517: dataIn2 = 32'd0; 
32'd5518: dataIn2 = 32'd0; 
32'd5519: dataIn2 = 32'd1; 
32'd5520: dataIn2 = 32'd1; 
32'd5521: dataIn2 = 32'd1; 
32'd5522: dataIn2 = 32'd1; 
32'd5523: dataIn2 = 32'd1; 
32'd5524: dataIn2 = 32'd1; 
32'd5525: dataIn2 = 32'd1; 
32'd5526: dataIn2 = 32'd0; 
32'd5527: dataIn2 = 32'd1; 
32'd5528: dataIn2 = 32'd0; 
32'd5529: dataIn2 = 32'd1; 
32'd5530: dataIn2 = 32'd0; 
32'd5531: dataIn2 = 32'd1; 
32'd5532: dataIn2 = 32'd1; 
32'd5533: dataIn2 = 32'd1; 
32'd5534: dataIn2 = 32'd1; 
32'd5535: dataIn2 = 32'd1; 
32'd5536: dataIn2 = 32'd0; 
32'd5537: dataIn2 = 32'd0; 
32'd5538: dataIn2 = 32'd1; 
32'd5539: dataIn2 = 32'd1; 
32'd5540: dataIn2 = 32'd0; 
32'd5541: dataIn2 = 32'd0; 
32'd5542: dataIn2 = 32'd0; 
32'd5543: dataIn2 = 32'd1; 
32'd5544: dataIn2 = 32'd1; 
32'd5545: dataIn2 = 32'd1; 
32'd5546: dataIn2 = 32'd0; 
32'd5547: dataIn2 = 32'd1; 
32'd5548: dataIn2 = 32'd0; 
32'd5549: dataIn2 = 32'd0; 
32'd5550: dataIn2 = 32'd0; 
32'd5551: dataIn2 = 32'd0; 
32'd5552: dataIn2 = 32'd1; 
32'd5553: dataIn2 = 32'd0; 
32'd5554: dataIn2 = 32'd0; 
32'd5555: dataIn2 = 32'd0; 
32'd5556: dataIn2 = 32'd0; 
32'd5557: dataIn2 = 32'd0; 
32'd5558: dataIn2 = 32'd0; 
32'd5559: dataIn2 = 32'd0; 
32'd5560: dataIn2 = 32'd1; 
32'd5561: dataIn2 = 32'd1; 
32'd5562: dataIn2 = 32'd1; 
32'd5563: dataIn2 = 32'd0; 
32'd5564: dataIn2 = 32'd0; 
32'd5565: dataIn2 = 32'd1; 
32'd5566: dataIn2 = 32'd0; 
32'd5567: dataIn2 = 32'd1; 
32'd5568: dataIn2 = 32'd1; 
32'd5569: dataIn2 = 32'd1; 
32'd5570: dataIn2 = 32'd0; 
32'd5571: dataIn2 = 32'd0; 
32'd5572: dataIn2 = 32'd0; 
32'd5573: dataIn2 = 32'd0; 
32'd5574: dataIn2 = 32'd0; 
32'd5575: dataIn2 = 32'd0; 
32'd5576: dataIn2 = 32'd0; 
32'd5577: dataIn2 = 32'd0; 
32'd5578: dataIn2 = 32'd0; 
32'd5579: dataIn2 = 32'd0; 
32'd5580: dataIn2 = 32'd0; 
32'd5581: dataIn2 = 32'd0; 
32'd5582: dataIn2 = 32'd0; 
32'd5583: dataIn2 = 32'd0; 
32'd5584: dataIn2 = 32'd1; 
32'd5585: dataIn2 = 32'd0; 
32'd5586: dataIn2 = 32'd0; 
32'd5587: dataIn2 = 32'd0; 
32'd5588: dataIn2 = 32'd0; 
32'd5589: dataIn2 = 32'd0; 
32'd5590: dataIn2 = 32'd1; 
32'd5591: dataIn2 = 32'd0; 
32'd5592: dataIn2 = 32'd0; 
32'd5593: dataIn2 = 32'd1; 
32'd5594: dataIn2 = 32'd0; 
32'd5595: dataIn2 = 32'd0; 
32'd5596: dataIn2 = 32'd1; 
32'd5597: dataIn2 = 32'd0; 
32'd5598: dataIn2 = 32'd1; 
32'd5599: dataIn2 = 32'd0; 
32'd5600: dataIn2 = 32'd0; 
32'd5601: dataIn2 = 32'd0; 
32'd5602: dataIn2 = 32'd1; 
32'd5603: dataIn2 = 32'd0; 
32'd5604: dataIn2 = 32'd0; 
32'd5605: dataIn2 = 32'd1; 
32'd5606: dataIn2 = 32'd0; 
32'd5607: dataIn2 = 32'd1; 
32'd5608: dataIn2 = 32'd0; 
32'd5609: dataIn2 = 32'd1; 
32'd5610: dataIn2 = 32'd0; 
32'd5611: dataIn2 = 32'd1; 
32'd5612: dataIn2 = 32'd1; 
32'd5613: dataIn2 = 32'd1; 
32'd5614: dataIn2 = 32'd0; 
32'd5615: dataIn2 = 32'd0; 
32'd5616: dataIn2 = 32'd0; 
32'd5617: dataIn2 = 32'd0; 
32'd5618: dataIn2 = 32'd0; 
32'd5619: dataIn2 = 32'd0; 
32'd5620: dataIn2 = 32'd0; 
32'd5621: dataIn2 = 32'd1; 
32'd5622: dataIn2 = 32'd1; 
32'd5623: dataIn2 = 32'd1; 
32'd5624: dataIn2 = 32'd1; 
32'd5625: dataIn2 = 32'd0; 
32'd5626: dataIn2 = 32'd1; 
32'd5627: dataIn2 = 32'd0; 
32'd5628: dataIn2 = 32'd1; 
32'd5629: dataIn2 = 32'd1; 
32'd5630: dataIn2 = 32'd0; 
32'd5631: dataIn2 = 32'd1; 
32'd5632: dataIn2 = 32'd0; 
32'd5633: dataIn2 = 32'd0; 
32'd5634: dataIn2 = 32'd1; 
32'd5635: dataIn2 = 32'd0; 
32'd5636: dataIn2 = 32'd0; 
32'd5637: dataIn2 = 32'd0; 
32'd5638: dataIn2 = 32'd0; 
32'd5639: dataIn2 = 32'd0; 
32'd5640: dataIn2 = 32'd1; 
32'd5641: dataIn2 = 32'd0; 
32'd5642: dataIn2 = 32'd1; 
32'd5643: dataIn2 = 32'd0; 
32'd5644: dataIn2 = 32'd1; 
32'd5645: dataIn2 = 32'd0; 
32'd5646: dataIn2 = 32'd1; 
32'd5647: dataIn2 = 32'd1; 
32'd5648: dataIn2 = 32'd1; 
32'd5649: dataIn2 = 32'd1; 
32'd5650: dataIn2 = 32'd1; 
32'd5651: dataIn2 = 32'd0; 
32'd5652: dataIn2 = 32'd1; 
32'd5653: dataIn2 = 32'd0; 
32'd5654: dataIn2 = 32'd0; 
32'd5655: dataIn2 = 32'd0; 
32'd5656: dataIn2 = 32'd1; 
32'd5657: dataIn2 = 32'd1; 
32'd5658: dataIn2 = 32'd1; 
32'd5659: dataIn2 = 32'd1; 
32'd5660: dataIn2 = 32'd0; 
32'd5661: dataIn2 = 32'd0; 
32'd5662: dataIn2 = 32'd1; 
32'd5663: dataIn2 = 32'd1; 
32'd5664: dataIn2 = 32'd1; 
32'd5665: dataIn2 = 32'd0; 
32'd5666: dataIn2 = 32'd0; 
32'd5667: dataIn2 = 32'd0; 
32'd5668: dataIn2 = 32'd0; 
32'd5669: dataIn2 = 32'd1; 
32'd5670: dataIn2 = 32'd1; 
32'd5671: dataIn2 = 32'd1; 
32'd5672: dataIn2 = 32'd1; 
32'd5673: dataIn2 = 32'd0; 
32'd5674: dataIn2 = 32'd1; 
32'd5675: dataIn2 = 32'd1; 
32'd5676: dataIn2 = 32'd1; 
32'd5677: dataIn2 = 32'd1; 
32'd5678: dataIn2 = 32'd0; 
32'd5679: dataIn2 = 32'd0; 
32'd5680: dataIn2 = 32'd0; 
32'd5681: dataIn2 = 32'd0; 
32'd5682: dataIn2 = 32'd1; 
32'd5683: dataIn2 = 32'd0; 
32'd5684: dataIn2 = 32'd0; 
32'd5685: dataIn2 = 32'd0; 
32'd5686: dataIn2 = 32'd1; 
32'd5687: dataIn2 = 32'd1; 
32'd5688: dataIn2 = 32'd1; 
32'd5689: dataIn2 = 32'd1; 
32'd5690: dataIn2 = 32'd1; 
32'd5691: dataIn2 = 32'd1; 
32'd5692: dataIn2 = 32'd0; 
32'd5693: dataIn2 = 32'd0; 
32'd5694: dataIn2 = 32'd1; 
32'd5695: dataIn2 = 32'd0; 
32'd5696: dataIn2 = 32'd1; 
32'd5697: dataIn2 = 32'd1; 
32'd5698: dataIn2 = 32'd1; 
32'd5699: dataIn2 = 32'd1; 
32'd5700: dataIn2 = 32'd0; 
32'd5701: dataIn2 = 32'd1; 
32'd5702: dataIn2 = 32'd1; 
32'd5703: dataIn2 = 32'd1; 
32'd5704: dataIn2 = 32'd1; 
32'd5705: dataIn2 = 32'd1; 
32'd5706: dataIn2 = 32'd0; 
32'd5707: dataIn2 = 32'd1; 
32'd5708: dataIn2 = 32'd1; 
32'd5709: dataIn2 = 32'd0; 
32'd5710: dataIn2 = 32'd1; 
32'd5711: dataIn2 = 32'd1; 
32'd5712: dataIn2 = 32'd1; 
32'd5713: dataIn2 = 32'd1; 
32'd5714: dataIn2 = 32'd1; 
32'd5715: dataIn2 = 32'd1; 
32'd5716: dataIn2 = 32'd0; 
32'd5717: dataIn2 = 32'd0; 
32'd5718: dataIn2 = 32'd1; 
32'd5719: dataIn2 = 32'd0; 
32'd5720: dataIn2 = 32'd1; 
32'd5721: dataIn2 = 32'd1; 
32'd5722: dataIn2 = 32'd0; 
32'd5723: dataIn2 = 32'd1; 
32'd5724: dataIn2 = 32'd0; 
32'd5725: dataIn2 = 32'd1; 
32'd5726: dataIn2 = 32'd0; 
32'd5727: dataIn2 = 32'd1; 
32'd5728: dataIn2 = 32'd1; 
32'd5729: dataIn2 = 32'd0; 
32'd5730: dataIn2 = 32'd0; 
32'd5731: dataIn2 = 32'd1; 
32'd5732: dataIn2 = 32'd0; 
32'd5733: dataIn2 = 32'd1; 
32'd5734: dataIn2 = 32'd0; 
32'd5735: dataIn2 = 32'd1; 
32'd5736: dataIn2 = 32'd1; 
32'd5737: dataIn2 = 32'd1; 
32'd5738: dataIn2 = 32'd0; 
32'd5739: dataIn2 = 32'd0; 
32'd5740: dataIn2 = 32'd0; 
32'd5741: dataIn2 = 32'd1; 
32'd5742: dataIn2 = 32'd1; 
32'd5743: dataIn2 = 32'd1; 
32'd5744: dataIn2 = 32'd0; 
32'd5745: dataIn2 = 32'd1; 
32'd5746: dataIn2 = 32'd1; 
32'd5747: dataIn2 = 32'd0; 
32'd5748: dataIn2 = 32'd0; 
32'd5749: dataIn2 = 32'd0; 
32'd5750: dataIn2 = 32'd1; 
32'd5751: dataIn2 = 32'd1; 
32'd5752: dataIn2 = 32'd1; 
32'd5753: dataIn2 = 32'd0; 
32'd5754: dataIn2 = 32'd1; 
32'd5755: dataIn2 = 32'd1; 
32'd5756: dataIn2 = 32'd1; 
32'd5757: dataIn2 = 32'd0; 
32'd5758: dataIn2 = 32'd1; 
32'd5759: dataIn2 = 32'd0; 
32'd5760: dataIn2 = 32'd0; 
32'd5761: dataIn2 = 32'd1; 
32'd5762: dataIn2 = 32'd0; 
32'd5763: dataIn2 = 32'd0; 
32'd5764: dataIn2 = 32'd1; 
32'd5765: dataIn2 = 32'd1; 
32'd5766: dataIn2 = 32'd0; 
32'd5767: dataIn2 = 32'd0; 
32'd5768: dataIn2 = 32'd0; 
32'd5769: dataIn2 = 32'd1; 
32'd5770: dataIn2 = 32'd1; 
32'd5771: dataIn2 = 32'd1; 
32'd5772: dataIn2 = 32'd1; 
32'd5773: dataIn2 = 32'd1; 
32'd5774: dataIn2 = 32'd0; 
32'd5775: dataIn2 = 32'd1; 
32'd5776: dataIn2 = 32'd1; 
32'd5777: dataIn2 = 32'd0; 
32'd5778: dataIn2 = 32'd0; 
32'd5779: dataIn2 = 32'd0; 
32'd5780: dataIn2 = 32'd0; 
32'd5781: dataIn2 = 32'd1; 
32'd5782: dataIn2 = 32'd1; 
32'd5783: dataIn2 = 32'd0; 
32'd5784: dataIn2 = 32'd1; 
32'd5785: dataIn2 = 32'd0; 
32'd5786: dataIn2 = 32'd0; 
32'd5787: dataIn2 = 32'd1; 
32'd5788: dataIn2 = 32'd1; 
32'd5789: dataIn2 = 32'd1; 
32'd5790: dataIn2 = 32'd0; 
32'd5791: dataIn2 = 32'd1; 
32'd5792: dataIn2 = 32'd1; 
32'd5793: dataIn2 = 32'd1; 
32'd5794: dataIn2 = 32'd0; 
32'd5795: dataIn2 = 32'd0; 
32'd5796: dataIn2 = 32'd1; 
32'd5797: dataIn2 = 32'd1; 
32'd5798: dataIn2 = 32'd1; 
32'd5799: dataIn2 = 32'd0; 
32'd5800: dataIn2 = 32'd0; 
32'd5801: dataIn2 = 32'd1; 
32'd5802: dataIn2 = 32'd0; 
32'd5803: dataIn2 = 32'd1; 
32'd5804: dataIn2 = 32'd0; 
32'd5805: dataIn2 = 32'd1; 
32'd5806: dataIn2 = 32'd0; 
32'd5807: dataIn2 = 32'd0; 
32'd5808: dataIn2 = 32'd1; 
32'd5809: dataIn2 = 32'd0; 
32'd5810: dataIn2 = 32'd0; 
32'd5811: dataIn2 = 32'd1; 
32'd5812: dataIn2 = 32'd0; 
32'd5813: dataIn2 = 32'd0; 
32'd5814: dataIn2 = 32'd0; 
32'd5815: dataIn2 = 32'd0; 
32'd5816: dataIn2 = 32'd1; 
32'd5817: dataIn2 = 32'd0; 
32'd5818: dataIn2 = 32'd0; 
32'd5819: dataIn2 = 32'd0; 
32'd5820: dataIn2 = 32'd0; 
32'd5821: dataIn2 = 32'd0; 
32'd5822: dataIn2 = 32'd1; 
32'd5823: dataIn2 = 32'd1; 
32'd5824: dataIn2 = 32'd0; 
32'd5825: dataIn2 = 32'd0; 
32'd5826: dataIn2 = 32'd1; 
32'd5827: dataIn2 = 32'd1; 
32'd5828: dataIn2 = 32'd1; 
32'd5829: dataIn2 = 32'd1; 
32'd5830: dataIn2 = 32'd1; 
32'd5831: dataIn2 = 32'd1; 
32'd5832: dataIn2 = 32'd1; 
32'd5833: dataIn2 = 32'd1; 
32'd5834: dataIn2 = 32'd0; 
32'd5835: dataIn2 = 32'd0; 
32'd5836: dataIn2 = 32'd0; 
32'd5837: dataIn2 = 32'd1; 
32'd5838: dataIn2 = 32'd1; 
32'd5839: dataIn2 = 32'd1; 
32'd5840: dataIn2 = 32'd1; 
32'd5841: dataIn2 = 32'd1; 
32'd5842: dataIn2 = 32'd1; 
32'd5843: dataIn2 = 32'd1; 
32'd5844: dataIn2 = 32'd1; 
32'd5845: dataIn2 = 32'd1; 
32'd5846: dataIn2 = 32'd1; 
32'd5847: dataIn2 = 32'd0; 
32'd5848: dataIn2 = 32'd0; 
32'd5849: dataIn2 = 32'd1; 
32'd5850: dataIn2 = 32'd1; 
32'd5851: dataIn2 = 32'd1; 
32'd5852: dataIn2 = 32'd0; 
32'd5853: dataIn2 = 32'd0; 
32'd5854: dataIn2 = 32'd0; 
32'd5855: dataIn2 = 32'd0; 
32'd5856: dataIn2 = 32'd1; 
32'd5857: dataIn2 = 32'd0; 
32'd5858: dataIn2 = 32'd0; 
32'd5859: dataIn2 = 32'd0; 
32'd5860: dataIn2 = 32'd1; 
32'd5861: dataIn2 = 32'd1; 
32'd5862: dataIn2 = 32'd1; 
32'd5863: dataIn2 = 32'd0; 
32'd5864: dataIn2 = 32'd0; 
32'd5865: dataIn2 = 32'd0; 
32'd5866: dataIn2 = 32'd0; 
32'd5867: dataIn2 = 32'd0; 
32'd5868: dataIn2 = 32'd1; 
32'd5869: dataIn2 = 32'd0; 
32'd5870: dataIn2 = 32'd1; 
32'd5871: dataIn2 = 32'd1; 
32'd5872: dataIn2 = 32'd0; 
32'd5873: dataIn2 = 32'd0; 
32'd5874: dataIn2 = 32'd1; 
32'd5875: dataIn2 = 32'd1; 
32'd5876: dataIn2 = 32'd1; 
32'd5877: dataIn2 = 32'd0; 
32'd5878: dataIn2 = 32'd1; 
32'd5879: dataIn2 = 32'd0; 
32'd5880: dataIn2 = 32'd1; 
32'd5881: dataIn2 = 32'd1; 
32'd5882: dataIn2 = 32'd0; 
32'd5883: dataIn2 = 32'd0; 
32'd5884: dataIn2 = 32'd0; 
32'd5885: dataIn2 = 32'd0; 
32'd5886: dataIn2 = 32'd1; 
32'd5887: dataIn2 = 32'd1; 
32'd5888: dataIn2 = 32'd0; 
32'd5889: dataIn2 = 32'd1; 
32'd5890: dataIn2 = 32'd1; 
32'd5891: dataIn2 = 32'd0; 
32'd5892: dataIn2 = 32'd1; 
32'd5893: dataIn2 = 32'd0; 
32'd5894: dataIn2 = 32'd0; 
32'd5895: dataIn2 = 32'd0; 
32'd5896: dataIn2 = 32'd0; 
32'd5897: dataIn2 = 32'd0; 
32'd5898: dataIn2 = 32'd1; 
32'd5899: dataIn2 = 32'd1; 
32'd5900: dataIn2 = 32'd1; 
32'd5901: dataIn2 = 32'd1; 
32'd5902: dataIn2 = 32'd0; 
32'd5903: dataIn2 = 32'd1; 
32'd5904: dataIn2 = 32'd1; 
32'd5905: dataIn2 = 32'd0; 
32'd5906: dataIn2 = 32'd1; 
32'd5907: dataIn2 = 32'd0; 
32'd5908: dataIn2 = 32'd1; 
32'd5909: dataIn2 = 32'd0; 
32'd5910: dataIn2 = 32'd0; 
32'd5911: dataIn2 = 32'd1; 
32'd5912: dataIn2 = 32'd1; 
32'd5913: dataIn2 = 32'd1; 
32'd5914: dataIn2 = 32'd1; 
32'd5915: dataIn2 = 32'd1; 
32'd5916: dataIn2 = 32'd0; 
32'd5917: dataIn2 = 32'd0; 
32'd5918: dataIn2 = 32'd1; 
32'd5919: dataIn2 = 32'd0; 
32'd5920: dataIn2 = 32'd0; 
32'd5921: dataIn2 = 32'd1; 
32'd5922: dataIn2 = 32'd0; 
32'd5923: dataIn2 = 32'd1; 
32'd5924: dataIn2 = 32'd0; 
32'd5925: dataIn2 = 32'd1; 
32'd5926: dataIn2 = 32'd0; 
32'd5927: dataIn2 = 32'd1; 
32'd5928: dataIn2 = 32'd1; 
32'd5929: dataIn2 = 32'd1; 
32'd5930: dataIn2 = 32'd1; 
32'd5931: dataIn2 = 32'd0; 
32'd5932: dataIn2 = 32'd0; 
32'd5933: dataIn2 = 32'd1; 
32'd5934: dataIn2 = 32'd1; 
32'd5935: dataIn2 = 32'd0; 
32'd5936: dataIn2 = 32'd0; 
32'd5937: dataIn2 = 32'd0; 
32'd5938: dataIn2 = 32'd1; 
32'd5939: dataIn2 = 32'd0; 
32'd5940: dataIn2 = 32'd0; 
32'd5941: dataIn2 = 32'd0; 
32'd5942: dataIn2 = 32'd1; 
32'd5943: dataIn2 = 32'd1; 
32'd5944: dataIn2 = 32'd1; 
32'd5945: dataIn2 = 32'd0; 
32'd5946: dataIn2 = 32'd1; 
32'd5947: dataIn2 = 32'd0; 
32'd5948: dataIn2 = 32'd1; 
32'd5949: dataIn2 = 32'd0; 
32'd5950: dataIn2 = 32'd0; 
32'd5951: dataIn2 = 32'd0; 
32'd5952: dataIn2 = 32'd1; 
32'd5953: dataIn2 = 32'd0; 
32'd5954: dataIn2 = 32'd1; 
32'd5955: dataIn2 = 32'd1; 
32'd5956: dataIn2 = 32'd1; 
32'd5957: dataIn2 = 32'd1; 
32'd5958: dataIn2 = 32'd1; 
32'd5959: dataIn2 = 32'd0; 
32'd5960: dataIn2 = 32'd1; 
32'd5961: dataIn2 = 32'd1; 
32'd5962: dataIn2 = 32'd1; 
32'd5963: dataIn2 = 32'd0; 
32'd5964: dataIn2 = 32'd1; 
32'd5965: dataIn2 = 32'd0; 
32'd5966: dataIn2 = 32'd0; 
32'd5967: dataIn2 = 32'd1; 
32'd5968: dataIn2 = 32'd1; 
32'd5969: dataIn2 = 32'd1; 
32'd5970: dataIn2 = 32'd0; 
32'd5971: dataIn2 = 32'd0; 
32'd5972: dataIn2 = 32'd0; 
32'd5973: dataIn2 = 32'd1; 
32'd5974: dataIn2 = 32'd0; 
32'd5975: dataIn2 = 32'd0; 
32'd5976: dataIn2 = 32'd1; 
32'd5977: dataIn2 = 32'd0; 
32'd5978: dataIn2 = 32'd1; 
32'd5979: dataIn2 = 32'd1; 
32'd5980: dataIn2 = 32'd0; 
32'd5981: dataIn2 = 32'd0; 
32'd5982: dataIn2 = 32'd0; 
32'd5983: dataIn2 = 32'd1; 
32'd5984: dataIn2 = 32'd0; 
32'd5985: dataIn2 = 32'd1; 
32'd5986: dataIn2 = 32'd1; 
32'd5987: dataIn2 = 32'd0; 
32'd5988: dataIn2 = 32'd1; 
32'd5989: dataIn2 = 32'd0; 
32'd5990: dataIn2 = 32'd1; 
32'd5991: dataIn2 = 32'd1; 
32'd5992: dataIn2 = 32'd0; 
32'd5993: dataIn2 = 32'd1; 
32'd5994: dataIn2 = 32'd0; 
32'd5995: dataIn2 = 32'd1; 
32'd5996: dataIn2 = 32'd1; 
32'd5997: dataIn2 = 32'd0; 
32'd5998: dataIn2 = 32'd0; 
32'd5999: dataIn2 = 32'd1; 
32'd6000: dataIn2 = 32'd0; 
32'd6001: dataIn2 = 32'd0; 
32'd6002: dataIn2 = 32'd1; 
32'd6003: dataIn2 = 32'd1; 
32'd6004: dataIn2 = 32'd1; 
32'd6005: dataIn2 = 32'd1; 
32'd6006: dataIn2 = 32'd0; 
32'd6007: dataIn2 = 32'd1; 
32'd6008: dataIn2 = 32'd1; 
32'd6009: dataIn2 = 32'd1; 
32'd6010: dataIn2 = 32'd0; 
32'd6011: dataIn2 = 32'd1; 
32'd6012: dataIn2 = 32'd0; 
32'd6013: dataIn2 = 32'd0; 
32'd6014: dataIn2 = 32'd0; 
32'd6015: dataIn2 = 32'd0; 
32'd6016: dataIn2 = 32'd0; 
32'd6017: dataIn2 = 32'd0; 
32'd6018: dataIn2 = 32'd0; 
32'd6019: dataIn2 = 32'd0; 
32'd6020: dataIn2 = 32'd1; 
32'd6021: dataIn2 = 32'd0; 
32'd6022: dataIn2 = 32'd1; 
32'd6023: dataIn2 = 32'd0; 
32'd6024: dataIn2 = 32'd1; 
32'd6025: dataIn2 = 32'd1; 
32'd6026: dataIn2 = 32'd0; 
32'd6027: dataIn2 = 32'd0; 
32'd6028: dataIn2 = 32'd1; 
32'd6029: dataIn2 = 32'd0; 
32'd6030: dataIn2 = 32'd1; 
32'd6031: dataIn2 = 32'd0; 
32'd6032: dataIn2 = 32'd1; 
32'd6033: dataIn2 = 32'd1; 
32'd6034: dataIn2 = 32'd1; 
32'd6035: dataIn2 = 32'd1; 
32'd6036: dataIn2 = 32'd1; 
32'd6037: dataIn2 = 32'd1; 
32'd6038: dataIn2 = 32'd0; 
32'd6039: dataIn2 = 32'd0; 
32'd6040: dataIn2 = 32'd1; 
32'd6041: dataIn2 = 32'd1; 
32'd6042: dataIn2 = 32'd1; 
32'd6043: dataIn2 = 32'd0; 
32'd6044: dataIn2 = 32'd1; 
32'd6045: dataIn2 = 32'd0; 
32'd6046: dataIn2 = 32'd0; 
32'd6047: dataIn2 = 32'd1; 
32'd6048: dataIn2 = 32'd1; 
32'd6049: dataIn2 = 32'd1; 
32'd6050: dataIn2 = 32'd0; 
32'd6051: dataIn2 = 32'd0; 
32'd6052: dataIn2 = 32'd0; 
32'd6053: dataIn2 = 32'd0; 
32'd6054: dataIn2 = 32'd1; 
32'd6055: dataIn2 = 32'd0; 
32'd6056: dataIn2 = 32'd1; 
32'd6057: dataIn2 = 32'd1; 
32'd6058: dataIn2 = 32'd0; 
32'd6059: dataIn2 = 32'd1; 
32'd6060: dataIn2 = 32'd0; 
32'd6061: dataIn2 = 32'd1; 
32'd6062: dataIn2 = 32'd0; 
32'd6063: dataIn2 = 32'd1; 
32'd6064: dataIn2 = 32'd1; 
32'd6065: dataIn2 = 32'd1; 
32'd6066: dataIn2 = 32'd0; 
32'd6067: dataIn2 = 32'd0; 
32'd6068: dataIn2 = 32'd0; 
32'd6069: dataIn2 = 32'd0; 
32'd6070: dataIn2 = 32'd0; 
32'd6071: dataIn2 = 32'd1; 
32'd6072: dataIn2 = 32'd0; 
32'd6073: dataIn2 = 32'd1; 
32'd6074: dataIn2 = 32'd1; 
32'd6075: dataIn2 = 32'd1; 
32'd6076: dataIn2 = 32'd1; 
32'd6077: dataIn2 = 32'd1; 
32'd6078: dataIn2 = 32'd0; 
32'd6079: dataIn2 = 32'd1; 
32'd6080: dataIn2 = 32'd0; 
32'd6081: dataIn2 = 32'd1; 
32'd6082: dataIn2 = 32'd1; 
32'd6083: dataIn2 = 32'd1; 
32'd6084: dataIn2 = 32'd0; 
32'd6085: dataIn2 = 32'd0; 
32'd6086: dataIn2 = 32'd1; 
32'd6087: dataIn2 = 32'd0; 
32'd6088: dataIn2 = 32'd1; 
32'd6089: dataIn2 = 32'd1; 
32'd6090: dataIn2 = 32'd1; 
32'd6091: dataIn2 = 32'd0; 
32'd6092: dataIn2 = 32'd1; 
32'd6093: dataIn2 = 32'd0; 
32'd6094: dataIn2 = 32'd1; 
32'd6095: dataIn2 = 32'd0; 
32'd6096: dataIn2 = 32'd0; 
32'd6097: dataIn2 = 32'd0; 
32'd6098: dataIn2 = 32'd1; 
32'd6099: dataIn2 = 32'd0; 
32'd6100: dataIn2 = 32'd0; 
32'd6101: dataIn2 = 32'd1; 
32'd6102: dataIn2 = 32'd1; 
32'd6103: dataIn2 = 32'd0; 
32'd6104: dataIn2 = 32'd0; 
32'd6105: dataIn2 = 32'd0; 
32'd6106: dataIn2 = 32'd0; 
32'd6107: dataIn2 = 32'd0; 
32'd6108: dataIn2 = 32'd1; 
32'd6109: dataIn2 = 32'd0; 
32'd6110: dataIn2 = 32'd1; 
32'd6111: dataIn2 = 32'd0; 
32'd6112: dataIn2 = 32'd1; 
32'd6113: dataIn2 = 32'd0; 
32'd6114: dataIn2 = 32'd1; 
32'd6115: dataIn2 = 32'd0; 
32'd6116: dataIn2 = 32'd0; 
32'd6117: dataIn2 = 32'd0; 
32'd6118: dataIn2 = 32'd0; 
32'd6119: dataIn2 = 32'd1; 
32'd6120: dataIn2 = 32'd1; 
32'd6121: dataIn2 = 32'd1; 
32'd6122: dataIn2 = 32'd0; 
32'd6123: dataIn2 = 32'd1; 
32'd6124: dataIn2 = 32'd1; 
32'd6125: dataIn2 = 32'd1; 
32'd6126: dataIn2 = 32'd1; 
32'd6127: dataIn2 = 32'd1; 
32'd6128: dataIn2 = 32'd0; 
32'd6129: dataIn2 = 32'd0; 
32'd6130: dataIn2 = 32'd1; 
32'd6131: dataIn2 = 32'd0; 
32'd6132: dataIn2 = 32'd1; 
32'd6133: dataIn2 = 32'd0; 
32'd6134: dataIn2 = 32'd0; 
32'd6135: dataIn2 = 32'd1; 
32'd6136: dataIn2 = 32'd1; 
32'd6137: dataIn2 = 32'd0; 
32'd6138: dataIn2 = 32'd1; 
32'd6139: dataIn2 = 32'd1; 
32'd6140: dataIn2 = 32'd0; 
32'd6141: dataIn2 = 32'd1; 
32'd6142: dataIn2 = 32'd1; 
32'd6143: dataIn2 = 32'd0; 
32'd6144: dataIn2 = 32'd1; 
32'd6145: dataIn2 = 32'd0; 
32'd6146: dataIn2 = 32'd0; 
32'd6147: dataIn2 = 32'd0; 
32'd6148: dataIn2 = 32'd0; 
32'd6149: dataIn2 = 32'd0; 
32'd6150: dataIn2 = 32'd1; 
32'd6151: dataIn2 = 32'd1; 
32'd6152: dataIn2 = 32'd1; 
32'd6153: dataIn2 = 32'd0; 
32'd6154: dataIn2 = 32'd1; 
32'd6155: dataIn2 = 32'd1; 
32'd6156: dataIn2 = 32'd1; 
32'd6157: dataIn2 = 32'd0; 
32'd6158: dataIn2 = 32'd0; 
32'd6159: dataIn2 = 32'd0; 
32'd6160: dataIn2 = 32'd1; 
32'd6161: dataIn2 = 32'd0; 
32'd6162: dataIn2 = 32'd1; 
32'd6163: dataIn2 = 32'd0; 
32'd6164: dataIn2 = 32'd0; 
32'd6165: dataIn2 = 32'd0; 
32'd6166: dataIn2 = 32'd0; 
32'd6167: dataIn2 = 32'd0; 
32'd6168: dataIn2 = 32'd0; 
32'd6169: dataIn2 = 32'd0; 
32'd6170: dataIn2 = 32'd0; 
32'd6171: dataIn2 = 32'd1; 
32'd6172: dataIn2 = 32'd1; 
32'd6173: dataIn2 = 32'd1; 
32'd6174: dataIn2 = 32'd0; 
32'd6175: dataIn2 = 32'd1; 
32'd6176: dataIn2 = 32'd0; 
32'd6177: dataIn2 = 32'd0; 
32'd6178: dataIn2 = 32'd0; 
32'd6179: dataIn2 = 32'd1; 
32'd6180: dataIn2 = 32'd0; 
32'd6181: dataIn2 = 32'd1; 
32'd6182: dataIn2 = 32'd1; 
32'd6183: dataIn2 = 32'd0; 
32'd6184: dataIn2 = 32'd1; 
32'd6185: dataIn2 = 32'd1; 
32'd6186: dataIn2 = 32'd1; 
32'd6187: dataIn2 = 32'd1; 
32'd6188: dataIn2 = 32'd0; 
32'd6189: dataIn2 = 32'd1; 
32'd6190: dataIn2 = 32'd0; 
32'd6191: dataIn2 = 32'd1; 
32'd6192: dataIn2 = 32'd0; 
32'd6193: dataIn2 = 32'd0; 
32'd6194: dataIn2 = 32'd1; 
32'd6195: dataIn2 = 32'd1; 
32'd6196: dataIn2 = 32'd0; 
32'd6197: dataIn2 = 32'd1; 
32'd6198: dataIn2 = 32'd0; 
32'd6199: dataIn2 = 32'd0; 
32'd6200: dataIn2 = 32'd0; 
32'd6201: dataIn2 = 32'd0; 
32'd6202: dataIn2 = 32'd1; 
32'd6203: dataIn2 = 32'd1; 
32'd6204: dataIn2 = 32'd1; 
32'd6205: dataIn2 = 32'd1; 
32'd6206: dataIn2 = 32'd0; 
32'd6207: dataIn2 = 32'd1; 
32'd6208: dataIn2 = 32'd0; 
32'd6209: dataIn2 = 32'd1; 
32'd6210: dataIn2 = 32'd1; 
32'd6211: dataIn2 = 32'd0; 
32'd6212: dataIn2 = 32'd1; 
32'd6213: dataIn2 = 32'd1; 
32'd6214: dataIn2 = 32'd0; 
32'd6215: dataIn2 = 32'd0; 
32'd6216: dataIn2 = 32'd0; 
32'd6217: dataIn2 = 32'd0; 
32'd6218: dataIn2 = 32'd0; 
32'd6219: dataIn2 = 32'd1; 
32'd6220: dataIn2 = 32'd1; 
32'd6221: dataIn2 = 32'd0; 
32'd6222: dataIn2 = 32'd1; 
32'd6223: dataIn2 = 32'd1; 
32'd6224: dataIn2 = 32'd1; 
32'd6225: dataIn2 = 32'd0; 
32'd6226: dataIn2 = 32'd1; 
32'd6227: dataIn2 = 32'd1; 
32'd6228: dataIn2 = 32'd1; 
32'd6229: dataIn2 = 32'd1; 
32'd6230: dataIn2 = 32'd0; 
32'd6231: dataIn2 = 32'd0; 
32'd6232: dataIn2 = 32'd0; 
32'd6233: dataIn2 = 32'd0; 
32'd6234: dataIn2 = 32'd1; 
32'd6235: dataIn2 = 32'd0; 
32'd6236: dataIn2 = 32'd0; 
32'd6237: dataIn2 = 32'd0; 
32'd6238: dataIn2 = 32'd1; 
32'd6239: dataIn2 = 32'd0; 
32'd6240: dataIn2 = 32'd1; 
32'd6241: dataIn2 = 32'd1; 
32'd6242: dataIn2 = 32'd1; 
32'd6243: dataIn2 = 32'd1; 
32'd6244: dataIn2 = 32'd1; 
32'd6245: dataIn2 = 32'd0; 
32'd6246: dataIn2 = 32'd1; 
32'd6247: dataIn2 = 32'd0; 
32'd6248: dataIn2 = 32'd1; 
32'd6249: dataIn2 = 32'd1; 
32'd6250: dataIn2 = 32'd1; 
32'd6251: dataIn2 = 32'd1; 
32'd6252: dataIn2 = 32'd0; 
32'd6253: dataIn2 = 32'd1; 
32'd6254: dataIn2 = 32'd1; 
32'd6255: dataIn2 = 32'd0; 
32'd6256: dataIn2 = 32'd0; 
32'd6257: dataIn2 = 32'd1; 
32'd6258: dataIn2 = 32'd1; 
32'd6259: dataIn2 = 32'd0; 
32'd6260: dataIn2 = 32'd0; 
32'd6261: dataIn2 = 32'd1; 
32'd6262: dataIn2 = 32'd0; 
32'd6263: dataIn2 = 32'd1; 
32'd6264: dataIn2 = 32'd0; 
32'd6265: dataIn2 = 32'd0; 
32'd6266: dataIn2 = 32'd0; 
32'd6267: dataIn2 = 32'd1; 
32'd6268: dataIn2 = 32'd0; 
32'd6269: dataIn2 = 32'd1; 
32'd6270: dataIn2 = 32'd1; 
32'd6271: dataIn2 = 32'd1; 
32'd6272: dataIn2 = 32'd1; 
32'd6273: dataIn2 = 32'd1; 
32'd6274: dataIn2 = 32'd0; 
32'd6275: dataIn2 = 32'd1; 
32'd6276: dataIn2 = 32'd1; 
32'd6277: dataIn2 = 32'd1; 
32'd6278: dataIn2 = 32'd1; 
32'd6279: dataIn2 = 32'd0; 
32'd6280: dataIn2 = 32'd0; 
32'd6281: dataIn2 = 32'd1; 
32'd6282: dataIn2 = 32'd1; 
32'd6283: dataIn2 = 32'd1; 
32'd6284: dataIn2 = 32'd1; 
32'd6285: dataIn2 = 32'd1; 
32'd6286: dataIn2 = 32'd0; 
32'd6287: dataIn2 = 32'd1; 
32'd6288: dataIn2 = 32'd1; 
32'd6289: dataIn2 = 32'd0; 
32'd6290: dataIn2 = 32'd0; 
32'd6291: dataIn2 = 32'd0; 
32'd6292: dataIn2 = 32'd1; 
32'd6293: dataIn2 = 32'd1; 
32'd6294: dataIn2 = 32'd1; 
32'd6295: dataIn2 = 32'd0; 
32'd6296: dataIn2 = 32'd1; 
32'd6297: dataIn2 = 32'd0; 
32'd6298: dataIn2 = 32'd1; 
32'd6299: dataIn2 = 32'd0; 
32'd6300: dataIn2 = 32'd1; 
32'd6301: dataIn2 = 32'd1; 
32'd6302: dataIn2 = 32'd0; 
32'd6303: dataIn2 = 32'd0; 
32'd6304: dataIn2 = 32'd1; 
32'd6305: dataIn2 = 32'd0; 
32'd6306: dataIn2 = 32'd0; 
32'd6307: dataIn2 = 32'd0; 
32'd6308: dataIn2 = 32'd1; 
32'd6309: dataIn2 = 32'd0; 
32'd6310: dataIn2 = 32'd1; 
32'd6311: dataIn2 = 32'd0; 
32'd6312: dataIn2 = 32'd0; 
32'd6313: dataIn2 = 32'd1; 
32'd6314: dataIn2 = 32'd0; 
32'd6315: dataIn2 = 32'd0; 
32'd6316: dataIn2 = 32'd0; 
32'd6317: dataIn2 = 32'd1; 
32'd6318: dataIn2 = 32'd1; 
32'd6319: dataIn2 = 32'd1; 
32'd6320: dataIn2 = 32'd0; 
32'd6321: dataIn2 = 32'd1; 
32'd6322: dataIn2 = 32'd1; 
32'd6323: dataIn2 = 32'd1; 
32'd6324: dataIn2 = 32'd0; 
32'd6325: dataIn2 = 32'd0; 
32'd6326: dataIn2 = 32'd0; 
32'd6327: dataIn2 = 32'd0; 
32'd6328: dataIn2 = 32'd0; 
32'd6329: dataIn2 = 32'd0; 
32'd6330: dataIn2 = 32'd1; 
32'd6331: dataIn2 = 32'd0; 
32'd6332: dataIn2 = 32'd0; 
32'd6333: dataIn2 = 32'd0; 
32'd6334: dataIn2 = 32'd0; 
32'd6335: dataIn2 = 32'd1; 
32'd6336: dataIn2 = 32'd0; 
32'd6337: dataIn2 = 32'd1; 
32'd6338: dataIn2 = 32'd0; 
32'd6339: dataIn2 = 32'd1; 
32'd6340: dataIn2 = 32'd0; 
32'd6341: dataIn2 = 32'd1; 
32'd6342: dataIn2 = 32'd0; 
32'd6343: dataIn2 = 32'd1; 
32'd6344: dataIn2 = 32'd1; 
32'd6345: dataIn2 = 32'd0; 
32'd6346: dataIn2 = 32'd1; 
32'd6347: dataIn2 = 32'd0; 
32'd6348: dataIn2 = 32'd0; 
32'd6349: dataIn2 = 32'd1; 
32'd6350: dataIn2 = 32'd1; 
32'd6351: dataIn2 = 32'd1; 
32'd6352: dataIn2 = 32'd0; 
32'd6353: dataIn2 = 32'd1; 
32'd6354: dataIn2 = 32'd0; 
32'd6355: dataIn2 = 32'd1; 
32'd6356: dataIn2 = 32'd1; 
32'd6357: dataIn2 = 32'd0; 
32'd6358: dataIn2 = 32'd1; 
32'd6359: dataIn2 = 32'd0; 
32'd6360: dataIn2 = 32'd1; 
32'd6361: dataIn2 = 32'd0; 
32'd6362: dataIn2 = 32'd0; 
32'd6363: dataIn2 = 32'd0; 
32'd6364: dataIn2 = 32'd0; 
32'd6365: dataIn2 = 32'd1; 
32'd6366: dataIn2 = 32'd1; 
32'd6367: dataIn2 = 32'd0; 
32'd6368: dataIn2 = 32'd0; 
32'd6369: dataIn2 = 32'd0; 
32'd6370: dataIn2 = 32'd1; 
32'd6371: dataIn2 = 32'd0; 
32'd6372: dataIn2 = 32'd0; 
32'd6373: dataIn2 = 32'd1; 
32'd6374: dataIn2 = 32'd0; 
32'd6375: dataIn2 = 32'd1; 
32'd6376: dataIn2 = 32'd0; 
32'd6377: dataIn2 = 32'd0; 
32'd6378: dataIn2 = 32'd1; 
32'd6379: dataIn2 = 32'd1; 
32'd6380: dataIn2 = 32'd1; 
32'd6381: dataIn2 = 32'd1; 
32'd6382: dataIn2 = 32'd0; 
32'd6383: dataIn2 = 32'd1; 
32'd6384: dataIn2 = 32'd1; 
32'd6385: dataIn2 = 32'd0; 
32'd6386: dataIn2 = 32'd0; 
32'd6387: dataIn2 = 32'd1; 
32'd6388: dataIn2 = 32'd1; 
32'd6389: dataIn2 = 32'd1; 
32'd6390: dataIn2 = 32'd0; 
32'd6391: dataIn2 = 32'd1; 
32'd6392: dataIn2 = 32'd1; 
32'd6393: dataIn2 = 32'd0; 
32'd6394: dataIn2 = 32'd0; 
32'd6395: dataIn2 = 32'd0; 
32'd6396: dataIn2 = 32'd0; 
32'd6397: dataIn2 = 32'd0; 
32'd6398: dataIn2 = 32'd1; 
32'd6399: dataIn2 = 32'd1; 
32'd6400: dataIn2 = 32'd0; 
32'd6401: dataIn2 = 32'd1; 
32'd6402: dataIn2 = 32'd0; 
32'd6403: dataIn2 = 32'd0; 
32'd6404: dataIn2 = 32'd1; 
32'd6405: dataIn2 = 32'd1; 
32'd6406: dataIn2 = 32'd0; 
32'd6407: dataIn2 = 32'd1; 
32'd6408: dataIn2 = 32'd1; 
32'd6409: dataIn2 = 32'd0; 
32'd6410: dataIn2 = 32'd1; 
32'd6411: dataIn2 = 32'd0; 
32'd6412: dataIn2 = 32'd1; 
32'd6413: dataIn2 = 32'd0; 
32'd6414: dataIn2 = 32'd1; 
32'd6415: dataIn2 = 32'd0; 
32'd6416: dataIn2 = 32'd0; 
32'd6417: dataIn2 = 32'd1; 
32'd6418: dataIn2 = 32'd1; 
32'd6419: dataIn2 = 32'd0; 
32'd6420: dataIn2 = 32'd1; 
32'd6421: dataIn2 = 32'd0; 
32'd6422: dataIn2 = 32'd1; 
32'd6423: dataIn2 = 32'd0; 
32'd6424: dataIn2 = 32'd0; 
32'd6425: dataIn2 = 32'd1; 
32'd6426: dataIn2 = 32'd0; 
32'd6427: dataIn2 = 32'd0; 
32'd6428: dataIn2 = 32'd0; 
32'd6429: dataIn2 = 32'd0; 
32'd6430: dataIn2 = 32'd0; 
32'd6431: dataIn2 = 32'd1; 
32'd6432: dataIn2 = 32'd1; 
32'd6433: dataIn2 = 32'd0; 
32'd6434: dataIn2 = 32'd0; 
32'd6435: dataIn2 = 32'd0; 
32'd6436: dataIn2 = 32'd0; 
32'd6437: dataIn2 = 32'd0; 
32'd6438: dataIn2 = 32'd0; 
32'd6439: dataIn2 = 32'd1; 
32'd6440: dataIn2 = 32'd0; 
32'd6441: dataIn2 = 32'd1; 
32'd6442: dataIn2 = 32'd1; 
32'd6443: dataIn2 = 32'd1; 
32'd6444: dataIn2 = 32'd1; 
32'd6445: dataIn2 = 32'd0; 
32'd6446: dataIn2 = 32'd1; 
32'd6447: dataIn2 = 32'd1; 
32'd6448: dataIn2 = 32'd0; 
32'd6449: dataIn2 = 32'd1; 
32'd6450: dataIn2 = 32'd1; 
32'd6451: dataIn2 = 32'd1; 
32'd6452: dataIn2 = 32'd0; 
32'd6453: dataIn2 = 32'd1; 
32'd6454: dataIn2 = 32'd0; 
32'd6455: dataIn2 = 32'd1; 
32'd6456: dataIn2 = 32'd1; 
32'd6457: dataIn2 = 32'd0; 
32'd6458: dataIn2 = 32'd1; 
32'd6459: dataIn2 = 32'd1; 
32'd6460: dataIn2 = 32'd0; 
32'd6461: dataIn2 = 32'd1; 
32'd6462: dataIn2 = 32'd0; 
32'd6463: dataIn2 = 32'd0; 
32'd6464: dataIn2 = 32'd0; 
32'd6465: dataIn2 = 32'd1; 
32'd6466: dataIn2 = 32'd1; 
32'd6467: dataIn2 = 32'd0; 
32'd6468: dataIn2 = 32'd0; 
32'd6469: dataIn2 = 32'd0; 
32'd6470: dataIn2 = 32'd1; 
32'd6471: dataIn2 = 32'd0; 
32'd6472: dataIn2 = 32'd1; 
32'd6473: dataIn2 = 32'd0; 
32'd6474: dataIn2 = 32'd1; 
32'd6475: dataIn2 = 32'd1; 
32'd6476: dataIn2 = 32'd0; 
32'd6477: dataIn2 = 32'd1; 
32'd6478: dataIn2 = 32'd1; 
32'd6479: dataIn2 = 32'd1; 
32'd6480: dataIn2 = 32'd0; 
32'd6481: dataIn2 = 32'd0; 
32'd6482: dataIn2 = 32'd0; 
32'd6483: dataIn2 = 32'd1; 
32'd6484: dataIn2 = 32'd1; 
32'd6485: dataIn2 = 32'd1; 
32'd6486: dataIn2 = 32'd1; 
32'd6487: dataIn2 = 32'd1; 
32'd6488: dataIn2 = 32'd0; 
32'd6489: dataIn2 = 32'd1; 
32'd6490: dataIn2 = 32'd0; 
32'd6491: dataIn2 = 32'd1; 
32'd6492: dataIn2 = 32'd1; 
32'd6493: dataIn2 = 32'd1; 
32'd6494: dataIn2 = 32'd0; 
32'd6495: dataIn2 = 32'd1; 
32'd6496: dataIn2 = 32'd0; 
32'd6497: dataIn2 = 32'd1; 
32'd6498: dataIn2 = 32'd0; 
32'd6499: dataIn2 = 32'd1; 
32'd6500: dataIn2 = 32'd0; 
32'd6501: dataIn2 = 32'd1; 
32'd6502: dataIn2 = 32'd1; 
32'd6503: dataIn2 = 32'd0; 
32'd6504: dataIn2 = 32'd0; 
32'd6505: dataIn2 = 32'd0; 
32'd6506: dataIn2 = 32'd0; 
32'd6507: dataIn2 = 32'd0; 
32'd6508: dataIn2 = 32'd0; 
32'd6509: dataIn2 = 32'd0; 
32'd6510: dataIn2 = 32'd1; 
32'd6511: dataIn2 = 32'd0; 
32'd6512: dataIn2 = 32'd1; 
32'd6513: dataIn2 = 32'd0; 
32'd6514: dataIn2 = 32'd1; 
32'd6515: dataIn2 = 32'd0; 
32'd6516: dataIn2 = 32'd0; 
32'd6517: dataIn2 = 32'd1; 
32'd6518: dataIn2 = 32'd0; 
32'd6519: dataIn2 = 32'd0; 
32'd6520: dataIn2 = 32'd0; 
32'd6521: dataIn2 = 32'd0; 
32'd6522: dataIn2 = 32'd0; 
32'd6523: dataIn2 = 32'd1; 
32'd6524: dataIn2 = 32'd0; 
32'd6525: dataIn2 = 32'd0; 
32'd6526: dataIn2 = 32'd0; 
32'd6527: dataIn2 = 32'd0; 
32'd6528: dataIn2 = 32'd0; 
32'd6529: dataIn2 = 32'd1; 
32'd6530: dataIn2 = 32'd0; 
32'd6531: dataIn2 = 32'd0; 
32'd6532: dataIn2 = 32'd1; 
32'd6533: dataIn2 = 32'd1; 
32'd6534: dataIn2 = 32'd1; 
32'd6535: dataIn2 = 32'd1; 
32'd6536: dataIn2 = 32'd0; 
32'd6537: dataIn2 = 32'd1; 
32'd6538: dataIn2 = 32'd0; 
32'd6539: dataIn2 = 32'd1; 
32'd6540: dataIn2 = 32'd1; 
32'd6541: dataIn2 = 32'd0; 
32'd6542: dataIn2 = 32'd0; 
32'd6543: dataIn2 = 32'd0; 
32'd6544: dataIn2 = 32'd0; 
32'd6545: dataIn2 = 32'd0; 
32'd6546: dataIn2 = 32'd1; 
32'd6547: dataIn2 = 32'd0; 
32'd6548: dataIn2 = 32'd1; 
32'd6549: dataIn2 = 32'd0; 
32'd6550: dataIn2 = 32'd1; 
32'd6551: dataIn2 = 32'd0; 
32'd6552: dataIn2 = 32'd1; 
32'd6553: dataIn2 = 32'd1; 
32'd6554: dataIn2 = 32'd0; 
32'd6555: dataIn2 = 32'd1; 
32'd6556: dataIn2 = 32'd1; 
32'd6557: dataIn2 = 32'd0; 
32'd6558: dataIn2 = 32'd1; 
32'd6559: dataIn2 = 32'd1; 
32'd6560: dataIn2 = 32'd0; 
32'd6561: dataIn2 = 32'd1; 
32'd6562: dataIn2 = 32'd1; 
32'd6563: dataIn2 = 32'd1; 
32'd6564: dataIn2 = 32'd0; 
32'd6565: dataIn2 = 32'd1; 
32'd6566: dataIn2 = 32'd0; 
32'd6567: dataIn2 = 32'd0; 
32'd6568: dataIn2 = 32'd1; 
32'd6569: dataIn2 = 32'd0; 
32'd6570: dataIn2 = 32'd0; 
32'd6571: dataIn2 = 32'd1; 
32'd6572: dataIn2 = 32'd0; 
32'd6573: dataIn2 = 32'd0; 
32'd6574: dataIn2 = 32'd0; 
32'd6575: dataIn2 = 32'd1; 
32'd6576: dataIn2 = 32'd1; 
32'd6577: dataIn2 = 32'd0; 
32'd6578: dataIn2 = 32'd1; 
32'd6579: dataIn2 = 32'd0; 
32'd6580: dataIn2 = 32'd0; 
32'd6581: dataIn2 = 32'd1; 
32'd6582: dataIn2 = 32'd0; 
32'd6583: dataIn2 = 32'd0; 
32'd6584: dataIn2 = 32'd0; 
32'd6585: dataIn2 = 32'd0; 
32'd6586: dataIn2 = 32'd0; 
32'd6587: dataIn2 = 32'd1; 
32'd6588: dataIn2 = 32'd0; 
32'd6589: dataIn2 = 32'd1; 
32'd6590: dataIn2 = 32'd0; 
32'd6591: dataIn2 = 32'd1; 
32'd6592: dataIn2 = 32'd0; 
32'd6593: dataIn2 = 32'd0; 
32'd6594: dataIn2 = 32'd0; 
32'd6595: dataIn2 = 32'd0; 
32'd6596: dataIn2 = 32'd0; 
32'd6597: dataIn2 = 32'd0; 
32'd6598: dataIn2 = 32'd0; 
32'd6599: dataIn2 = 32'd0; 
32'd6600: dataIn2 = 32'd0; 
32'd6601: dataIn2 = 32'd1; 
32'd6602: dataIn2 = 32'd1; 
32'd6603: dataIn2 = 32'd1; 
32'd6604: dataIn2 = 32'd0; 
32'd6605: dataIn2 = 32'd1; 
32'd6606: dataIn2 = 32'd0; 
32'd6607: dataIn2 = 32'd1; 
32'd6608: dataIn2 = 32'd1; 
32'd6609: dataIn2 = 32'd1; 
32'd6610: dataIn2 = 32'd0; 
32'd6611: dataIn2 = 32'd0; 
32'd6612: dataIn2 = 32'd1; 
32'd6613: dataIn2 = 32'd1; 
32'd6614: dataIn2 = 32'd1; 
32'd6615: dataIn2 = 32'd0; 
32'd6616: dataIn2 = 32'd0; 
32'd6617: dataIn2 = 32'd1; 
32'd6618: dataIn2 = 32'd1; 
32'd6619: dataIn2 = 32'd1; 
32'd6620: dataIn2 = 32'd0; 
32'd6621: dataIn2 = 32'd0; 
32'd6622: dataIn2 = 32'd0; 
32'd6623: dataIn2 = 32'd0; 
32'd6624: dataIn2 = 32'd1; 
32'd6625: dataIn2 = 32'd1; 
32'd6626: dataIn2 = 32'd0; 
32'd6627: dataIn2 = 32'd1; 
32'd6628: dataIn2 = 32'd1; 
32'd6629: dataIn2 = 32'd0; 
32'd6630: dataIn2 = 32'd0; 
32'd6631: dataIn2 = 32'd1; 
32'd6632: dataIn2 = 32'd0; 
32'd6633: dataIn2 = 32'd0; 
32'd6634: dataIn2 = 32'd0; 
32'd6635: dataIn2 = 32'd0; 
32'd6636: dataIn2 = 32'd1; 
32'd6637: dataIn2 = 32'd1; 
32'd6638: dataIn2 = 32'd1; 
32'd6639: dataIn2 = 32'd1; 
32'd6640: dataIn2 = 32'd1; 
32'd6641: dataIn2 = 32'd0; 
32'd6642: dataIn2 = 32'd1; 
32'd6643: dataIn2 = 32'd0; 
32'd6644: dataIn2 = 32'd0; 
32'd6645: dataIn2 = 32'd0; 
32'd6646: dataIn2 = 32'd1; 
32'd6647: dataIn2 = 32'd0; 
32'd6648: dataIn2 = 32'd0; 
32'd6649: dataIn2 = 32'd0; 
32'd6650: dataIn2 = 32'd1; 
32'd6651: dataIn2 = 32'd1; 
32'd6652: dataIn2 = 32'd1; 
32'd6653: dataIn2 = 32'd0; 
32'd6654: dataIn2 = 32'd0; 
32'd6655: dataIn2 = 32'd0; 
32'd6656: dataIn2 = 32'd0; 
32'd6657: dataIn2 = 32'd1; 
32'd6658: dataIn2 = 32'd1; 
32'd6659: dataIn2 = 32'd1; 
32'd6660: dataIn2 = 32'd0; 
32'd6661: dataIn2 = 32'd0; 
32'd6662: dataIn2 = 32'd0; 
32'd6663: dataIn2 = 32'd0; 
32'd6664: dataIn2 = 32'd0; 
32'd6665: dataIn2 = 32'd0; 
32'd6666: dataIn2 = 32'd0; 
32'd6667: dataIn2 = 32'd1; 
32'd6668: dataIn2 = 32'd1; 
32'd6669: dataIn2 = 32'd0; 
32'd6670: dataIn2 = 32'd1; 
32'd6671: dataIn2 = 32'd1; 
32'd6672: dataIn2 = 32'd0; 
32'd6673: dataIn2 = 32'd0; 
32'd6674: dataIn2 = 32'd1; 
32'd6675: dataIn2 = 32'd1; 
32'd6676: dataIn2 = 32'd1; 
32'd6677: dataIn2 = 32'd1; 
32'd6678: dataIn2 = 32'd0; 
32'd6679: dataIn2 = 32'd1; 
32'd6680: dataIn2 = 32'd1; 
32'd6681: dataIn2 = 32'd1; 
32'd6682: dataIn2 = 32'd1; 
32'd6683: dataIn2 = 32'd0; 
32'd6684: dataIn2 = 32'd0; 
32'd6685: dataIn2 = 32'd1; 
32'd6686: dataIn2 = 32'd1; 
32'd6687: dataIn2 = 32'd0; 
32'd6688: dataIn2 = 32'd0; 
32'd6689: dataIn2 = 32'd1; 
32'd6690: dataIn2 = 32'd0; 
32'd6691: dataIn2 = 32'd0; 
32'd6692: dataIn2 = 32'd0; 
32'd6693: dataIn2 = 32'd1; 
32'd6694: dataIn2 = 32'd1; 
32'd6695: dataIn2 = 32'd0; 
32'd6696: dataIn2 = 32'd1; 
32'd6697: dataIn2 = 32'd1; 
32'd6698: dataIn2 = 32'd0; 
32'd6699: dataIn2 = 32'd1; 
32'd6700: dataIn2 = 32'd0; 
32'd6701: dataIn2 = 32'd1; 
32'd6702: dataIn2 = 32'd1; 
32'd6703: dataIn2 = 32'd1; 
32'd6704: dataIn2 = 32'd1; 
32'd6705: dataIn2 = 32'd0; 
32'd6706: dataIn2 = 32'd0; 
32'd6707: dataIn2 = 32'd0; 
32'd6708: dataIn2 = 32'd1; 
32'd6709: dataIn2 = 32'd0; 
32'd6710: dataIn2 = 32'd0; 
32'd6711: dataIn2 = 32'd0; 
32'd6712: dataIn2 = 32'd1; 
32'd6713: dataIn2 = 32'd0; 
32'd6714: dataIn2 = 32'd1; 
32'd6715: dataIn2 = 32'd1; 
32'd6716: dataIn2 = 32'd1; 
32'd6717: dataIn2 = 32'd1; 
32'd6718: dataIn2 = 32'd0; 
32'd6719: dataIn2 = 32'd0; 
32'd6720: dataIn2 = 32'd1; 
32'd6721: dataIn2 = 32'd0; 
32'd6722: dataIn2 = 32'd1; 
32'd6723: dataIn2 = 32'd1; 
32'd6724: dataIn2 = 32'd1; 
32'd6725: dataIn2 = 32'd1; 
32'd6726: dataIn2 = 32'd0; 
32'd6727: dataIn2 = 32'd0; 
32'd6728: dataIn2 = 32'd0; 
32'd6729: dataIn2 = 32'd1; 
32'd6730: dataIn2 = 32'd0; 
32'd6731: dataIn2 = 32'd0; 
32'd6732: dataIn2 = 32'd0; 
32'd6733: dataIn2 = 32'd1; 
32'd6734: dataIn2 = 32'd0; 
32'd6735: dataIn2 = 32'd1; 
32'd6736: dataIn2 = 32'd1; 
32'd6737: dataIn2 = 32'd0; 
32'd6738: dataIn2 = 32'd1; 
32'd6739: dataIn2 = 32'd0; 
32'd6740: dataIn2 = 32'd0; 
32'd6741: dataIn2 = 32'd0; 
32'd6742: dataIn2 = 32'd0; 
32'd6743: dataIn2 = 32'd1; 
32'd6744: dataIn2 = 32'd1; 
32'd6745: dataIn2 = 32'd1; 
32'd6746: dataIn2 = 32'd0; 
32'd6747: dataIn2 = 32'd0; 
32'd6748: dataIn2 = 32'd1; 
32'd6749: dataIn2 = 32'd0; 
32'd6750: dataIn2 = 32'd1; 
32'd6751: dataIn2 = 32'd1; 
32'd6752: dataIn2 = 32'd0; 
32'd6753: dataIn2 = 32'd1; 
32'd6754: dataIn2 = 32'd1; 
32'd6755: dataIn2 = 32'd1; 
32'd6756: dataIn2 = 32'd1; 
32'd6757: dataIn2 = 32'd0; 
32'd6758: dataIn2 = 32'd1; 
32'd6759: dataIn2 = 32'd1; 
32'd6760: dataIn2 = 32'd0; 
32'd6761: dataIn2 = 32'd1; 
32'd6762: dataIn2 = 32'd0; 
32'd6763: dataIn2 = 32'd1; 
32'd6764: dataIn2 = 32'd1; 
32'd6765: dataIn2 = 32'd0; 
32'd6766: dataIn2 = 32'd0; 
32'd6767: dataIn2 = 32'd0; 
32'd6768: dataIn2 = 32'd1; 
32'd6769: dataIn2 = 32'd1; 
32'd6770: dataIn2 = 32'd0; 
32'd6771: dataIn2 = 32'd0; 
32'd6772: dataIn2 = 32'd1; 
32'd6773: dataIn2 = 32'd1; 
32'd6774: dataIn2 = 32'd0; 
32'd6775: dataIn2 = 32'd0; 
32'd6776: dataIn2 = 32'd1; 
32'd6777: dataIn2 = 32'd1; 
32'd6778: dataIn2 = 32'd0; 
32'd6779: dataIn2 = 32'd1; 
32'd6780: dataIn2 = 32'd1; 
32'd6781: dataIn2 = 32'd1; 
32'd6782: dataIn2 = 32'd1; 
32'd6783: dataIn2 = 32'd1; 
32'd6784: dataIn2 = 32'd1; 
32'd6785: dataIn2 = 32'd1; 
32'd6786: dataIn2 = 32'd0; 
32'd6787: dataIn2 = 32'd1; 
32'd6788: dataIn2 = 32'd0; 
32'd6789: dataIn2 = 32'd1; 
32'd6790: dataIn2 = 32'd0; 
32'd6791: dataIn2 = 32'd1; 
32'd6792: dataIn2 = 32'd1; 
32'd6793: dataIn2 = 32'd0; 
32'd6794: dataIn2 = 32'd1; 
32'd6795: dataIn2 = 32'd0; 
32'd6796: dataIn2 = 32'd1; 
32'd6797: dataIn2 = 32'd0; 
32'd6798: dataIn2 = 32'd1; 
32'd6799: dataIn2 = 32'd0; 
32'd6800: dataIn2 = 32'd1; 
32'd6801: dataIn2 = 32'd1; 
32'd6802: dataIn2 = 32'd1; 
32'd6803: dataIn2 = 32'd0; 
32'd6804: dataIn2 = 32'd1; 
32'd6805: dataIn2 = 32'd1; 
32'd6806: dataIn2 = 32'd1; 
32'd6807: dataIn2 = 32'd1; 
32'd6808: dataIn2 = 32'd0; 
32'd6809: dataIn2 = 32'd0; 
32'd6810: dataIn2 = 32'd1; 
32'd6811: dataIn2 = 32'd0; 
32'd6812: dataIn2 = 32'd0; 
32'd6813: dataIn2 = 32'd1; 
32'd6814: dataIn2 = 32'd1; 
32'd6815: dataIn2 = 32'd1; 
32'd6816: dataIn2 = 32'd1; 
32'd6817: dataIn2 = 32'd0; 
32'd6818: dataIn2 = 32'd1; 
32'd6819: dataIn2 = 32'd1; 
32'd6820: dataIn2 = 32'd0; 
32'd6821: dataIn2 = 32'd0; 
32'd6822: dataIn2 = 32'd0; 
32'd6823: dataIn2 = 32'd0; 
32'd6824: dataIn2 = 32'd0; 
32'd6825: dataIn2 = 32'd1; 
32'd6826: dataIn2 = 32'd1; 
32'd6827: dataIn2 = 32'd0; 
32'd6828: dataIn2 = 32'd0; 
32'd6829: dataIn2 = 32'd1; 
32'd6830: dataIn2 = 32'd1; 
32'd6831: dataIn2 = 32'd1; 
32'd6832: dataIn2 = 32'd1; 
32'd6833: dataIn2 = 32'd1; 
32'd6834: dataIn2 = 32'd1; 
32'd6835: dataIn2 = 32'd0; 
32'd6836: dataIn2 = 32'd0; 
32'd6837: dataIn2 = 32'd0; 
32'd6838: dataIn2 = 32'd1; 
32'd6839: dataIn2 = 32'd0; 
32'd6840: dataIn2 = 32'd0; 
32'd6841: dataIn2 = 32'd0; 
32'd6842: dataIn2 = 32'd0; 
32'd6843: dataIn2 = 32'd0; 
32'd6844: dataIn2 = 32'd1; 
32'd6845: dataIn2 = 32'd0; 
32'd6846: dataIn2 = 32'd1; 
32'd6847: dataIn2 = 32'd0; 
32'd6848: dataIn2 = 32'd1; 
32'd6849: dataIn2 = 32'd0; 
32'd6850: dataIn2 = 32'd0; 
32'd6851: dataIn2 = 32'd0; 
32'd6852: dataIn2 = 32'd0; 
32'd6853: dataIn2 = 32'd1; 
32'd6854: dataIn2 = 32'd1; 
32'd6855: dataIn2 = 32'd0; 
32'd6856: dataIn2 = 32'd1; 
32'd6857: dataIn2 = 32'd0; 
32'd6858: dataIn2 = 32'd1; 
32'd6859: dataIn2 = 32'd0; 
32'd6860: dataIn2 = 32'd0; 
32'd6861: dataIn2 = 32'd0; 
32'd6862: dataIn2 = 32'd1; 
32'd6863: dataIn2 = 32'd1; 
32'd6864: dataIn2 = 32'd1; 
32'd6865: dataIn2 = 32'd0; 
32'd6866: dataIn2 = 32'd0; 
32'd6867: dataIn2 = 32'd0; 
32'd6868: dataIn2 = 32'd0; 
32'd6869: dataIn2 = 32'd0; 
32'd6870: dataIn2 = 32'd0; 
32'd6871: dataIn2 = 32'd0; 
32'd6872: dataIn2 = 32'd1; 
32'd6873: dataIn2 = 32'd1; 
32'd6874: dataIn2 = 32'd0; 
32'd6875: dataIn2 = 32'd1; 
32'd6876: dataIn2 = 32'd1; 
32'd6877: dataIn2 = 32'd1; 
32'd6878: dataIn2 = 32'd0; 
32'd6879: dataIn2 = 32'd1; 
32'd6880: dataIn2 = 32'd0; 
32'd6881: dataIn2 = 32'd1; 
32'd6882: dataIn2 = 32'd1; 
32'd6883: dataIn2 = 32'd1; 
32'd6884: dataIn2 = 32'd1; 
32'd6885: dataIn2 = 32'd0; 
32'd6886: dataIn2 = 32'd0; 
32'd6887: dataIn2 = 32'd0; 
32'd6888: dataIn2 = 32'd1; 
32'd6889: dataIn2 = 32'd1; 
32'd6890: dataIn2 = 32'd0; 
32'd6891: dataIn2 = 32'd1; 
32'd6892: dataIn2 = 32'd0; 
32'd6893: dataIn2 = 32'd0; 
32'd6894: dataIn2 = 32'd0; 
32'd6895: dataIn2 = 32'd1; 
32'd6896: dataIn2 = 32'd0; 
32'd6897: dataIn2 = 32'd0; 
32'd6898: dataIn2 = 32'd1; 
32'd6899: dataIn2 = 32'd1; 
32'd6900: dataIn2 = 32'd0; 
32'd6901: dataIn2 = 32'd1; 
32'd6902: dataIn2 = 32'd1; 
32'd6903: dataIn2 = 32'd0; 
32'd6904: dataIn2 = 32'd0; 
32'd6905: dataIn2 = 32'd1; 
32'd6906: dataIn2 = 32'd0; 
32'd6907: dataIn2 = 32'd1; 
32'd6908: dataIn2 = 32'd0; 
32'd6909: dataIn2 = 32'd1; 
32'd6910: dataIn2 = 32'd1; 
32'd6911: dataIn2 = 32'd0; 
32'd6912: dataIn2 = 32'd0; 
32'd6913: dataIn2 = 32'd0; 
32'd6914: dataIn2 = 32'd0; 
32'd6915: dataIn2 = 32'd1; 
32'd6916: dataIn2 = 32'd0; 
32'd6917: dataIn2 = 32'd0; 
32'd6918: dataIn2 = 32'd0; 
32'd6919: dataIn2 = 32'd1; 
32'd6920: dataIn2 = 32'd0; 
32'd6921: dataIn2 = 32'd0; 
32'd6922: dataIn2 = 32'd0; 
32'd6923: dataIn2 = 32'd0; 
32'd6924: dataIn2 = 32'd0; 
32'd6925: dataIn2 = 32'd1; 
32'd6926: dataIn2 = 32'd0; 
32'd6927: dataIn2 = 32'd1; 
32'd6928: dataIn2 = 32'd0; 
32'd6929: dataIn2 = 32'd1; 
32'd6930: dataIn2 = 32'd1; 
32'd6931: dataIn2 = 32'd1; 
32'd6932: dataIn2 = 32'd0; 
32'd6933: dataIn2 = 32'd0; 
32'd6934: dataIn2 = 32'd1; 
32'd6935: dataIn2 = 32'd0; 
32'd6936: dataIn2 = 32'd0; 
32'd6937: dataIn2 = 32'd1; 
32'd6938: dataIn2 = 32'd0; 
32'd6939: dataIn2 = 32'd1; 
32'd6940: dataIn2 = 32'd0; 
32'd6941: dataIn2 = 32'd1; 
32'd6942: dataIn2 = 32'd1; 
32'd6943: dataIn2 = 32'd1; 
32'd6944: dataIn2 = 32'd1; 
32'd6945: dataIn2 = 32'd0; 
32'd6946: dataIn2 = 32'd0; 
32'd6947: dataIn2 = 32'd1; 
32'd6948: dataIn2 = 32'd1; 
32'd6949: dataIn2 = 32'd0; 
32'd6950: dataIn2 = 32'd0; 
32'd6951: dataIn2 = 32'd1; 
32'd6952: dataIn2 = 32'd0; 
32'd6953: dataIn2 = 32'd1; 
32'd6954: dataIn2 = 32'd1; 
32'd6955: dataIn2 = 32'd1; 
32'd6956: dataIn2 = 32'd0; 
32'd6957: dataIn2 = 32'd0; 
32'd6958: dataIn2 = 32'd0; 
32'd6959: dataIn2 = 32'd0; 
32'd6960: dataIn2 = 32'd1; 
32'd6961: dataIn2 = 32'd0; 
32'd6962: dataIn2 = 32'd0; 
32'd6963: dataIn2 = 32'd1; 
32'd6964: dataIn2 = 32'd1; 
32'd6965: dataIn2 = 32'd0; 
32'd6966: dataIn2 = 32'd1; 
32'd6967: dataIn2 = 32'd0; 
32'd6968: dataIn2 = 32'd0; 
32'd6969: dataIn2 = 32'd0; 
32'd6970: dataIn2 = 32'd1; 
32'd6971: dataIn2 = 32'd0; 
32'd6972: dataIn2 = 32'd0; 
32'd6973: dataIn2 = 32'd0; 
32'd6974: dataIn2 = 32'd0; 
32'd6975: dataIn2 = 32'd1; 
32'd6976: dataIn2 = 32'd0; 
32'd6977: dataIn2 = 32'd1; 
32'd6978: dataIn2 = 32'd0; 
32'd6979: dataIn2 = 32'd0; 
32'd6980: dataIn2 = 32'd0; 
32'd6981: dataIn2 = 32'd0; 
32'd6982: dataIn2 = 32'd1; 
32'd6983: dataIn2 = 32'd1; 
32'd6984: dataIn2 = 32'd1; 
32'd6985: dataIn2 = 32'd0; 
32'd6986: dataIn2 = 32'd1; 
32'd6987: dataIn2 = 32'd0; 
32'd6988: dataIn2 = 32'd0; 
32'd6989: dataIn2 = 32'd0; 
32'd6990: dataIn2 = 32'd1; 
32'd6991: dataIn2 = 32'd0; 
32'd6992: dataIn2 = 32'd0; 
32'd6993: dataIn2 = 32'd1; 
32'd6994: dataIn2 = 32'd1; 
32'd6995: dataIn2 = 32'd0; 
32'd6996: dataIn2 = 32'd1; 
32'd6997: dataIn2 = 32'd1; 
32'd6998: dataIn2 = 32'd1; 
32'd6999: dataIn2 = 32'd0; 
32'd7000: dataIn2 = 32'd0; 
32'd7001: dataIn2 = 32'd0; 
32'd7002: dataIn2 = 32'd0; 
32'd7003: dataIn2 = 32'd0; 
32'd7004: dataIn2 = 32'd0; 
32'd7005: dataIn2 = 32'd1; 
32'd7006: dataIn2 = 32'd1; 
32'd7007: dataIn2 = 32'd1; 
32'd7008: dataIn2 = 32'd0; 
32'd7009: dataIn2 = 32'd0; 
32'd7010: dataIn2 = 32'd1; 
32'd7011: dataIn2 = 32'd0; 
32'd7012: dataIn2 = 32'd1; 
32'd7013: dataIn2 = 32'd1; 
32'd7014: dataIn2 = 32'd0; 
32'd7015: dataIn2 = 32'd0; 
32'd7016: dataIn2 = 32'd1; 
32'd7017: dataIn2 = 32'd0; 
32'd7018: dataIn2 = 32'd1; 
32'd7019: dataIn2 = 32'd0; 
32'd7020: dataIn2 = 32'd0; 
32'd7021: dataIn2 = 32'd1; 
32'd7022: dataIn2 = 32'd1; 
32'd7023: dataIn2 = 32'd1; 
32'd7024: dataIn2 = 32'd0; 
32'd7025: dataIn2 = 32'd0; 
32'd7026: dataIn2 = 32'd0; 
32'd7027: dataIn2 = 32'd0; 
32'd7028: dataIn2 = 32'd1; 
32'd7029: dataIn2 = 32'd1; 
32'd7030: dataIn2 = 32'd0; 
32'd7031: dataIn2 = 32'd0; 
32'd7032: dataIn2 = 32'd1; 
32'd7033: dataIn2 = 32'd1; 
32'd7034: dataIn2 = 32'd1; 
32'd7035: dataIn2 = 32'd0; 
32'd7036: dataIn2 = 32'd1; 
32'd7037: dataIn2 = 32'd0; 
32'd7038: dataIn2 = 32'd1; 
32'd7039: dataIn2 = 32'd0; 
32'd7040: dataIn2 = 32'd0; 
32'd7041: dataIn2 = 32'd1; 
32'd7042: dataIn2 = 32'd1; 
32'd7043: dataIn2 = 32'd0; 
32'd7044: dataIn2 = 32'd1; 
32'd7045: dataIn2 = 32'd1; 
32'd7046: dataIn2 = 32'd1; 
32'd7047: dataIn2 = 32'd1; 
32'd7048: dataIn2 = 32'd1; 
32'd7049: dataIn2 = 32'd0; 
32'd7050: dataIn2 = 32'd0; 
32'd7051: dataIn2 = 32'd0; 
32'd7052: dataIn2 = 32'd1; 
32'd7053: dataIn2 = 32'd0; 
32'd7054: dataIn2 = 32'd1; 
32'd7055: dataIn2 = 32'd1; 
32'd7056: dataIn2 = 32'd0; 
32'd7057: dataIn2 = 32'd0; 
32'd7058: dataIn2 = 32'd1; 
32'd7059: dataIn2 = 32'd0; 
32'd7060: dataIn2 = 32'd1; 
32'd7061: dataIn2 = 32'd0; 
32'd7062: dataIn2 = 32'd1; 
32'd7063: dataIn2 = 32'd0; 
32'd7064: dataIn2 = 32'd0; 
32'd7065: dataIn2 = 32'd1; 
32'd7066: dataIn2 = 32'd1; 
32'd7067: dataIn2 = 32'd0; 
32'd7068: dataIn2 = 32'd1; 
32'd7069: dataIn2 = 32'd0; 
32'd7070: dataIn2 = 32'd0; 
32'd7071: dataIn2 = 32'd1; 
32'd7072: dataIn2 = 32'd1; 
32'd7073: dataIn2 = 32'd1; 
32'd7074: dataIn2 = 32'd0; 
32'd7075: dataIn2 = 32'd1; 
32'd7076: dataIn2 = 32'd1; 
32'd7077: dataIn2 = 32'd0; 
32'd7078: dataIn2 = 32'd0; 
32'd7079: dataIn2 = 32'd0; 
32'd7080: dataIn2 = 32'd0; 
32'd7081: dataIn2 = 32'd1; 
32'd7082: dataIn2 = 32'd0; 
32'd7083: dataIn2 = 32'd1; 
32'd7084: dataIn2 = 32'd1; 
32'd7085: dataIn2 = 32'd0; 
32'd7086: dataIn2 = 32'd1; 
32'd7087: dataIn2 = 32'd0; 
32'd7088: dataIn2 = 32'd0; 
32'd7089: dataIn2 = 32'd1; 
32'd7090: dataIn2 = 32'd1; 
32'd7091: dataIn2 = 32'd1; 
32'd7092: dataIn2 = 32'd1; 
32'd7093: dataIn2 = 32'd0; 
32'd7094: dataIn2 = 32'd1; 
32'd7095: dataIn2 = 32'd0; 
32'd7096: dataIn2 = 32'd1; 
32'd7097: dataIn2 = 32'd0; 
32'd7098: dataIn2 = 32'd1; 
32'd7099: dataIn2 = 32'd1; 
32'd7100: dataIn2 = 32'd1; 
32'd7101: dataIn2 = 32'd0; 
32'd7102: dataIn2 = 32'd0; 
32'd7103: dataIn2 = 32'd0; 
32'd7104: dataIn2 = 32'd0; 
32'd7105: dataIn2 = 32'd1; 
32'd7106: dataIn2 = 32'd1; 
32'd7107: dataIn2 = 32'd1; 
32'd7108: dataIn2 = 32'd1; 
32'd7109: dataIn2 = 32'd1; 
32'd7110: dataIn2 = 32'd1; 
32'd7111: dataIn2 = 32'd0; 
32'd7112: dataIn2 = 32'd0; 
32'd7113: dataIn2 = 32'd1; 
32'd7114: dataIn2 = 32'd1; 
32'd7115: dataIn2 = 32'd1; 
32'd7116: dataIn2 = 32'd1; 
32'd7117: dataIn2 = 32'd0; 
32'd7118: dataIn2 = 32'd0; 
32'd7119: dataIn2 = 32'd1; 
32'd7120: dataIn2 = 32'd0; 
32'd7121: dataIn2 = 32'd1; 
32'd7122: dataIn2 = 32'd0; 
32'd7123: dataIn2 = 32'd0; 
32'd7124: dataIn2 = 32'd1; 
32'd7125: dataIn2 = 32'd1; 
32'd7126: dataIn2 = 32'd1; 
32'd7127: dataIn2 = 32'd0; 
32'd7128: dataIn2 = 32'd1; 
32'd7129: dataIn2 = 32'd0; 
32'd7130: dataIn2 = 32'd0; 
32'd7131: dataIn2 = 32'd1; 
32'd7132: dataIn2 = 32'd1; 
32'd7133: dataIn2 = 32'd0; 
32'd7134: dataIn2 = 32'd1; 
32'd7135: dataIn2 = 32'd0; 
32'd7136: dataIn2 = 32'd0; 
32'd7137: dataIn2 = 32'd1; 
32'd7138: dataIn2 = 32'd0; 
32'd7139: dataIn2 = 32'd1; 
32'd7140: dataIn2 = 32'd0; 
32'd7141: dataIn2 = 32'd0; 
32'd7142: dataIn2 = 32'd0; 
32'd7143: dataIn2 = 32'd1; 
32'd7144: dataIn2 = 32'd1; 
32'd7145: dataIn2 = 32'd0; 
32'd7146: dataIn2 = 32'd0; 
32'd7147: dataIn2 = 32'd0; 
32'd7148: dataIn2 = 32'd1; 
32'd7149: dataIn2 = 32'd1; 
32'd7150: dataIn2 = 32'd0; 
32'd7151: dataIn2 = 32'd1; 
32'd7152: dataIn2 = 32'd1; 
32'd7153: dataIn2 = 32'd0; 
32'd7154: dataIn2 = 32'd1; 
32'd7155: dataIn2 = 32'd0; 
32'd7156: dataIn2 = 32'd0; 
32'd7157: dataIn2 = 32'd0; 
32'd7158: dataIn2 = 32'd0; 
32'd7159: dataIn2 = 32'd0; 
32'd7160: dataIn2 = 32'd0; 
32'd7161: dataIn2 = 32'd1; 
32'd7162: dataIn2 = 32'd1; 
32'd7163: dataIn2 = 32'd1; 
32'd7164: dataIn2 = 32'd0; 
32'd7165: dataIn2 = 32'd1; 
32'd7166: dataIn2 = 32'd1; 
32'd7167: dataIn2 = 32'd1; 
32'd7168: dataIn2 = 32'd0; 
32'd7169: dataIn2 = 32'd0; 
32'd7170: dataIn2 = 32'd1; 
32'd7171: dataIn2 = 32'd0; 
32'd7172: dataIn2 = 32'd0; 
32'd7173: dataIn2 = 32'd1; 
32'd7174: dataIn2 = 32'd1; 
32'd7175: dataIn2 = 32'd0; 
32'd7176: dataIn2 = 32'd0; 
32'd7177: dataIn2 = 32'd1; 
32'd7178: dataIn2 = 32'd0; 
32'd7179: dataIn2 = 32'd0; 
32'd7180: dataIn2 = 32'd1; 
32'd7181: dataIn2 = 32'd0; 
32'd7182: dataIn2 = 32'd0; 
32'd7183: dataIn2 = 32'd0; 
32'd7184: dataIn2 = 32'd0; 
32'd7185: dataIn2 = 32'd0; 
32'd7186: dataIn2 = 32'd0; 
32'd7187: dataIn2 = 32'd1; 
32'd7188: dataIn2 = 32'd0; 
32'd7189: dataIn2 = 32'd0; 
32'd7190: dataIn2 = 32'd1; 
32'd7191: dataIn2 = 32'd0; 
32'd7192: dataIn2 = 32'd0; 
32'd7193: dataIn2 = 32'd0; 
32'd7194: dataIn2 = 32'd0; 
32'd7195: dataIn2 = 32'd1; 
32'd7196: dataIn2 = 32'd0; 
32'd7197: dataIn2 = 32'd0; 
32'd7198: dataIn2 = 32'd1; 
32'd7199: dataIn2 = 32'd0; 
32'd7200: dataIn2 = 32'd1; 
32'd7201: dataIn2 = 32'd1; 
32'd7202: dataIn2 = 32'd0; 
32'd7203: dataIn2 = 32'd0; 
32'd7204: dataIn2 = 32'd0; 
32'd7205: dataIn2 = 32'd0; 
32'd7206: dataIn2 = 32'd0; 
32'd7207: dataIn2 = 32'd1; 
32'd7208: dataIn2 = 32'd0; 
32'd7209: dataIn2 = 32'd1; 
32'd7210: dataIn2 = 32'd1; 
32'd7211: dataIn2 = 32'd1; 
32'd7212: dataIn2 = 32'd1; 
32'd7213: dataIn2 = 32'd0; 
32'd7214: dataIn2 = 32'd0; 
32'd7215: dataIn2 = 32'd0; 
32'd7216: dataIn2 = 32'd0; 
32'd7217: dataIn2 = 32'd0; 
32'd7218: dataIn2 = 32'd0; 
32'd7219: dataIn2 = 32'd1; 
32'd7220: dataIn2 = 32'd1; 
32'd7221: dataIn2 = 32'd1; 
32'd7222: dataIn2 = 32'd0; 
32'd7223: dataIn2 = 32'd1; 
32'd7224: dataIn2 = 32'd1; 
32'd7225: dataIn2 = 32'd0; 
32'd7226: dataIn2 = 32'd1; 
32'd7227: dataIn2 = 32'd1; 
32'd7228: dataIn2 = 32'd0; 
32'd7229: dataIn2 = 32'd0; 
32'd7230: dataIn2 = 32'd1; 
32'd7231: dataIn2 = 32'd0; 
32'd7232: dataIn2 = 32'd1; 
32'd7233: dataIn2 = 32'd1; 
32'd7234: dataIn2 = 32'd1; 
32'd7235: dataIn2 = 32'd0; 
32'd7236: dataIn2 = 32'd1; 
32'd7237: dataIn2 = 32'd1; 
32'd7238: dataIn2 = 32'd1; 
32'd7239: dataIn2 = 32'd1; 
32'd7240: dataIn2 = 32'd1; 
32'd7241: dataIn2 = 32'd1; 
32'd7242: dataIn2 = 32'd0; 
32'd7243: dataIn2 = 32'd0; 
32'd7244: dataIn2 = 32'd0; 
32'd7245: dataIn2 = 32'd0; 
32'd7246: dataIn2 = 32'd1; 
32'd7247: dataIn2 = 32'd1; 
32'd7248: dataIn2 = 32'd1; 
32'd7249: dataIn2 = 32'd0; 
32'd7250: dataIn2 = 32'd1; 
32'd7251: dataIn2 = 32'd0; 
32'd7252: dataIn2 = 32'd0; 
32'd7253: dataIn2 = 32'd1; 
32'd7254: dataIn2 = 32'd1; 
32'd7255: dataIn2 = 32'd0; 
32'd7256: dataIn2 = 32'd0; 
32'd7257: dataIn2 = 32'd1; 
32'd7258: dataIn2 = 32'd1; 
32'd7259: dataIn2 = 32'd0; 
32'd7260: dataIn2 = 32'd1; 
32'd7261: dataIn2 = 32'd1; 
32'd7262: dataIn2 = 32'd1; 
32'd7263: dataIn2 = 32'd1; 
32'd7264: dataIn2 = 32'd1; 
32'd7265: dataIn2 = 32'd0; 
32'd7266: dataIn2 = 32'd1; 
32'd7267: dataIn2 = 32'd0; 
32'd7268: dataIn2 = 32'd1; 
32'd7269: dataIn2 = 32'd0; 
32'd7270: dataIn2 = 32'd0; 
32'd7271: dataIn2 = 32'd1; 
32'd7272: dataIn2 = 32'd1; 
32'd7273: dataIn2 = 32'd0; 
32'd7274: dataIn2 = 32'd1; 
32'd7275: dataIn2 = 32'd0; 
32'd7276: dataIn2 = 32'd1; 
32'd7277: dataIn2 = 32'd1; 
32'd7278: dataIn2 = 32'd1; 
32'd7279: dataIn2 = 32'd0; 
32'd7280: dataIn2 = 32'd0; 
32'd7281: dataIn2 = 32'd1; 
32'd7282: dataIn2 = 32'd0; 
32'd7283: dataIn2 = 32'd0; 
32'd7284: dataIn2 = 32'd1; 
32'd7285: dataIn2 = 32'd1; 
32'd7286: dataIn2 = 32'd0; 
32'd7287: dataIn2 = 32'd0; 
32'd7288: dataIn2 = 32'd1; 
32'd7289: dataIn2 = 32'd0; 
32'd7290: dataIn2 = 32'd1; 
32'd7291: dataIn2 = 32'd1; 
32'd7292: dataIn2 = 32'd1; 
32'd7293: dataIn2 = 32'd1; 
32'd7294: dataIn2 = 32'd1; 
32'd7295: dataIn2 = 32'd1; 
32'd7296: dataIn2 = 32'd1; 
32'd7297: dataIn2 = 32'd0; 
32'd7298: dataIn2 = 32'd1; 
32'd7299: dataIn2 = 32'd1; 
32'd7300: dataIn2 = 32'd0; 
32'd7301: dataIn2 = 32'd0; 
32'd7302: dataIn2 = 32'd1; 
32'd7303: dataIn2 = 32'd0; 
32'd7304: dataIn2 = 32'd0; 
32'd7305: dataIn2 = 32'd1; 
32'd7306: dataIn2 = 32'd1; 
32'd7307: dataIn2 = 32'd1; 
32'd7308: dataIn2 = 32'd1; 
32'd7309: dataIn2 = 32'd1; 
32'd7310: dataIn2 = 32'd0; 
32'd7311: dataIn2 = 32'd0; 
32'd7312: dataIn2 = 32'd0; 
32'd7313: dataIn2 = 32'd0; 
32'd7314: dataIn2 = 32'd0; 
32'd7315: dataIn2 = 32'd0; 
32'd7316: dataIn2 = 32'd1; 
32'd7317: dataIn2 = 32'd1; 
32'd7318: dataIn2 = 32'd1; 
32'd7319: dataIn2 = 32'd0; 
32'd7320: dataIn2 = 32'd0; 
32'd7321: dataIn2 = 32'd0; 
32'd7322: dataIn2 = 32'd1; 
32'd7323: dataIn2 = 32'd0; 
32'd7324: dataIn2 = 32'd0; 
32'd7325: dataIn2 = 32'd0; 
32'd7326: dataIn2 = 32'd1; 
32'd7327: dataIn2 = 32'd1; 
32'd7328: dataIn2 = 32'd1; 
32'd7329: dataIn2 = 32'd0; 
32'd7330: dataIn2 = 32'd0; 
32'd7331: dataIn2 = 32'd0; 
32'd7332: dataIn2 = 32'd1; 
32'd7333: dataIn2 = 32'd0; 
32'd7334: dataIn2 = 32'd0; 
32'd7335: dataIn2 = 32'd1; 
32'd7336: dataIn2 = 32'd0; 
32'd7337: dataIn2 = 32'd0; 
32'd7338: dataIn2 = 32'd1; 
32'd7339: dataIn2 = 32'd0; 
32'd7340: dataIn2 = 32'd1; 
32'd7341: dataIn2 = 32'd0; 
32'd7342: dataIn2 = 32'd0; 
32'd7343: dataIn2 = 32'd1; 
32'd7344: dataIn2 = 32'd1; 
32'd7345: dataIn2 = 32'd0; 
32'd7346: dataIn2 = 32'd1; 
32'd7347: dataIn2 = 32'd1; 
32'd7348: dataIn2 = 32'd0; 
32'd7349: dataIn2 = 32'd1; 
32'd7350: dataIn2 = 32'd1; 
32'd7351: dataIn2 = 32'd0; 
32'd7352: dataIn2 = 32'd0; 
32'd7353: dataIn2 = 32'd1; 
32'd7354: dataIn2 = 32'd0; 
32'd7355: dataIn2 = 32'd0; 
32'd7356: dataIn2 = 32'd1; 
32'd7357: dataIn2 = 32'd1; 
32'd7358: dataIn2 = 32'd0; 
32'd7359: dataIn2 = 32'd1; 
32'd7360: dataIn2 = 32'd1; 
32'd7361: dataIn2 = 32'd1; 
32'd7362: dataIn2 = 32'd1; 
32'd7363: dataIn2 = 32'd1; 
32'd7364: dataIn2 = 32'd1; 
32'd7365: dataIn2 = 32'd0; 
32'd7366: dataIn2 = 32'd1; 
32'd7367: dataIn2 = 32'd0; 
32'd7368: dataIn2 = 32'd0; 
32'd7369: dataIn2 = 32'd0; 
32'd7370: dataIn2 = 32'd1; 
32'd7371: dataIn2 = 32'd0; 
32'd7372: dataIn2 = 32'd0; 
32'd7373: dataIn2 = 32'd1; 
32'd7374: dataIn2 = 32'd0; 
32'd7375: dataIn2 = 32'd0; 
32'd7376: dataIn2 = 32'd0; 
32'd7377: dataIn2 = 32'd0; 
32'd7378: dataIn2 = 32'd0; 
32'd7379: dataIn2 = 32'd0; 
32'd7380: dataIn2 = 32'd1; 
32'd7381: dataIn2 = 32'd0; 
32'd7382: dataIn2 = 32'd0; 
32'd7383: dataIn2 = 32'd1; 
32'd7384: dataIn2 = 32'd0; 
32'd7385: dataIn2 = 32'd1; 
32'd7386: dataIn2 = 32'd0; 
32'd7387: dataIn2 = 32'd0; 
32'd7388: dataIn2 = 32'd1; 
32'd7389: dataIn2 = 32'd0; 
32'd7390: dataIn2 = 32'd0; 
32'd7391: dataIn2 = 32'd0; 
32'd7392: dataIn2 = 32'd1; 
32'd7393: dataIn2 = 32'd1; 
32'd7394: dataIn2 = 32'd1; 
32'd7395: dataIn2 = 32'd1; 
32'd7396: dataIn2 = 32'd1; 
32'd7397: dataIn2 = 32'd1; 
32'd7398: dataIn2 = 32'd1; 
32'd7399: dataIn2 = 32'd1; 
32'd7400: dataIn2 = 32'd1; 
32'd7401: dataIn2 = 32'd0; 
32'd7402: dataIn2 = 32'd0; 
32'd7403: dataIn2 = 32'd1; 
32'd7404: dataIn2 = 32'd1; 
32'd7405: dataIn2 = 32'd1; 
32'd7406: dataIn2 = 32'd1; 
32'd7407: dataIn2 = 32'd1; 
32'd7408: dataIn2 = 32'd1; 
32'd7409: dataIn2 = 32'd0; 
32'd7410: dataIn2 = 32'd1; 
32'd7411: dataIn2 = 32'd0; 
32'd7412: dataIn2 = 32'd0; 
32'd7413: dataIn2 = 32'd0; 
32'd7414: dataIn2 = 32'd1; 
32'd7415: dataIn2 = 32'd1; 
32'd7416: dataIn2 = 32'd1; 
32'd7417: dataIn2 = 32'd1; 
32'd7418: dataIn2 = 32'd0; 
32'd7419: dataIn2 = 32'd1; 
32'd7420: dataIn2 = 32'd1; 
32'd7421: dataIn2 = 32'd1; 
32'd7422: dataIn2 = 32'd0; 
32'd7423: dataIn2 = 32'd0; 
32'd7424: dataIn2 = 32'd0; 
32'd7425: dataIn2 = 32'd0; 
32'd7426: dataIn2 = 32'd1; 
32'd7427: dataIn2 = 32'd0; 
32'd7428: dataIn2 = 32'd1; 
32'd7429: dataIn2 = 32'd1; 
32'd7430: dataIn2 = 32'd0; 
32'd7431: dataIn2 = 32'd1; 
32'd7432: dataIn2 = 32'd1; 
32'd7433: dataIn2 = 32'd1; 
32'd7434: dataIn2 = 32'd0; 
32'd7435: dataIn2 = 32'd1; 
32'd7436: dataIn2 = 32'd0; 
32'd7437: dataIn2 = 32'd0; 
32'd7438: dataIn2 = 32'd1; 
32'd7439: dataIn2 = 32'd0; 
32'd7440: dataIn2 = 32'd1; 
32'd7441: dataIn2 = 32'd1; 
32'd7442: dataIn2 = 32'd1; 
32'd7443: dataIn2 = 32'd0; 
32'd7444: dataIn2 = 32'd0; 
32'd7445: dataIn2 = 32'd1; 
32'd7446: dataIn2 = 32'd0; 
32'd7447: dataIn2 = 32'd1; 
32'd7448: dataIn2 = 32'd0; 
32'd7449: dataIn2 = 32'd0; 
32'd7450: dataIn2 = 32'd0; 
32'd7451: dataIn2 = 32'd1; 
32'd7452: dataIn2 = 32'd1; 
32'd7453: dataIn2 = 32'd0; 
32'd7454: dataIn2 = 32'd1; 
32'd7455: dataIn2 = 32'd1; 
32'd7456: dataIn2 = 32'd1; 
32'd7457: dataIn2 = 32'd0; 
32'd7458: dataIn2 = 32'd1; 
32'd7459: dataIn2 = 32'd1; 
32'd7460: dataIn2 = 32'd0; 
32'd7461: dataIn2 = 32'd1; 
32'd7462: dataIn2 = 32'd0; 
32'd7463: dataIn2 = 32'd0; 
32'd7464: dataIn2 = 32'd1; 
32'd7465: dataIn2 = 32'd1; 
32'd7466: dataIn2 = 32'd1; 
32'd7467: dataIn2 = 32'd0; 
32'd7468: dataIn2 = 32'd1; 
32'd7469: dataIn2 = 32'd0; 
32'd7470: dataIn2 = 32'd1; 
32'd7471: dataIn2 = 32'd0; 
32'd7472: dataIn2 = 32'd1; 
32'd7473: dataIn2 = 32'd0; 
32'd7474: dataIn2 = 32'd0; 
32'd7475: dataIn2 = 32'd0; 
32'd7476: dataIn2 = 32'd1; 
32'd7477: dataIn2 = 32'd1; 
32'd7478: dataIn2 = 32'd1; 
32'd7479: dataIn2 = 32'd1; 
32'd7480: dataIn2 = 32'd0; 
32'd7481: dataIn2 = 32'd0; 
32'd7482: dataIn2 = 32'd0; 
32'd7483: dataIn2 = 32'd1; 
32'd7484: dataIn2 = 32'd0; 
32'd7485: dataIn2 = 32'd1; 
32'd7486: dataIn2 = 32'd0; 
32'd7487: dataIn2 = 32'd0; 
32'd7488: dataIn2 = 32'd0; 
32'd7489: dataIn2 = 32'd0; 
32'd7490: dataIn2 = 32'd1; 
32'd7491: dataIn2 = 32'd0; 
32'd7492: dataIn2 = 32'd0; 
32'd7493: dataIn2 = 32'd1; 
32'd7494: dataIn2 = 32'd0; 
32'd7495: dataIn2 = 32'd0; 
32'd7496: dataIn2 = 32'd1; 
32'd7497: dataIn2 = 32'd0; 
32'd7498: dataIn2 = 32'd0; 
32'd7499: dataIn2 = 32'd1; 
32'd7500: dataIn2 = 32'd1; 
32'd7501: dataIn2 = 32'd0; 
32'd7502: dataIn2 = 32'd1; 
32'd7503: dataIn2 = 32'd1; 
32'd7504: dataIn2 = 32'd1; 
32'd7505: dataIn2 = 32'd1; 
32'd7506: dataIn2 = 32'd1; 
32'd7507: dataIn2 = 32'd0; 
32'd7508: dataIn2 = 32'd0; 
32'd7509: dataIn2 = 32'd1; 
32'd7510: dataIn2 = 32'd0; 
32'd7511: dataIn2 = 32'd0; 
32'd7512: dataIn2 = 32'd1; 
32'd7513: dataIn2 = 32'd1; 
32'd7514: dataIn2 = 32'd1; 
32'd7515: dataIn2 = 32'd0; 
32'd7516: dataIn2 = 32'd1; 
32'd7517: dataIn2 = 32'd0; 
32'd7518: dataIn2 = 32'd1; 
32'd7519: dataIn2 = 32'd1; 
32'd7520: dataIn2 = 32'd0; 
32'd7521: dataIn2 = 32'd1; 
32'd7522: dataIn2 = 32'd1; 
32'd7523: dataIn2 = 32'd1; 
32'd7524: dataIn2 = 32'd1; 
32'd7525: dataIn2 = 32'd0; 
32'd7526: dataIn2 = 32'd1; 
32'd7527: dataIn2 = 32'd0; 
32'd7528: dataIn2 = 32'd1; 
32'd7529: dataIn2 = 32'd0; 
32'd7530: dataIn2 = 32'd1; 
32'd7531: dataIn2 = 32'd0; 
32'd7532: dataIn2 = 32'd0; 
32'd7533: dataIn2 = 32'd0; 
32'd7534: dataIn2 = 32'd0; 
32'd7535: dataIn2 = 32'd0; 
32'd7536: dataIn2 = 32'd1; 
32'd7537: dataIn2 = 32'd0; 
32'd7538: dataIn2 = 32'd1; 
32'd7539: dataIn2 = 32'd0; 
32'd7540: dataIn2 = 32'd0; 
32'd7541: dataIn2 = 32'd0; 
32'd7542: dataIn2 = 32'd1; 
32'd7543: dataIn2 = 32'd0; 
32'd7544: dataIn2 = 32'd1; 
32'd7545: dataIn2 = 32'd1; 
32'd7546: dataIn2 = 32'd0; 
32'd7547: dataIn2 = 32'd1; 
32'd7548: dataIn2 = 32'd0; 
32'd7549: dataIn2 = 32'd1; 
32'd7550: dataIn2 = 32'd1; 
32'd7551: dataIn2 = 32'd0; 
32'd7552: dataIn2 = 32'd1; 
32'd7553: dataIn2 = 32'd1; 
32'd7554: dataIn2 = 32'd0; 
32'd7555: dataIn2 = 32'd1; 
32'd7556: dataIn2 = 32'd0; 
32'd7557: dataIn2 = 32'd1; 
32'd7558: dataIn2 = 32'd1; 
32'd7559: dataIn2 = 32'd0; 
32'd7560: dataIn2 = 32'd0; 
32'd7561: dataIn2 = 32'd0; 
32'd7562: dataIn2 = 32'd1; 
32'd7563: dataIn2 = 32'd0; 
32'd7564: dataIn2 = 32'd1; 
32'd7565: dataIn2 = 32'd0; 
32'd7566: dataIn2 = 32'd0; 
32'd7567: dataIn2 = 32'd0; 
32'd7568: dataIn2 = 32'd0; 
32'd7569: dataIn2 = 32'd0; 
32'd7570: dataIn2 = 32'd1; 
32'd7571: dataIn2 = 32'd1; 
32'd7572: dataIn2 = 32'd1; 
32'd7573: dataIn2 = 32'd1; 
32'd7574: dataIn2 = 32'd1; 
32'd7575: dataIn2 = 32'd0; 
32'd7576: dataIn2 = 32'd1; 
32'd7577: dataIn2 = 32'd0; 
32'd7578: dataIn2 = 32'd0; 
32'd7579: dataIn2 = 32'd1; 
32'd7580: dataIn2 = 32'd0; 
32'd7581: dataIn2 = 32'd0; 
32'd7582: dataIn2 = 32'd1; 
32'd7583: dataIn2 = 32'd1; 
32'd7584: dataIn2 = 32'd0; 
32'd7585: dataIn2 = 32'd0; 
32'd7586: dataIn2 = 32'd0; 
32'd7587: dataIn2 = 32'd1; 
32'd7588: dataIn2 = 32'd1; 
32'd7589: dataIn2 = 32'd0; 
32'd7590: dataIn2 = 32'd1; 
32'd7591: dataIn2 = 32'd1; 
32'd7592: dataIn2 = 32'd0; 
32'd7593: dataIn2 = 32'd1; 
32'd7594: dataIn2 = 32'd1; 
32'd7595: dataIn2 = 32'd1; 
32'd7596: dataIn2 = 32'd1; 
32'd7597: dataIn2 = 32'd1; 
32'd7598: dataIn2 = 32'd1; 
32'd7599: dataIn2 = 32'd1; 
32'd7600: dataIn2 = 32'd1; 
32'd7601: dataIn2 = 32'd0; 
32'd7602: dataIn2 = 32'd1; 
32'd7603: dataIn2 = 32'd0; 
32'd7604: dataIn2 = 32'd1; 
32'd7605: dataIn2 = 32'd0; 
32'd7606: dataIn2 = 32'd0; 
32'd7607: dataIn2 = 32'd1; 
32'd7608: dataIn2 = 32'd1; 
32'd7609: dataIn2 = 32'd0; 
32'd7610: dataIn2 = 32'd1; 
32'd7611: dataIn2 = 32'd1; 
32'd7612: dataIn2 = 32'd0; 
32'd7613: dataIn2 = 32'd1; 
32'd7614: dataIn2 = 32'd0; 
32'd7615: dataIn2 = 32'd1; 
32'd7616: dataIn2 = 32'd0; 
32'd7617: dataIn2 = 32'd0; 
32'd7618: dataIn2 = 32'd1; 
32'd7619: dataIn2 = 32'd1; 
32'd7620: dataIn2 = 32'd1; 
32'd7621: dataIn2 = 32'd0; 
32'd7622: dataIn2 = 32'd0; 
32'd7623: dataIn2 = 32'd0; 
32'd7624: dataIn2 = 32'd0; 
32'd7625: dataIn2 = 32'd1; 
32'd7626: dataIn2 = 32'd0; 
32'd7627: dataIn2 = 32'd0; 
32'd7628: dataIn2 = 32'd0; 
32'd7629: dataIn2 = 32'd1; 
32'd7630: dataIn2 = 32'd0; 
32'd7631: dataIn2 = 32'd1; 
32'd7632: dataIn2 = 32'd0; 
32'd7633: dataIn2 = 32'd0; 
32'd7634: dataIn2 = 32'd0; 
32'd7635: dataIn2 = 32'd0; 
32'd7636: dataIn2 = 32'd0; 
32'd7637: dataIn2 = 32'd1; 
32'd7638: dataIn2 = 32'd1; 
32'd7639: dataIn2 = 32'd1; 
32'd7640: dataIn2 = 32'd1; 
32'd7641: dataIn2 = 32'd1; 
32'd7642: dataIn2 = 32'd1; 
32'd7643: dataIn2 = 32'd1; 
32'd7644: dataIn2 = 32'd1; 
32'd7645: dataIn2 = 32'd1; 
32'd7646: dataIn2 = 32'd1; 
32'd7647: dataIn2 = 32'd1; 
32'd7648: dataIn2 = 32'd0; 
32'd7649: dataIn2 = 32'd1; 
32'd7650: dataIn2 = 32'd0; 
32'd7651: dataIn2 = 32'd0; 
32'd7652: dataIn2 = 32'd0; 
32'd7653: dataIn2 = 32'd1; 
32'd7654: dataIn2 = 32'd0; 
32'd7655: dataIn2 = 32'd1; 
32'd7656: dataIn2 = 32'd0; 
32'd7657: dataIn2 = 32'd0; 
32'd7658: dataIn2 = 32'd1; 
32'd7659: dataIn2 = 32'd1; 
32'd7660: dataIn2 = 32'd1; 
32'd7661: dataIn2 = 32'd1; 
32'd7662: dataIn2 = 32'd1; 
32'd7663: dataIn2 = 32'd0; 
32'd7664: dataIn2 = 32'd1; 
32'd7665: dataIn2 = 32'd0; 
32'd7666: dataIn2 = 32'd0; 
32'd7667: dataIn2 = 32'd0; 
32'd7668: dataIn2 = 32'd0; 
32'd7669: dataIn2 = 32'd0; 
32'd7670: dataIn2 = 32'd1; 
32'd7671: dataIn2 = 32'd1; 
32'd7672: dataIn2 = 32'd0; 
32'd7673: dataIn2 = 32'd0; 
32'd7674: dataIn2 = 32'd1; 
32'd7675: dataIn2 = 32'd0; 
32'd7676: dataIn2 = 32'd0; 
32'd7677: dataIn2 = 32'd0; 
32'd7678: dataIn2 = 32'd0; 
32'd7679: dataIn2 = 32'd0; 
32'd7680: dataIn2 = 32'd1; 
32'd7681: dataIn2 = 32'd1; 
32'd7682: dataIn2 = 32'd0; 
32'd7683: dataIn2 = 32'd0; 
32'd7684: dataIn2 = 32'd0; 
32'd7685: dataIn2 = 32'd0; 
32'd7686: dataIn2 = 32'd1; 
32'd7687: dataIn2 = 32'd0; 
32'd7688: dataIn2 = 32'd0; 
32'd7689: dataIn2 = 32'd1; 
32'd7690: dataIn2 = 32'd1; 
32'd7691: dataIn2 = 32'd1; 
32'd7692: dataIn2 = 32'd1; 
32'd7693: dataIn2 = 32'd1; 
32'd7694: dataIn2 = 32'd1; 
32'd7695: dataIn2 = 32'd1; 
32'd7696: dataIn2 = 32'd0; 
32'd7697: dataIn2 = 32'd0; 
32'd7698: dataIn2 = 32'd0; 
32'd7699: dataIn2 = 32'd1; 
32'd7700: dataIn2 = 32'd1; 
32'd7701: dataIn2 = 32'd1; 
32'd7702: dataIn2 = 32'd0; 
32'd7703: dataIn2 = 32'd0; 
32'd7704: dataIn2 = 32'd0; 
32'd7705: dataIn2 = 32'd0; 
32'd7706: dataIn2 = 32'd0; 
32'd7707: dataIn2 = 32'd1; 
32'd7708: dataIn2 = 32'd1; 
32'd7709: dataIn2 = 32'd1; 
32'd7710: dataIn2 = 32'd0; 
32'd7711: dataIn2 = 32'd1; 
32'd7712: dataIn2 = 32'd0; 
32'd7713: dataIn2 = 32'd1; 
32'd7714: dataIn2 = 32'd1; 
32'd7715: dataIn2 = 32'd0; 
32'd7716: dataIn2 = 32'd1; 
32'd7717: dataIn2 = 32'd0; 
32'd7718: dataIn2 = 32'd1; 
32'd7719: dataIn2 = 32'd1; 
32'd7720: dataIn2 = 32'd0; 
32'd7721: dataIn2 = 32'd0; 
32'd7722: dataIn2 = 32'd1; 
32'd7723: dataIn2 = 32'd0; 
32'd7724: dataIn2 = 32'd0; 
32'd7725: dataIn2 = 32'd1; 
32'd7726: dataIn2 = 32'd1; 
32'd7727: dataIn2 = 32'd1; 
32'd7728: dataIn2 = 32'd1; 
32'd7729: dataIn2 = 32'd1; 
32'd7730: dataIn2 = 32'd1; 
32'd7731: dataIn2 = 32'd1; 
32'd7732: dataIn2 = 32'd0; 
32'd7733: dataIn2 = 32'd0; 
32'd7734: dataIn2 = 32'd0; 
32'd7735: dataIn2 = 32'd0; 
32'd7736: dataIn2 = 32'd1; 
32'd7737: dataIn2 = 32'd0; 
32'd7738: dataIn2 = 32'd1; 
32'd7739: dataIn2 = 32'd0; 
32'd7740: dataIn2 = 32'd1; 
32'd7741: dataIn2 = 32'd1; 
32'd7742: dataIn2 = 32'd1; 
32'd7743: dataIn2 = 32'd0; 
32'd7744: dataIn2 = 32'd0; 
32'd7745: dataIn2 = 32'd1; 
32'd7746: dataIn2 = 32'd1; 
32'd7747: dataIn2 = 32'd0; 
32'd7748: dataIn2 = 32'd1; 
32'd7749: dataIn2 = 32'd1; 
32'd7750: dataIn2 = 32'd1; 
32'd7751: dataIn2 = 32'd1; 
32'd7752: dataIn2 = 32'd0; 
32'd7753: dataIn2 = 32'd1; 
32'd7754: dataIn2 = 32'd1; 
32'd7755: dataIn2 = 32'd0; 
32'd7756: dataIn2 = 32'd0; 
32'd7757: dataIn2 = 32'd0; 
32'd7758: dataIn2 = 32'd1; 
32'd7759: dataIn2 = 32'd0; 
32'd7760: dataIn2 = 32'd1; 
32'd7761: dataIn2 = 32'd1; 
32'd7762: dataIn2 = 32'd1; 
32'd7763: dataIn2 = 32'd1; 
32'd7764: dataIn2 = 32'd0; 
32'd7765: dataIn2 = 32'd0; 
32'd7766: dataIn2 = 32'd0; 
32'd7767: dataIn2 = 32'd1; 
32'd7768: dataIn2 = 32'd1; 
32'd7769: dataIn2 = 32'd1; 
32'd7770: dataIn2 = 32'd0; 
32'd7771: dataIn2 = 32'd1; 
32'd7772: dataIn2 = 32'd1; 
32'd7773: dataIn2 = 32'd1; 
32'd7774: dataIn2 = 32'd1; 
32'd7775: dataIn2 = 32'd0; 
32'd7776: dataIn2 = 32'd0; 
32'd7777: dataIn2 = 32'd0; 
32'd7778: dataIn2 = 32'd0; 
32'd7779: dataIn2 = 32'd1; 
32'd7780: dataIn2 = 32'd1; 
32'd7781: dataIn2 = 32'd1; 
32'd7782: dataIn2 = 32'd0; 
32'd7783: dataIn2 = 32'd1; 
32'd7784: dataIn2 = 32'd1; 
32'd7785: dataIn2 = 32'd1; 
32'd7786: dataIn2 = 32'd1; 
32'd7787: dataIn2 = 32'd0; 
32'd7788: dataIn2 = 32'd1; 
32'd7789: dataIn2 = 32'd0; 
32'd7790: dataIn2 = 32'd1; 
32'd7791: dataIn2 = 32'd1; 
32'd7792: dataIn2 = 32'd0; 
32'd7793: dataIn2 = 32'd1; 
32'd7794: dataIn2 = 32'd0; 
32'd7795: dataIn2 = 32'd1; 
32'd7796: dataIn2 = 32'd1; 
32'd7797: dataIn2 = 32'd1; 
32'd7798: dataIn2 = 32'd0; 
32'd7799: dataIn2 = 32'd1; 
32'd7800: dataIn2 = 32'd1; 
32'd7801: dataIn2 = 32'd0; 
32'd7802: dataIn2 = 32'd0; 
32'd7803: dataIn2 = 32'd1; 
32'd7804: dataIn2 = 32'd0; 
32'd7805: dataIn2 = 32'd0; 
32'd7806: dataIn2 = 32'd1; 
32'd7807: dataIn2 = 32'd1; 
32'd7808: dataIn2 = 32'd0; 
32'd7809: dataIn2 = 32'd0; 
32'd7810: dataIn2 = 32'd0; 
32'd7811: dataIn2 = 32'd1; 
32'd7812: dataIn2 = 32'd0; 
32'd7813: dataIn2 = 32'd0; 
32'd7814: dataIn2 = 32'd0; 
32'd7815: dataIn2 = 32'd1; 
32'd7816: dataIn2 = 32'd0; 
32'd7817: dataIn2 = 32'd1; 
32'd7818: dataIn2 = 32'd1; 
32'd7819: dataIn2 = 32'd0; 
32'd7820: dataIn2 = 32'd1; 
32'd7821: dataIn2 = 32'd0; 
32'd7822: dataIn2 = 32'd0; 
32'd7823: dataIn2 = 32'd1; 
32'd7824: dataIn2 = 32'd1; 
32'd7825: dataIn2 = 32'd1; 
32'd7826: dataIn2 = 32'd0; 
32'd7827: dataIn2 = 32'd0; 
32'd7828: dataIn2 = 32'd1; 
32'd7829: dataIn2 = 32'd0; 
32'd7830: dataIn2 = 32'd1; 
32'd7831: dataIn2 = 32'd0; 
32'd7832: dataIn2 = 32'd0; 
32'd7833: dataIn2 = 32'd1; 
32'd7834: dataIn2 = 32'd0; 
32'd7835: dataIn2 = 32'd1; 
32'd7836: dataIn2 = 32'd0; 
32'd7837: dataIn2 = 32'd1; 
32'd7838: dataIn2 = 32'd1; 
32'd7839: dataIn2 = 32'd0; 
32'd7840: dataIn2 = 32'd1; 
32'd7841: dataIn2 = 32'd1; 
32'd7842: dataIn2 = 32'd0; 
32'd7843: dataIn2 = 32'd0; 
32'd7844: dataIn2 = 32'd1; 
32'd7845: dataIn2 = 32'd1; 
32'd7846: dataIn2 = 32'd0; 
32'd7847: dataIn2 = 32'd0; 
32'd7848: dataIn2 = 32'd0; 
32'd7849: dataIn2 = 32'd1; 
32'd7850: dataIn2 = 32'd0; 
32'd7851: dataIn2 = 32'd0; 
32'd7852: dataIn2 = 32'd0; 
32'd7853: dataIn2 = 32'd1; 
32'd7854: dataIn2 = 32'd1; 
32'd7855: dataIn2 = 32'd0; 
32'd7856: dataIn2 = 32'd1; 
32'd7857: dataIn2 = 32'd1; 
32'd7858: dataIn2 = 32'd0; 
32'd7859: dataIn2 = 32'd1; 
32'd7860: dataIn2 = 32'd0; 
32'd7861: dataIn2 = 32'd0; 
32'd7862: dataIn2 = 32'd0; 
32'd7863: dataIn2 = 32'd0; 
32'd7864: dataIn2 = 32'd1; 
32'd7865: dataIn2 = 32'd1; 
32'd7866: dataIn2 = 32'd1; 
32'd7867: dataIn2 = 32'd0; 
32'd7868: dataIn2 = 32'd1; 
32'd7869: dataIn2 = 32'd0; 
32'd7870: dataIn2 = 32'd1; 
32'd7871: dataIn2 = 32'd0; 
32'd7872: dataIn2 = 32'd0; 
32'd7873: dataIn2 = 32'd0; 
32'd7874: dataIn2 = 32'd0; 
32'd7875: dataIn2 = 32'd1; 
32'd7876: dataIn2 = 32'd0; 
32'd7877: dataIn2 = 32'd1; 
32'd7878: dataIn2 = 32'd1; 
32'd7879: dataIn2 = 32'd0; 
32'd7880: dataIn2 = 32'd0; 
32'd7881: dataIn2 = 32'd1; 
32'd7882: dataIn2 = 32'd0; 
32'd7883: dataIn2 = 32'd1; 
32'd7884: dataIn2 = 32'd1; 
32'd7885: dataIn2 = 32'd0; 
32'd7886: dataIn2 = 32'd0; 
32'd7887: dataIn2 = 32'd1; 
32'd7888: dataIn2 = 32'd0; 
32'd7889: dataIn2 = 32'd0; 
32'd7890: dataIn2 = 32'd0; 
32'd7891: dataIn2 = 32'd1; 
32'd7892: dataIn2 = 32'd0; 
32'd7893: dataIn2 = 32'd1; 
32'd7894: dataIn2 = 32'd0; 
32'd7895: dataIn2 = 32'd1; 
32'd7896: dataIn2 = 32'd0; 
32'd7897: dataIn2 = 32'd0; 
32'd7898: dataIn2 = 32'd0; 
32'd7899: dataIn2 = 32'd1; 
32'd7900: dataIn2 = 32'd0; 
32'd7901: dataIn2 = 32'd1; 
32'd7902: dataIn2 = 32'd1; 
32'd7903: dataIn2 = 32'd1; 
32'd7904: dataIn2 = 32'd1; 
32'd7905: dataIn2 = 32'd1; 
32'd7906: dataIn2 = 32'd0; 
32'd7907: dataIn2 = 32'd1; 
32'd7908: dataIn2 = 32'd0; 
32'd7909: dataIn2 = 32'd0; 
32'd7910: dataIn2 = 32'd0; 
32'd7911: dataIn2 = 32'd1; 
32'd7912: dataIn2 = 32'd1; 
32'd7913: dataIn2 = 32'd0; 
32'd7914: dataIn2 = 32'd0; 
32'd7915: dataIn2 = 32'd0; 
32'd7916: dataIn2 = 32'd1; 
32'd7917: dataIn2 = 32'd0; 
32'd7918: dataIn2 = 32'd0; 
32'd7919: dataIn2 = 32'd0; 
32'd7920: dataIn2 = 32'd0; 
32'd7921: dataIn2 = 32'd1; 
32'd7922: dataIn2 = 32'd1; 
32'd7923: dataIn2 = 32'd1; 
32'd7924: dataIn2 = 32'd0; 
32'd7925: dataIn2 = 32'd1; 
32'd7926: dataIn2 = 32'd1; 
32'd7927: dataIn2 = 32'd1; 
32'd7928: dataIn2 = 32'd0; 
32'd7929: dataIn2 = 32'd0; 
32'd7930: dataIn2 = 32'd1; 
32'd7931: dataIn2 = 32'd0; 
32'd7932: dataIn2 = 32'd0; 
32'd7933: dataIn2 = 32'd0; 
32'd7934: dataIn2 = 32'd1; 
32'd7935: dataIn2 = 32'd1; 
32'd7936: dataIn2 = 32'd0; 
32'd7937: dataIn2 = 32'd0; 
32'd7938: dataIn2 = 32'd1; 
32'd7939: dataIn2 = 32'd0; 
32'd7940: dataIn2 = 32'd0; 
32'd7941: dataIn2 = 32'd1; 
32'd7942: dataIn2 = 32'd1; 
32'd7943: dataIn2 = 32'd0; 
32'd7944: dataIn2 = 32'd1; 
32'd7945: dataIn2 = 32'd1; 
32'd7946: dataIn2 = 32'd0; 
32'd7947: dataIn2 = 32'd0; 
32'd7948: dataIn2 = 32'd0; 
32'd7949: dataIn2 = 32'd1; 
32'd7950: dataIn2 = 32'd0; 
32'd7951: dataIn2 = 32'd0; 
32'd7952: dataIn2 = 32'd1; 
32'd7953: dataIn2 = 32'd0; 
32'd7954: dataIn2 = 32'd1; 
32'd7955: dataIn2 = 32'd1; 
32'd7956: dataIn2 = 32'd1; 
32'd7957: dataIn2 = 32'd0; 
32'd7958: dataIn2 = 32'd0; 
32'd7959: dataIn2 = 32'd1; 
32'd7960: dataIn2 = 32'd0; 
32'd7961: dataIn2 = 32'd0; 
32'd7962: dataIn2 = 32'd0; 
32'd7963: dataIn2 = 32'd1; 
32'd7964: dataIn2 = 32'd0; 
32'd7965: dataIn2 = 32'd1; 
32'd7966: dataIn2 = 32'd1; 
32'd7967: dataIn2 = 32'd1; 
32'd7968: dataIn2 = 32'd0; 
32'd7969: dataIn2 = 32'd1; 
32'd7970: dataIn2 = 32'd1; 
32'd7971: dataIn2 = 32'd1; 
32'd7972: dataIn2 = 32'd0; 
32'd7973: dataIn2 = 32'd1; 
32'd7974: dataIn2 = 32'd1; 
32'd7975: dataIn2 = 32'd0; 
32'd7976: dataIn2 = 32'd0; 
32'd7977: dataIn2 = 32'd0; 
32'd7978: dataIn2 = 32'd1; 
32'd7979: dataIn2 = 32'd0; 
32'd7980: dataIn2 = 32'd1; 
32'd7981: dataIn2 = 32'd0; 
32'd7982: dataIn2 = 32'd1; 
32'd7983: dataIn2 = 32'd0; 
32'd7984: dataIn2 = 32'd1; 
32'd7985: dataIn2 = 32'd1; 
32'd7986: dataIn2 = 32'd1; 
32'd7987: dataIn2 = 32'd1; 
32'd7988: dataIn2 = 32'd0; 
32'd7989: dataIn2 = 32'd1; 
32'd7990: dataIn2 = 32'd0; 
32'd7991: dataIn2 = 32'd0; 
32'd7992: dataIn2 = 32'd0; 
32'd7993: dataIn2 = 32'd1; 
32'd7994: dataIn2 = 32'd0; 
32'd7995: dataIn2 = 32'd0; 
32'd7996: dataIn2 = 32'd1; 
32'd7997: dataIn2 = 32'd0; 
32'd7998: dataIn2 = 32'd0; 
32'd7999: dataIn2 = 32'd1; 
32'd8000: dataIn2 = 32'd0; 
32'd8001: dataIn2 = 32'd0; 
32'd8002: dataIn2 = 32'd1; 
32'd8003: dataIn2 = 32'd1; 
32'd8004: dataIn2 = 32'd1; 
32'd8005: dataIn2 = 32'd1; 
32'd8006: dataIn2 = 32'd1; 
32'd8007: dataIn2 = 32'd0; 
32'd8008: dataIn2 = 32'd0; 
32'd8009: dataIn2 = 32'd1; 
32'd8010: dataIn2 = 32'd1; 
32'd8011: dataIn2 = 32'd1; 
32'd8012: dataIn2 = 32'd1; 
32'd8013: dataIn2 = 32'd0; 
32'd8014: dataIn2 = 32'd0; 
32'd8015: dataIn2 = 32'd0; 
32'd8016: dataIn2 = 32'd1; 
32'd8017: dataIn2 = 32'd1; 
32'd8018: dataIn2 = 32'd0; 
32'd8019: dataIn2 = 32'd1; 
32'd8020: dataIn2 = 32'd0; 
32'd8021: dataIn2 = 32'd0; 
32'd8022: dataIn2 = 32'd0; 
32'd8023: dataIn2 = 32'd1; 
32'd8024: dataIn2 = 32'd0; 
32'd8025: dataIn2 = 32'd0; 
32'd8026: dataIn2 = 32'd1; 
32'd8027: dataIn2 = 32'd0; 
32'd8028: dataIn2 = 32'd1; 
32'd8029: dataIn2 = 32'd1; 
32'd8030: dataIn2 = 32'd0; 
32'd8031: dataIn2 = 32'd0; 
32'd8032: dataIn2 = 32'd1; 
32'd8033: dataIn2 = 32'd0; 
32'd8034: dataIn2 = 32'd0; 
32'd8035: dataIn2 = 32'd1; 
32'd8036: dataIn2 = 32'd0; 
32'd8037: dataIn2 = 32'd0; 
32'd8038: dataIn2 = 32'd1; 
32'd8039: dataIn2 = 32'd1; 
32'd8040: dataIn2 = 32'd0; 
32'd8041: dataIn2 = 32'd1; 
32'd8042: dataIn2 = 32'd1; 
32'd8043: dataIn2 = 32'd0; 
32'd8044: dataIn2 = 32'd1; 
32'd8045: dataIn2 = 32'd1; 
32'd8046: dataIn2 = 32'd0; 
32'd8047: dataIn2 = 32'd1; 
32'd8048: dataIn2 = 32'd0; 
32'd8049: dataIn2 = 32'd0; 
32'd8050: dataIn2 = 32'd1; 
32'd8051: dataIn2 = 32'd1; 
32'd8052: dataIn2 = 32'd0; 
32'd8053: dataIn2 = 32'd1; 
32'd8054: dataIn2 = 32'd0; 
32'd8055: dataIn2 = 32'd1; 
32'd8056: dataIn2 = 32'd0; 
32'd8057: dataIn2 = 32'd1; 
32'd8058: dataIn2 = 32'd1; 
32'd8059: dataIn2 = 32'd0; 
32'd8060: dataIn2 = 32'd1; 
32'd8061: dataIn2 = 32'd1; 
32'd8062: dataIn2 = 32'd1; 
32'd8063: dataIn2 = 32'd1; 
32'd8064: dataIn2 = 32'd0; 
32'd8065: dataIn2 = 32'd1; 
32'd8066: dataIn2 = 32'd0; 
32'd8067: dataIn2 = 32'd0; 
32'd8068: dataIn2 = 32'd0; 
32'd8069: dataIn2 = 32'd1; 
32'd8070: dataIn2 = 32'd1; 
32'd8071: dataIn2 = 32'd0; 
32'd8072: dataIn2 = 32'd1; 
32'd8073: dataIn2 = 32'd1; 
32'd8074: dataIn2 = 32'd1; 
32'd8075: dataIn2 = 32'd1; 
32'd8076: dataIn2 = 32'd1; 
32'd8077: dataIn2 = 32'd1; 
32'd8078: dataIn2 = 32'd0; 
32'd8079: dataIn2 = 32'd1; 
32'd8080: dataIn2 = 32'd1; 
32'd8081: dataIn2 = 32'd1; 
32'd8082: dataIn2 = 32'd0; 
32'd8083: dataIn2 = 32'd1; 
32'd8084: dataIn2 = 32'd1; 
32'd8085: dataIn2 = 32'd1; 
32'd8086: dataIn2 = 32'd0; 
32'd8087: dataIn2 = 32'd1; 
32'd8088: dataIn2 = 32'd0; 
32'd8089: dataIn2 = 32'd1; 
32'd8090: dataIn2 = 32'd0; 
32'd8091: dataIn2 = 32'd1; 
32'd8092: dataIn2 = 32'd0; 
32'd8093: dataIn2 = 32'd0; 
32'd8094: dataIn2 = 32'd1; 
32'd8095: dataIn2 = 32'd1; 
32'd8096: dataIn2 = 32'd1; 
32'd8097: dataIn2 = 32'd0; 
32'd8098: dataIn2 = 32'd1; 
32'd8099: dataIn2 = 32'd0; 
32'd8100: dataIn2 = 32'd1; 
32'd8101: dataIn2 = 32'd1; 
32'd8102: dataIn2 = 32'd0; 
32'd8103: dataIn2 = 32'd0; 
32'd8104: dataIn2 = 32'd0; 
32'd8105: dataIn2 = 32'd1; 
32'd8106: dataIn2 = 32'd0; 
32'd8107: dataIn2 = 32'd0; 
32'd8108: dataIn2 = 32'd0; 
32'd8109: dataIn2 = 32'd0; 
32'd8110: dataIn2 = 32'd1; 
32'd8111: dataIn2 = 32'd1; 
32'd8112: dataIn2 = 32'd1; 
32'd8113: dataIn2 = 32'd0; 
32'd8114: dataIn2 = 32'd0; 
32'd8115: dataIn2 = 32'd0; 
32'd8116: dataIn2 = 32'd1; 
32'd8117: dataIn2 = 32'd1; 
32'd8118: dataIn2 = 32'd1; 
32'd8119: dataIn2 = 32'd0; 
32'd8120: dataIn2 = 32'd0; 
32'd8121: dataIn2 = 32'd1; 
32'd8122: dataIn2 = 32'd0; 
32'd8123: dataIn2 = 32'd1; 
32'd8124: dataIn2 = 32'd0; 
32'd8125: dataIn2 = 32'd1; 
32'd8126: dataIn2 = 32'd0; 
32'd8127: dataIn2 = 32'd1; 
32'd8128: dataIn2 = 32'd1; 
32'd8129: dataIn2 = 32'd0; 
32'd8130: dataIn2 = 32'd1; 
32'd8131: dataIn2 = 32'd1; 
32'd8132: dataIn2 = 32'd0; 
32'd8133: dataIn2 = 32'd0; 
32'd8134: dataIn2 = 32'd1; 
32'd8135: dataIn2 = 32'd0; 
32'd8136: dataIn2 = 32'd0; 
32'd8137: dataIn2 = 32'd1; 
32'd8138: dataIn2 = 32'd0; 
32'd8139: dataIn2 = 32'd1; 
32'd8140: dataIn2 = 32'd1; 
32'd8141: dataIn2 = 32'd1; 
32'd8142: dataIn2 = 32'd0; 
32'd8143: dataIn2 = 32'd0; 
32'd8144: dataIn2 = 32'd1; 
32'd8145: dataIn2 = 32'd0; 
32'd8146: dataIn2 = 32'd1; 
32'd8147: dataIn2 = 32'd1; 
32'd8148: dataIn2 = 32'd0; 
32'd8149: dataIn2 = 32'd0; 
32'd8150: dataIn2 = 32'd0; 
32'd8151: dataIn2 = 32'd0; 
32'd8152: dataIn2 = 32'd1; 
32'd8153: dataIn2 = 32'd1; 
32'd8154: dataIn2 = 32'd1; 
32'd8155: dataIn2 = 32'd1; 
32'd8156: dataIn2 = 32'd1; 
32'd8157: dataIn2 = 32'd0; 
32'd8158: dataIn2 = 32'd0; 
32'd8159: dataIn2 = 32'd1; 
32'd8160: dataIn2 = 32'd0; 
32'd8161: dataIn2 = 32'd1; 
32'd8162: dataIn2 = 32'd1; 
32'd8163: dataIn2 = 32'd0; 
32'd8164: dataIn2 = 32'd0; 
32'd8165: dataIn2 = 32'd0; 
32'd8166: dataIn2 = 32'd0; 
32'd8167: dataIn2 = 32'd0; 
32'd8168: dataIn2 = 32'd1; 
32'd8169: dataIn2 = 32'd1; 
32'd8170: dataIn2 = 32'd0; 
32'd8171: dataIn2 = 32'd0; 
32'd8172: dataIn2 = 32'd1; 
32'd8173: dataIn2 = 32'd1; 
32'd8174: dataIn2 = 32'd0; 
32'd8175: dataIn2 = 32'd1; 
32'd8176: dataIn2 = 32'd1; 
32'd8177: dataIn2 = 32'd0; 
32'd8178: dataIn2 = 32'd1; 
32'd8179: dataIn2 = 32'd0; 
32'd8180: dataIn2 = 32'd0; 
32'd8181: dataIn2 = 32'd1; 
32'd8182: dataIn2 = 32'd0; 
32'd8183: dataIn2 = 32'd0; 
32'd8184: dataIn2 = 32'd1; 
32'd8185: dataIn2 = 32'd1; 
32'd8186: dataIn2 = 32'd1; 
32'd8187: dataIn2 = 32'd1; 
32'd8188: dataIn2 = 32'd0; 
32'd8189: dataIn2 = 32'd1; 
32'd8190: dataIn2 = 32'd1; 
32'd8191: dataIn2 = 32'd0; 
32'd8192: dataIn2 = 32'd0; 
32'd8193: dataIn2 = 32'd1; 
32'd8194: dataIn2 = 32'd0; 
32'd8195: dataIn2 = 32'd0; 
32'd8196: dataIn2 = 32'd0; 
32'd8197: dataIn2 = 32'd1; 
32'd8198: dataIn2 = 32'd1; 
32'd8199: dataIn2 = 32'd0; 
32'd8200: dataIn2 = 32'd1; 
32'd8201: dataIn2 = 32'd0; 
32'd8202: dataIn2 = 32'd0; 
32'd8203: dataIn2 = 32'd0; 
32'd8204: dataIn2 = 32'd1; 
32'd8205: dataIn2 = 32'd1; 
32'd8206: dataIn2 = 32'd0; 
32'd8207: dataIn2 = 32'd1; 
32'd8208: dataIn2 = 32'd1; 
32'd8209: dataIn2 = 32'd1; 
32'd8210: dataIn2 = 32'd1; 
32'd8211: dataIn2 = 32'd0; 
32'd8212: dataIn2 = 32'd0; 
32'd8213: dataIn2 = 32'd0; 
32'd8214: dataIn2 = 32'd1; 
32'd8215: dataIn2 = 32'd0; 
32'd8216: dataIn2 = 32'd1; 
32'd8217: dataIn2 = 32'd1; 
32'd8218: dataIn2 = 32'd1; 
32'd8219: dataIn2 = 32'd1; 
32'd8220: dataIn2 = 32'd0; 
32'd8221: dataIn2 = 32'd0; 
32'd8222: dataIn2 = 32'd0; 
32'd8223: dataIn2 = 32'd1; 
32'd8224: dataIn2 = 32'd0; 
32'd8225: dataIn2 = 32'd1; 
32'd8226: dataIn2 = 32'd1; 
32'd8227: dataIn2 = 32'd1; 
32'd8228: dataIn2 = 32'd1; 
32'd8229: dataIn2 = 32'd1; 
32'd8230: dataIn2 = 32'd0; 
32'd8231: dataIn2 = 32'd0; 
32'd8232: dataIn2 = 32'd0; 
32'd8233: dataIn2 = 32'd1; 
32'd8234: dataIn2 = 32'd1; 
32'd8235: dataIn2 = 32'd0; 
32'd8236: dataIn2 = 32'd0; 
32'd8237: dataIn2 = 32'd0; 
32'd8238: dataIn2 = 32'd1; 
32'd8239: dataIn2 = 32'd0; 
32'd8240: dataIn2 = 32'd0; 
32'd8241: dataIn2 = 32'd1; 
32'd8242: dataIn2 = 32'd0; 
32'd8243: dataIn2 = 32'd0; 
32'd8244: dataIn2 = 32'd1; 
32'd8245: dataIn2 = 32'd0; 
32'd8246: dataIn2 = 32'd0; 
32'd8247: dataIn2 = 32'd0; 
32'd8248: dataIn2 = 32'd1; 
32'd8249: dataIn2 = 32'd1; 
32'd8250: dataIn2 = 32'd0; 
32'd8251: dataIn2 = 32'd1; 
32'd8252: dataIn2 = 32'd0; 
32'd8253: dataIn2 = 32'd0; 
32'd8254: dataIn2 = 32'd0; 
32'd8255: dataIn2 = 32'd0; 
32'd8256: dataIn2 = 32'd0; 
32'd8257: dataIn2 = 32'd1; 
32'd8258: dataIn2 = 32'd1; 
32'd8259: dataIn2 = 32'd0; 
32'd8260: dataIn2 = 32'd1; 
32'd8261: dataIn2 = 32'd1; 
32'd8262: dataIn2 = 32'd0; 
32'd8263: dataIn2 = 32'd1; 
32'd8264: dataIn2 = 32'd0; 
32'd8265: dataIn2 = 32'd0; 
32'd8266: dataIn2 = 32'd1; 
32'd8267: dataIn2 = 32'd0; 
32'd8268: dataIn2 = 32'd0; 
32'd8269: dataIn2 = 32'd1; 
32'd8270: dataIn2 = 32'd0; 
32'd8271: dataIn2 = 32'd1; 
32'd8272: dataIn2 = 32'd1; 
32'd8273: dataIn2 = 32'd0; 
32'd8274: dataIn2 = 32'd0; 
32'd8275: dataIn2 = 32'd0; 
32'd8276: dataIn2 = 32'd1; 
32'd8277: dataIn2 = 32'd0; 
32'd8278: dataIn2 = 32'd0; 
32'd8279: dataIn2 = 32'd0; 
32'd8280: dataIn2 = 32'd0; 
32'd8281: dataIn2 = 32'd0; 
32'd8282: dataIn2 = 32'd1; 
32'd8283: dataIn2 = 32'd0; 
32'd8284: dataIn2 = 32'd0; 
32'd8285: dataIn2 = 32'd1; 
32'd8286: dataIn2 = 32'd1; 
32'd8287: dataIn2 = 32'd0; 
32'd8288: dataIn2 = 32'd1; 
32'd8289: dataIn2 = 32'd1; 
32'd8290: dataIn2 = 32'd0; 
32'd8291: dataIn2 = 32'd0; 
32'd8292: dataIn2 = 32'd1; 
32'd8293: dataIn2 = 32'd1; 
32'd8294: dataIn2 = 32'd1; 
32'd8295: dataIn2 = 32'd0; 
32'd8296: dataIn2 = 32'd0; 
32'd8297: dataIn2 = 32'd0; 
32'd8298: dataIn2 = 32'd0; 
32'd8299: dataIn2 = 32'd0; 
32'd8300: dataIn2 = 32'd1; 
32'd8301: dataIn2 = 32'd1; 
32'd8302: dataIn2 = 32'd0; 
32'd8303: dataIn2 = 32'd0; 
32'd8304: dataIn2 = 32'd1; 
32'd8305: dataIn2 = 32'd1; 
32'd8306: dataIn2 = 32'd0; 
32'd8307: dataIn2 = 32'd0; 
32'd8308: dataIn2 = 32'd0; 
32'd8309: dataIn2 = 32'd1; 
32'd8310: dataIn2 = 32'd0; 
32'd8311: dataIn2 = 32'd1; 
32'd8312: dataIn2 = 32'd0; 
32'd8313: dataIn2 = 32'd1; 
32'd8314: dataIn2 = 32'd1; 
32'd8315: dataIn2 = 32'd0; 
32'd8316: dataIn2 = 32'd1; 
32'd8317: dataIn2 = 32'd0; 
32'd8318: dataIn2 = 32'd1; 
32'd8319: dataIn2 = 32'd1; 
32'd8320: dataIn2 = 32'd1; 
32'd8321: dataIn2 = 32'd1; 
32'd8322: dataIn2 = 32'd0; 
32'd8323: dataIn2 = 32'd1; 
32'd8324: dataIn2 = 32'd1; 
32'd8325: dataIn2 = 32'd0; 
32'd8326: dataIn2 = 32'd0; 
32'd8327: dataIn2 = 32'd0; 
32'd8328: dataIn2 = 32'd0; 
32'd8329: dataIn2 = 32'd0; 
32'd8330: dataIn2 = 32'd1; 
32'd8331: dataIn2 = 32'd1; 
32'd8332: dataIn2 = 32'd1; 
32'd8333: dataIn2 = 32'd1; 
32'd8334: dataIn2 = 32'd1; 
32'd8335: dataIn2 = 32'd0; 
32'd8336: dataIn2 = 32'd0; 
32'd8337: dataIn2 = 32'd1; 
32'd8338: dataIn2 = 32'd0; 
32'd8339: dataIn2 = 32'd1; 
32'd8340: dataIn2 = 32'd0; 
32'd8341: dataIn2 = 32'd1; 
32'd8342: dataIn2 = 32'd0; 
32'd8343: dataIn2 = 32'd1; 
32'd8344: dataIn2 = 32'd1; 
32'd8345: dataIn2 = 32'd1; 
32'd8346: dataIn2 = 32'd0; 
32'd8347: dataIn2 = 32'd1; 
32'd8348: dataIn2 = 32'd1; 
32'd8349: dataIn2 = 32'd1; 
32'd8350: dataIn2 = 32'd1; 
32'd8351: dataIn2 = 32'd0; 
32'd8352: dataIn2 = 32'd0; 
32'd8353: dataIn2 = 32'd0; 
32'd8354: dataIn2 = 32'd0; 
32'd8355: dataIn2 = 32'd0; 
32'd8356: dataIn2 = 32'd1; 
32'd8357: dataIn2 = 32'd1; 
32'd8358: dataIn2 = 32'd1; 
32'd8359: dataIn2 = 32'd0; 
32'd8360: dataIn2 = 32'd1; 
32'd8361: dataIn2 = 32'd1; 
32'd8362: dataIn2 = 32'd0; 
32'd8363: dataIn2 = 32'd0; 
32'd8364: dataIn2 = 32'd1; 
32'd8365: dataIn2 = 32'd1; 
32'd8366: dataIn2 = 32'd1; 
32'd8367: dataIn2 = 32'd0; 
32'd8368: dataIn2 = 32'd0; 
32'd8369: dataIn2 = 32'd0; 
32'd8370: dataIn2 = 32'd0; 
32'd8371: dataIn2 = 32'd1; 
32'd8372: dataIn2 = 32'd1; 
32'd8373: dataIn2 = 32'd0; 
32'd8374: dataIn2 = 32'd0; 
32'd8375: dataIn2 = 32'd0; 
32'd8376: dataIn2 = 32'd1; 
32'd8377: dataIn2 = 32'd1; 
32'd8378: dataIn2 = 32'd0; 
32'd8379: dataIn2 = 32'd1; 
32'd8380: dataIn2 = 32'd1; 
32'd8381: dataIn2 = 32'd0; 
32'd8382: dataIn2 = 32'd0; 
32'd8383: dataIn2 = 32'd1; 
32'd8384: dataIn2 = 32'd0; 
32'd8385: dataIn2 = 32'd1; 
32'd8386: dataIn2 = 32'd1; 
32'd8387: dataIn2 = 32'd0; 
32'd8388: dataIn2 = 32'd0; 
32'd8389: dataIn2 = 32'd0; 
32'd8390: dataIn2 = 32'd0; 
32'd8391: dataIn2 = 32'd0; 
32'd8392: dataIn2 = 32'd1; 
32'd8393: dataIn2 = 32'd1; 
32'd8394: dataIn2 = 32'd1; 
32'd8395: dataIn2 = 32'd0; 
32'd8396: dataIn2 = 32'd1; 
32'd8397: dataIn2 = 32'd1; 
32'd8398: dataIn2 = 32'd1; 
32'd8399: dataIn2 = 32'd0; 
32'd8400: dataIn2 = 32'd0; 
32'd8401: dataIn2 = 32'd1; 
32'd8402: dataIn2 = 32'd1; 
32'd8403: dataIn2 = 32'd1; 
32'd8404: dataIn2 = 32'd1; 
32'd8405: dataIn2 = 32'd0; 
32'd8406: dataIn2 = 32'd0; 
32'd8407: dataIn2 = 32'd0; 
32'd8408: dataIn2 = 32'd1; 
32'd8409: dataIn2 = 32'd0; 
32'd8410: dataIn2 = 32'd0; 
32'd8411: dataIn2 = 32'd0; 
32'd8412: dataIn2 = 32'd1; 
32'd8413: dataIn2 = 32'd1; 
32'd8414: dataIn2 = 32'd0; 
32'd8415: dataIn2 = 32'd1; 
32'd8416: dataIn2 = 32'd0; 
32'd8417: dataIn2 = 32'd0; 
32'd8418: dataIn2 = 32'd0; 
32'd8419: dataIn2 = 32'd1; 
32'd8420: dataIn2 = 32'd0; 
32'd8421: dataIn2 = 32'd0; 
32'd8422: dataIn2 = 32'd1; 
32'd8423: dataIn2 = 32'd1; 
32'd8424: dataIn2 = 32'd0; 
32'd8425: dataIn2 = 32'd0; 
32'd8426: dataIn2 = 32'd0; 
32'd8427: dataIn2 = 32'd0; 
32'd8428: dataIn2 = 32'd0; 
32'd8429: dataIn2 = 32'd0; 
32'd8430: dataIn2 = 32'd1; 
32'd8431: dataIn2 = 32'd1; 
32'd8432: dataIn2 = 32'd1; 
32'd8433: dataIn2 = 32'd1; 
32'd8434: dataIn2 = 32'd1; 
32'd8435: dataIn2 = 32'd0; 
32'd8436: dataIn2 = 32'd0; 
32'd8437: dataIn2 = 32'd0; 
32'd8438: dataIn2 = 32'd1; 
32'd8439: dataIn2 = 32'd1; 
32'd8440: dataIn2 = 32'd1; 
32'd8441: dataIn2 = 32'd1; 
32'd8442: dataIn2 = 32'd0; 
32'd8443: dataIn2 = 32'd0; 
32'd8444: dataIn2 = 32'd0; 
32'd8445: dataIn2 = 32'd0; 
32'd8446: dataIn2 = 32'd1; 
32'd8447: dataIn2 = 32'd1; 
32'd8448: dataIn2 = 32'd0; 
32'd8449: dataIn2 = 32'd1; 
32'd8450: dataIn2 = 32'd0; 
32'd8451: dataIn2 = 32'd0; 
32'd8452: dataIn2 = 32'd1; 
32'd8453: dataIn2 = 32'd1; 
32'd8454: dataIn2 = 32'd0; 
32'd8455: dataIn2 = 32'd0; 
32'd8456: dataIn2 = 32'd0; 
32'd8457: dataIn2 = 32'd0; 
32'd8458: dataIn2 = 32'd0; 
32'd8459: dataIn2 = 32'd0; 
32'd8460: dataIn2 = 32'd0; 
32'd8461: dataIn2 = 32'd1; 
32'd8462: dataIn2 = 32'd1; 
32'd8463: dataIn2 = 32'd1; 
32'd8464: dataIn2 = 32'd1; 
32'd8465: dataIn2 = 32'd0; 
32'd8466: dataIn2 = 32'd0; 
32'd8467: dataIn2 = 32'd1; 
32'd8468: dataIn2 = 32'd0; 
32'd8469: dataIn2 = 32'd0; 
32'd8470: dataIn2 = 32'd0; 
32'd8471: dataIn2 = 32'd1; 
32'd8472: dataIn2 = 32'd0; 
32'd8473: dataIn2 = 32'd1; 
32'd8474: dataIn2 = 32'd1; 
32'd8475: dataIn2 = 32'd0; 
32'd8476: dataIn2 = 32'd0; 
32'd8477: dataIn2 = 32'd1; 
32'd8478: dataIn2 = 32'd0; 
32'd8479: dataIn2 = 32'd1; 
32'd8480: dataIn2 = 32'd1; 
32'd8481: dataIn2 = 32'd1; 
32'd8482: dataIn2 = 32'd0; 
32'd8483: dataIn2 = 32'd1; 
32'd8484: dataIn2 = 32'd1; 
32'd8485: dataIn2 = 32'd0; 
32'd8486: dataIn2 = 32'd1; 
32'd8487: dataIn2 = 32'd1; 
32'd8488: dataIn2 = 32'd0; 
32'd8489: dataIn2 = 32'd1; 
32'd8490: dataIn2 = 32'd1; 
32'd8491: dataIn2 = 32'd0; 
32'd8492: dataIn2 = 32'd0; 
32'd8493: dataIn2 = 32'd0; 
32'd8494: dataIn2 = 32'd0; 
32'd8495: dataIn2 = 32'd0; 
32'd8496: dataIn2 = 32'd0; 
32'd8497: dataIn2 = 32'd1; 
32'd8498: dataIn2 = 32'd0; 
32'd8499: dataIn2 = 32'd0; 
32'd8500: dataIn2 = 32'd0; 
32'd8501: dataIn2 = 32'd1; 
32'd8502: dataIn2 = 32'd0; 
32'd8503: dataIn2 = 32'd1; 
32'd8504: dataIn2 = 32'd1; 
32'd8505: dataIn2 = 32'd0; 
32'd8506: dataIn2 = 32'd1; 
32'd8507: dataIn2 = 32'd1; 
32'd8508: dataIn2 = 32'd0; 
32'd8509: dataIn2 = 32'd1; 
32'd8510: dataIn2 = 32'd0; 
32'd8511: dataIn2 = 32'd1; 
32'd8512: dataIn2 = 32'd0; 
32'd8513: dataIn2 = 32'd1; 
32'd8514: dataIn2 = 32'd0; 
32'd8515: dataIn2 = 32'd1; 
32'd8516: dataIn2 = 32'd0; 
32'd8517: dataIn2 = 32'd0; 
32'd8518: dataIn2 = 32'd0; 
32'd8519: dataIn2 = 32'd1; 
32'd8520: dataIn2 = 32'd1; 
32'd8521: dataIn2 = 32'd1; 
32'd8522: dataIn2 = 32'd0; 
32'd8523: dataIn2 = 32'd1; 
32'd8524: dataIn2 = 32'd1; 
32'd8525: dataIn2 = 32'd0; 
32'd8526: dataIn2 = 32'd0; 
32'd8527: dataIn2 = 32'd0; 
32'd8528: dataIn2 = 32'd0; 
32'd8529: dataIn2 = 32'd1; 
32'd8530: dataIn2 = 32'd0; 
32'd8531: dataIn2 = 32'd0; 
32'd8532: dataIn2 = 32'd1; 
32'd8533: dataIn2 = 32'd0; 
32'd8534: dataIn2 = 32'd0; 
32'd8535: dataIn2 = 32'd1; 
32'd8536: dataIn2 = 32'd0; 
32'd8537: dataIn2 = 32'd0; 
32'd8538: dataIn2 = 32'd0; 
32'd8539: dataIn2 = 32'd1; 
32'd8540: dataIn2 = 32'd0; 
32'd8541: dataIn2 = 32'd0; 
32'd8542: dataIn2 = 32'd0; 
32'd8543: dataIn2 = 32'd1; 
32'd8544: dataIn2 = 32'd0; 
32'd8545: dataIn2 = 32'd1; 
32'd8546: dataIn2 = 32'd0; 
32'd8547: dataIn2 = 32'd0; 
32'd8548: dataIn2 = 32'd1; 
32'd8549: dataIn2 = 32'd1; 
32'd8550: dataIn2 = 32'd0; 
32'd8551: dataIn2 = 32'd1; 
32'd8552: dataIn2 = 32'd0; 
32'd8553: dataIn2 = 32'd0; 
32'd8554: dataIn2 = 32'd0; 
32'd8555: dataIn2 = 32'd0; 
32'd8556: dataIn2 = 32'd0; 
32'd8557: dataIn2 = 32'd0; 
32'd8558: dataIn2 = 32'd1; 
32'd8559: dataIn2 = 32'd1; 
32'd8560: dataIn2 = 32'd0; 
32'd8561: dataIn2 = 32'd0; 
32'd8562: dataIn2 = 32'd1; 
32'd8563: dataIn2 = 32'd0; 
32'd8564: dataIn2 = 32'd1; 
32'd8565: dataIn2 = 32'd0; 
32'd8566: dataIn2 = 32'd1; 
32'd8567: dataIn2 = 32'd1; 
32'd8568: dataIn2 = 32'd1; 
32'd8569: dataIn2 = 32'd1; 
32'd8570: dataIn2 = 32'd1; 
32'd8571: dataIn2 = 32'd1; 
32'd8572: dataIn2 = 32'd1; 
32'd8573: dataIn2 = 32'd0; 
32'd8574: dataIn2 = 32'd1; 
32'd8575: dataIn2 = 32'd0; 
32'd8576: dataIn2 = 32'd1; 
32'd8577: dataIn2 = 32'd1; 
32'd8578: dataIn2 = 32'd0; 
32'd8579: dataIn2 = 32'd0; 
32'd8580: dataIn2 = 32'd1; 
32'd8581: dataIn2 = 32'd0; 
32'd8582: dataIn2 = 32'd1; 
32'd8583: dataIn2 = 32'd0; 
32'd8584: dataIn2 = 32'd0; 
32'd8585: dataIn2 = 32'd0; 
32'd8586: dataIn2 = 32'd1; 
32'd8587: dataIn2 = 32'd1; 
32'd8588: dataIn2 = 32'd1; 
32'd8589: dataIn2 = 32'd1; 
32'd8590: dataIn2 = 32'd1; 
32'd8591: dataIn2 = 32'd0; 
32'd8592: dataIn2 = 32'd1; 
32'd8593: dataIn2 = 32'd1; 
32'd8594: dataIn2 = 32'd0; 
32'd8595: dataIn2 = 32'd1; 
32'd8596: dataIn2 = 32'd0; 
32'd8597: dataIn2 = 32'd1; 
32'd8598: dataIn2 = 32'd0; 
32'd8599: dataIn2 = 32'd1; 
32'd8600: dataIn2 = 32'd1; 
32'd8601: dataIn2 = 32'd0; 
32'd8602: dataIn2 = 32'd0; 
32'd8603: dataIn2 = 32'd1; 
32'd8604: dataIn2 = 32'd1; 
32'd8605: dataIn2 = 32'd0; 
32'd8606: dataIn2 = 32'd1; 
32'd8607: dataIn2 = 32'd0; 
32'd8608: dataIn2 = 32'd1; 
32'd8609: dataIn2 = 32'd0; 
32'd8610: dataIn2 = 32'd0; 
32'd8611: dataIn2 = 32'd0; 
32'd8612: dataIn2 = 32'd1; 
32'd8613: dataIn2 = 32'd0; 
32'd8614: dataIn2 = 32'd0; 
32'd8615: dataIn2 = 32'd1; 
32'd8616: dataIn2 = 32'd0; 
32'd8617: dataIn2 = 32'd1; 
32'd8618: dataIn2 = 32'd0; 
32'd8619: dataIn2 = 32'd1; 
32'd8620: dataIn2 = 32'd1; 
32'd8621: dataIn2 = 32'd0; 
32'd8622: dataIn2 = 32'd0; 
32'd8623: dataIn2 = 32'd1; 
32'd8624: dataIn2 = 32'd1; 
32'd8625: dataIn2 = 32'd0; 
32'd8626: dataIn2 = 32'd0; 
32'd8627: dataIn2 = 32'd1; 
32'd8628: dataIn2 = 32'd0; 
32'd8629: dataIn2 = 32'd1; 
32'd8630: dataIn2 = 32'd1; 
32'd8631: dataIn2 = 32'd1; 
32'd8632: dataIn2 = 32'd0; 
32'd8633: dataIn2 = 32'd0; 
32'd8634: dataIn2 = 32'd0; 
32'd8635: dataIn2 = 32'd1; 
32'd8636: dataIn2 = 32'd0; 
32'd8637: dataIn2 = 32'd1; 
32'd8638: dataIn2 = 32'd1; 
32'd8639: dataIn2 = 32'd1; 
32'd8640: dataIn2 = 32'd1; 
32'd8641: dataIn2 = 32'd0; 
32'd8642: dataIn2 = 32'd0; 
32'd8643: dataIn2 = 32'd1; 
32'd8644: dataIn2 = 32'd0; 
32'd8645: dataIn2 = 32'd0; 
32'd8646: dataIn2 = 32'd1; 
32'd8647: dataIn2 = 32'd0; 
32'd8648: dataIn2 = 32'd0; 
32'd8649: dataIn2 = 32'd0; 
32'd8650: dataIn2 = 32'd0; 
32'd8651: dataIn2 = 32'd0; 
32'd8652: dataIn2 = 32'd0; 
32'd8653: dataIn2 = 32'd1; 
32'd8654: dataIn2 = 32'd0; 
32'd8655: dataIn2 = 32'd0; 
32'd8656: dataIn2 = 32'd0; 
32'd8657: dataIn2 = 32'd1; 
32'd8658: dataIn2 = 32'd0; 
32'd8659: dataIn2 = 32'd0; 
32'd8660: dataIn2 = 32'd0; 
32'd8661: dataIn2 = 32'd1; 
32'd8662: dataIn2 = 32'd1; 
32'd8663: dataIn2 = 32'd0; 
32'd8664: dataIn2 = 32'd1; 
32'd8665: dataIn2 = 32'd0; 
32'd8666: dataIn2 = 32'd1; 
32'd8667: dataIn2 = 32'd1; 
32'd8668: dataIn2 = 32'd1; 
32'd8669: dataIn2 = 32'd0; 
32'd8670: dataIn2 = 32'd0; 
32'd8671: dataIn2 = 32'd0; 
32'd8672: dataIn2 = 32'd0; 
32'd8673: dataIn2 = 32'd1; 
32'd8674: dataIn2 = 32'd0; 
32'd8675: dataIn2 = 32'd1; 
32'd8676: dataIn2 = 32'd0; 
32'd8677: dataIn2 = 32'd1; 
32'd8678: dataIn2 = 32'd0; 
32'd8679: dataIn2 = 32'd1; 
32'd8680: dataIn2 = 32'd0; 
32'd8681: dataIn2 = 32'd1; 
32'd8682: dataIn2 = 32'd1; 
32'd8683: dataIn2 = 32'd0; 
32'd8684: dataIn2 = 32'd1; 
32'd8685: dataIn2 = 32'd0; 
32'd8686: dataIn2 = 32'd1; 
32'd8687: dataIn2 = 32'd1; 
32'd8688: dataIn2 = 32'd1; 
32'd8689: dataIn2 = 32'd0; 
32'd8690: dataIn2 = 32'd0; 
32'd8691: dataIn2 = 32'd0; 
32'd8692: dataIn2 = 32'd0; 
32'd8693: dataIn2 = 32'd1; 
32'd8694: dataIn2 = 32'd0; 
32'd8695: dataIn2 = 32'd0; 
32'd8696: dataIn2 = 32'd1; 
32'd8697: dataIn2 = 32'd1; 
32'd8698: dataIn2 = 32'd1; 
32'd8699: dataIn2 = 32'd0; 
32'd8700: dataIn2 = 32'd1; 
32'd8701: dataIn2 = 32'd0; 
32'd8702: dataIn2 = 32'd0; 
32'd8703: dataIn2 = 32'd1; 
32'd8704: dataIn2 = 32'd0; 
32'd8705: dataIn2 = 32'd0; 
32'd8706: dataIn2 = 32'd1; 
32'd8707: dataIn2 = 32'd1; 
32'd8708: dataIn2 = 32'd1; 
32'd8709: dataIn2 = 32'd0; 
32'd8710: dataIn2 = 32'd0; 
32'd8711: dataIn2 = 32'd0; 
32'd8712: dataIn2 = 32'd1; 
32'd8713: dataIn2 = 32'd0; 
32'd8714: dataIn2 = 32'd0; 
32'd8715: dataIn2 = 32'd0; 
32'd8716: dataIn2 = 32'd1; 
32'd8717: dataIn2 = 32'd0; 
32'd8718: dataIn2 = 32'd0; 
32'd8719: dataIn2 = 32'd0; 
32'd8720: dataIn2 = 32'd1; 
32'd8721: dataIn2 = 32'd0; 
32'd8722: dataIn2 = 32'd1; 
32'd8723: dataIn2 = 32'd1; 
32'd8724: dataIn2 = 32'd1; 
32'd8725: dataIn2 = 32'd1; 
32'd8726: dataIn2 = 32'd0; 
32'd8727: dataIn2 = 32'd1; 
32'd8728: dataIn2 = 32'd0; 
32'd8729: dataIn2 = 32'd0; 
32'd8730: dataIn2 = 32'd1; 
32'd8731: dataIn2 = 32'd0; 
32'd8732: dataIn2 = 32'd1; 
32'd8733: dataIn2 = 32'd0; 
32'd8734: dataIn2 = 32'd1; 
32'd8735: dataIn2 = 32'd0; 
32'd8736: dataIn2 = 32'd1; 
32'd8737: dataIn2 = 32'd1; 
32'd8738: dataIn2 = 32'd1; 
32'd8739: dataIn2 = 32'd1; 
32'd8740: dataIn2 = 32'd0; 
32'd8741: dataIn2 = 32'd0; 
32'd8742: dataIn2 = 32'd1; 
32'd8743: dataIn2 = 32'd1; 
32'd8744: dataIn2 = 32'd1; 
32'd8745: dataIn2 = 32'd1; 
32'd8746: dataIn2 = 32'd1; 
32'd8747: dataIn2 = 32'd0; 
32'd8748: dataIn2 = 32'd0; 
32'd8749: dataIn2 = 32'd0; 
32'd8750: dataIn2 = 32'd1; 
32'd8751: dataIn2 = 32'd0; 
32'd8752: dataIn2 = 32'd1; 
32'd8753: dataIn2 = 32'd0; 
32'd8754: dataIn2 = 32'd0; 
32'd8755: dataIn2 = 32'd0; 
32'd8756: dataIn2 = 32'd1; 
32'd8757: dataIn2 = 32'd0; 
32'd8758: dataIn2 = 32'd0; 
32'd8759: dataIn2 = 32'd1; 
32'd8760: dataIn2 = 32'd0; 
32'd8761: dataIn2 = 32'd1; 
32'd8762: dataIn2 = 32'd0; 
32'd8763: dataIn2 = 32'd1; 
32'd8764: dataIn2 = 32'd1; 
32'd8765: dataIn2 = 32'd0; 
32'd8766: dataIn2 = 32'd0; 
32'd8767: dataIn2 = 32'd0; 
32'd8768: dataIn2 = 32'd0; 
32'd8769: dataIn2 = 32'd1; 
32'd8770: dataIn2 = 32'd1; 
32'd8771: dataIn2 = 32'd0; 
32'd8772: dataIn2 = 32'd0; 
32'd8773: dataIn2 = 32'd0; 
32'd8774: dataIn2 = 32'd0; 
32'd8775: dataIn2 = 32'd1; 
32'd8776: dataIn2 = 32'd1; 
32'd8777: dataIn2 = 32'd0; 
32'd8778: dataIn2 = 32'd1; 
32'd8779: dataIn2 = 32'd0; 
32'd8780: dataIn2 = 32'd0; 
32'd8781: dataIn2 = 32'd0; 
32'd8782: dataIn2 = 32'd1; 
32'd8783: dataIn2 = 32'd1; 
32'd8784: dataIn2 = 32'd0; 
32'd8785: dataIn2 = 32'd1; 
32'd8786: dataIn2 = 32'd0; 
32'd8787: dataIn2 = 32'd1; 
32'd8788: dataIn2 = 32'd0; 
32'd8789: dataIn2 = 32'd1; 
32'd8790: dataIn2 = 32'd1; 
32'd8791: dataIn2 = 32'd0; 
32'd8792: dataIn2 = 32'd0; 
32'd8793: dataIn2 = 32'd0; 
32'd8794: dataIn2 = 32'd0; 
32'd8795: dataIn2 = 32'd1; 
32'd8796: dataIn2 = 32'd1; 
32'd8797: dataIn2 = 32'd1; 
32'd8798: dataIn2 = 32'd1; 
32'd8799: dataIn2 = 32'd0; 
32'd8800: dataIn2 = 32'd1; 
32'd8801: dataIn2 = 32'd1; 
32'd8802: dataIn2 = 32'd0; 
32'd8803: dataIn2 = 32'd0; 
32'd8804: dataIn2 = 32'd0; 
32'd8805: dataIn2 = 32'd1; 
32'd8806: dataIn2 = 32'd0; 
32'd8807: dataIn2 = 32'd1; 
32'd8808: dataIn2 = 32'd1; 
32'd8809: dataIn2 = 32'd0; 
32'd8810: dataIn2 = 32'd1; 
32'd8811: dataIn2 = 32'd1; 
32'd8812: dataIn2 = 32'd1; 
32'd8813: dataIn2 = 32'd1; 
32'd8814: dataIn2 = 32'd0; 
32'd8815: dataIn2 = 32'd1; 
32'd8816: dataIn2 = 32'd0; 
32'd8817: dataIn2 = 32'd1; 
32'd8818: dataIn2 = 32'd0; 
32'd8819: dataIn2 = 32'd1; 
32'd8820: dataIn2 = 32'd0; 
32'd8821: dataIn2 = 32'd1; 
32'd8822: dataIn2 = 32'd1; 
32'd8823: dataIn2 = 32'd0; 
32'd8824: dataIn2 = 32'd1; 
32'd8825: dataIn2 = 32'd1; 
32'd8826: dataIn2 = 32'd0; 
32'd8827: dataIn2 = 32'd0; 
32'd8828: dataIn2 = 32'd1; 
32'd8829: dataIn2 = 32'd0; 
32'd8830: dataIn2 = 32'd0; 
32'd8831: dataIn2 = 32'd1; 
32'd8832: dataIn2 = 32'd0; 
32'd8833: dataIn2 = 32'd1; 
32'd8834: dataIn2 = 32'd1; 
32'd8835: dataIn2 = 32'd0; 
32'd8836: dataIn2 = 32'd0; 
32'd8837: dataIn2 = 32'd0; 
32'd8838: dataIn2 = 32'd1; 
32'd8839: dataIn2 = 32'd0; 
32'd8840: dataIn2 = 32'd0; 
32'd8841: dataIn2 = 32'd0; 
32'd8842: dataIn2 = 32'd0; 
32'd8843: dataIn2 = 32'd1; 
32'd8844: dataIn2 = 32'd0; 
32'd8845: dataIn2 = 32'd1; 
32'd8846: dataIn2 = 32'd0; 
32'd8847: dataIn2 = 32'd1; 
32'd8848: dataIn2 = 32'd0; 
32'd8849: dataIn2 = 32'd0; 
32'd8850: dataIn2 = 32'd0; 
32'd8851: dataIn2 = 32'd1; 
32'd8852: dataIn2 = 32'd1; 
32'd8853: dataIn2 = 32'd0; 
32'd8854: dataIn2 = 32'd0; 
32'd8855: dataIn2 = 32'd1; 
32'd8856: dataIn2 = 32'd1; 
32'd8857: dataIn2 = 32'd0; 
32'd8858: dataIn2 = 32'd0; 
32'd8859: dataIn2 = 32'd1; 
32'd8860: dataIn2 = 32'd1; 
32'd8861: dataIn2 = 32'd1; 
32'd8862: dataIn2 = 32'd0; 
32'd8863: dataIn2 = 32'd0; 
32'd8864: dataIn2 = 32'd0; 
32'd8865: dataIn2 = 32'd1; 
32'd8866: dataIn2 = 32'd0; 
32'd8867: dataIn2 = 32'd0; 
32'd8868: dataIn2 = 32'd1; 
32'd8869: dataIn2 = 32'd1; 
32'd8870: dataIn2 = 32'd1; 
32'd8871: dataIn2 = 32'd0; 
32'd8872: dataIn2 = 32'd1; 
32'd8873: dataIn2 = 32'd1; 
32'd8874: dataIn2 = 32'd0; 
32'd8875: dataIn2 = 32'd1; 
32'd8876: dataIn2 = 32'd0; 
32'd8877: dataIn2 = 32'd0; 
32'd8878: dataIn2 = 32'd1; 
32'd8879: dataIn2 = 32'd0; 
32'd8880: dataIn2 = 32'd0; 
32'd8881: dataIn2 = 32'd1; 
32'd8882: dataIn2 = 32'd0; 
32'd8883: dataIn2 = 32'd0; 
32'd8884: dataIn2 = 32'd0; 
32'd8885: dataIn2 = 32'd0; 
32'd8886: dataIn2 = 32'd1; 
32'd8887: dataIn2 = 32'd1; 
32'd8888: dataIn2 = 32'd1; 
32'd8889: dataIn2 = 32'd0; 
32'd8890: dataIn2 = 32'd0; 
32'd8891: dataIn2 = 32'd0; 
32'd8892: dataIn2 = 32'd1; 
32'd8893: dataIn2 = 32'd1; 
32'd8894: dataIn2 = 32'd1; 
32'd8895: dataIn2 = 32'd0; 
32'd8896: dataIn2 = 32'd0; 
32'd8897: dataIn2 = 32'd0; 
32'd8898: dataIn2 = 32'd1; 
32'd8899: dataIn2 = 32'd0; 
32'd8900: dataIn2 = 32'd0; 
32'd8901: dataIn2 = 32'd1; 
32'd8902: dataIn2 = 32'd1; 
32'd8903: dataIn2 = 32'd0; 
32'd8904: dataIn2 = 32'd1; 
32'd8905: dataIn2 = 32'd1; 
32'd8906: dataIn2 = 32'd0; 
32'd8907: dataIn2 = 32'd1; 
32'd8908: dataIn2 = 32'd0; 
32'd8909: dataIn2 = 32'd0; 
32'd8910: dataIn2 = 32'd1; 
32'd8911: dataIn2 = 32'd0; 
32'd8912: dataIn2 = 32'd0; 
32'd8913: dataIn2 = 32'd0; 
32'd8914: dataIn2 = 32'd1; 
32'd8915: dataIn2 = 32'd1; 
32'd8916: dataIn2 = 32'd0; 
32'd8917: dataIn2 = 32'd0; 
32'd8918: dataIn2 = 32'd0; 
32'd8919: dataIn2 = 32'd1; 
32'd8920: dataIn2 = 32'd1; 
32'd8921: dataIn2 = 32'd1; 
32'd8922: dataIn2 = 32'd0; 
32'd8923: dataIn2 = 32'd1; 
32'd8924: dataIn2 = 32'd0; 
32'd8925: dataIn2 = 32'd1; 
32'd8926: dataIn2 = 32'd0; 
32'd8927: dataIn2 = 32'd1; 
32'd8928: dataIn2 = 32'd0; 
32'd8929: dataIn2 = 32'd1; 
32'd8930: dataIn2 = 32'd0; 
32'd8931: dataIn2 = 32'd1; 
32'd8932: dataIn2 = 32'd0; 
32'd8933: dataIn2 = 32'd0; 
32'd8934: dataIn2 = 32'd0; 
32'd8935: dataIn2 = 32'd0; 
32'd8936: dataIn2 = 32'd1; 
32'd8937: dataIn2 = 32'd0; 
32'd8938: dataIn2 = 32'd0; 
32'd8939: dataIn2 = 32'd1; 
32'd8940: dataIn2 = 32'd1; 
32'd8941: dataIn2 = 32'd1; 
32'd8942: dataIn2 = 32'd0; 
32'd8943: dataIn2 = 32'd0; 
32'd8944: dataIn2 = 32'd0; 
32'd8945: dataIn2 = 32'd1; 
32'd8946: dataIn2 = 32'd0; 
32'd8947: dataIn2 = 32'd0; 
32'd8948: dataIn2 = 32'd0; 
32'd8949: dataIn2 = 32'd0; 
32'd8950: dataIn2 = 32'd1; 
32'd8951: dataIn2 = 32'd1; 
32'd8952: dataIn2 = 32'd0; 
32'd8953: dataIn2 = 32'd1; 
32'd8954: dataIn2 = 32'd1; 
32'd8955: dataIn2 = 32'd0; 
32'd8956: dataIn2 = 32'd0; 
32'd8957: dataIn2 = 32'd0; 
32'd8958: dataIn2 = 32'd1; 
32'd8959: dataIn2 = 32'd0; 
32'd8960: dataIn2 = 32'd0; 
32'd8961: dataIn2 = 32'd0; 
32'd8962: dataIn2 = 32'd0; 
32'd8963: dataIn2 = 32'd0; 
32'd8964: dataIn2 = 32'd1; 
32'd8965: dataIn2 = 32'd1; 
32'd8966: dataIn2 = 32'd0; 
32'd8967: dataIn2 = 32'd0; 
32'd8968: dataIn2 = 32'd0; 
32'd8969: dataIn2 = 32'd1; 
32'd8970: dataIn2 = 32'd1; 
32'd8971: dataIn2 = 32'd0; 
32'd8972: dataIn2 = 32'd0; 
32'd8973: dataIn2 = 32'd0; 
32'd8974: dataIn2 = 32'd0; 
32'd8975: dataIn2 = 32'd1; 
32'd8976: dataIn2 = 32'd0; 
32'd8977: dataIn2 = 32'd0; 
32'd8978: dataIn2 = 32'd1; 
32'd8979: dataIn2 = 32'd0; 
32'd8980: dataIn2 = 32'd1; 
32'd8981: dataIn2 = 32'd1; 
32'd8982: dataIn2 = 32'd0; 
32'd8983: dataIn2 = 32'd1; 
32'd8984: dataIn2 = 32'd0; 
32'd8985: dataIn2 = 32'd1; 
32'd8986: dataIn2 = 32'd1; 
32'd8987: dataIn2 = 32'd0; 
32'd8988: dataIn2 = 32'd0; 
32'd8989: dataIn2 = 32'd1; 
32'd8990: dataIn2 = 32'd0; 
32'd8991: dataIn2 = 32'd1; 
32'd8992: dataIn2 = 32'd1; 
32'd8993: dataIn2 = 32'd0; 
32'd8994: dataIn2 = 32'd0; 
32'd8995: dataIn2 = 32'd1; 
32'd8996: dataIn2 = 32'd0; 
32'd8997: dataIn2 = 32'd1; 
32'd8998: dataIn2 = 32'd0; 
32'd8999: dataIn2 = 32'd1; 
32'd9000: dataIn2 = 32'd0; 
32'd9001: dataIn2 = 32'd1; 
32'd9002: dataIn2 = 32'd0; 
32'd9003: dataIn2 = 32'd1; 
32'd9004: dataIn2 = 32'd0; 
32'd9005: dataIn2 = 32'd1; 
32'd9006: dataIn2 = 32'd1; 
32'd9007: dataIn2 = 32'd1; 
32'd9008: dataIn2 = 32'd0; 
32'd9009: dataIn2 = 32'd0; 
32'd9010: dataIn2 = 32'd1; 
32'd9011: dataIn2 = 32'd0; 
32'd9012: dataIn2 = 32'd1; 
32'd9013: dataIn2 = 32'd0; 
32'd9014: dataIn2 = 32'd0; 
32'd9015: dataIn2 = 32'd1; 
32'd9016: dataIn2 = 32'd0; 
32'd9017: dataIn2 = 32'd0; 
32'd9018: dataIn2 = 32'd1; 
32'd9019: dataIn2 = 32'd0; 
32'd9020: dataIn2 = 32'd1; 
32'd9021: dataIn2 = 32'd1; 
32'd9022: dataIn2 = 32'd0; 
32'd9023: dataIn2 = 32'd1; 
32'd9024: dataIn2 = 32'd0; 
32'd9025: dataIn2 = 32'd0; 
32'd9026: dataIn2 = 32'd0; 
32'd9027: dataIn2 = 32'd1; 
32'd9028: dataIn2 = 32'd1; 
32'd9029: dataIn2 = 32'd0; 
32'd9030: dataIn2 = 32'd0; 
32'd9031: dataIn2 = 32'd0; 
32'd9032: dataIn2 = 32'd0; 
32'd9033: dataIn2 = 32'd1; 
32'd9034: dataIn2 = 32'd0; 
32'd9035: dataIn2 = 32'd1; 
32'd9036: dataIn2 = 32'd0; 
32'd9037: dataIn2 = 32'd0; 
32'd9038: dataIn2 = 32'd1; 
32'd9039: dataIn2 = 32'd1; 
32'd9040: dataIn2 = 32'd0; 
32'd9041: dataIn2 = 32'd0; 
32'd9042: dataIn2 = 32'd0; 
32'd9043: dataIn2 = 32'd0; 
32'd9044: dataIn2 = 32'd1; 
32'd9045: dataIn2 = 32'd1; 
32'd9046: dataIn2 = 32'd1; 
32'd9047: dataIn2 = 32'd0; 
32'd9048: dataIn2 = 32'd1; 
32'd9049: dataIn2 = 32'd1; 
32'd9050: dataIn2 = 32'd0; 
32'd9051: dataIn2 = 32'd1; 
32'd9052: dataIn2 = 32'd1; 
32'd9053: dataIn2 = 32'd0; 
32'd9054: dataIn2 = 32'd0; 
32'd9055: dataIn2 = 32'd0; 
32'd9056: dataIn2 = 32'd1; 
32'd9057: dataIn2 = 32'd1; 
32'd9058: dataIn2 = 32'd0; 
32'd9059: dataIn2 = 32'd0; 
32'd9060: dataIn2 = 32'd1; 
32'd9061: dataIn2 = 32'd0; 
32'd9062: dataIn2 = 32'd0; 
32'd9063: dataIn2 = 32'd1; 
32'd9064: dataIn2 = 32'd0; 
32'd9065: dataIn2 = 32'd0; 
32'd9066: dataIn2 = 32'd0; 
32'd9067: dataIn2 = 32'd1; 
32'd9068: dataIn2 = 32'd1; 
32'd9069: dataIn2 = 32'd1; 
32'd9070: dataIn2 = 32'd0; 
32'd9071: dataIn2 = 32'd0; 
32'd9072: dataIn2 = 32'd0; 
32'd9073: dataIn2 = 32'd1; 
32'd9074: dataIn2 = 32'd1; 
32'd9075: dataIn2 = 32'd0; 
32'd9076: dataIn2 = 32'd0; 
32'd9077: dataIn2 = 32'd0; 
32'd9078: dataIn2 = 32'd1; 
32'd9079: dataIn2 = 32'd1; 
32'd9080: dataIn2 = 32'd0; 
32'd9081: dataIn2 = 32'd1; 
32'd9082: dataIn2 = 32'd0; 
32'd9083: dataIn2 = 32'd1; 
32'd9084: dataIn2 = 32'd1; 
32'd9085: dataIn2 = 32'd1; 
32'd9086: dataIn2 = 32'd1; 
32'd9087: dataIn2 = 32'd0; 
32'd9088: dataIn2 = 32'd0; 
32'd9089: dataIn2 = 32'd1; 
32'd9090: dataIn2 = 32'd0; 
32'd9091: dataIn2 = 32'd0; 
32'd9092: dataIn2 = 32'd0; 
32'd9093: dataIn2 = 32'd0; 
32'd9094: dataIn2 = 32'd0; 
32'd9095: dataIn2 = 32'd1; 
32'd9096: dataIn2 = 32'd1; 
32'd9097: dataIn2 = 32'd1; 
32'd9098: dataIn2 = 32'd0; 
32'd9099: dataIn2 = 32'd1; 
32'd9100: dataIn2 = 32'd0; 
32'd9101: dataIn2 = 32'd0; 
32'd9102: dataIn2 = 32'd1; 
32'd9103: dataIn2 = 32'd0; 
32'd9104: dataIn2 = 32'd0; 
32'd9105: dataIn2 = 32'd1; 
32'd9106: dataIn2 = 32'd1; 
32'd9107: dataIn2 = 32'd1; 
32'd9108: dataIn2 = 32'd0; 
32'd9109: dataIn2 = 32'd0; 
32'd9110: dataIn2 = 32'd1; 
32'd9111: dataIn2 = 32'd0; 
32'd9112: dataIn2 = 32'd1; 
32'd9113: dataIn2 = 32'd1; 
32'd9114: dataIn2 = 32'd1; 
32'd9115: dataIn2 = 32'd0; 
32'd9116: dataIn2 = 32'd0; 
32'd9117: dataIn2 = 32'd0; 
32'd9118: dataIn2 = 32'd0; 
32'd9119: dataIn2 = 32'd0; 
32'd9120: dataIn2 = 32'd0; 
32'd9121: dataIn2 = 32'd1; 
32'd9122: dataIn2 = 32'd0; 
32'd9123: dataIn2 = 32'd0; 
32'd9124: dataIn2 = 32'd0; 
32'd9125: dataIn2 = 32'd1; 
32'd9126: dataIn2 = 32'd0; 
32'd9127: dataIn2 = 32'd1; 
32'd9128: dataIn2 = 32'd0; 
32'd9129: dataIn2 = 32'd1; 
32'd9130: dataIn2 = 32'd1; 
32'd9131: dataIn2 = 32'd0; 
32'd9132: dataIn2 = 32'd0; 
32'd9133: dataIn2 = 32'd0; 
32'd9134: dataIn2 = 32'd0; 
32'd9135: dataIn2 = 32'd0; 
32'd9136: dataIn2 = 32'd0; 
32'd9137: dataIn2 = 32'd0; 
32'd9138: dataIn2 = 32'd1; 
32'd9139: dataIn2 = 32'd1; 
32'd9140: dataIn2 = 32'd0; 
32'd9141: dataIn2 = 32'd0; 
32'd9142: dataIn2 = 32'd0; 
32'd9143: dataIn2 = 32'd1; 
32'd9144: dataIn2 = 32'd1; 
32'd9145: dataIn2 = 32'd1; 
32'd9146: dataIn2 = 32'd1; 
32'd9147: dataIn2 = 32'd1; 
32'd9148: dataIn2 = 32'd0; 
32'd9149: dataIn2 = 32'd0; 
32'd9150: dataIn2 = 32'd1; 
32'd9151: dataIn2 = 32'd0; 
32'd9152: dataIn2 = 32'd1; 
32'd9153: dataIn2 = 32'd1; 
32'd9154: dataIn2 = 32'd1; 
32'd9155: dataIn2 = 32'd1; 
32'd9156: dataIn2 = 32'd1; 
32'd9157: dataIn2 = 32'd0; 
32'd9158: dataIn2 = 32'd0; 
32'd9159: dataIn2 = 32'd1; 
32'd9160: dataIn2 = 32'd1; 
32'd9161: dataIn2 = 32'd1; 
32'd9162: dataIn2 = 32'd1; 
32'd9163: dataIn2 = 32'd0; 
32'd9164: dataIn2 = 32'd1; 
32'd9165: dataIn2 = 32'd1; 
32'd9166: dataIn2 = 32'd0; 
32'd9167: dataIn2 = 32'd0; 
32'd9168: dataIn2 = 32'd0; 
32'd9169: dataIn2 = 32'd1; 
32'd9170: dataIn2 = 32'd0; 
32'd9171: dataIn2 = 32'd0; 
32'd9172: dataIn2 = 32'd0; 
32'd9173: dataIn2 = 32'd1; 
32'd9174: dataIn2 = 32'd0; 
32'd9175: dataIn2 = 32'd1; 
32'd9176: dataIn2 = 32'd0; 
32'd9177: dataIn2 = 32'd1; 
32'd9178: dataIn2 = 32'd0; 
32'd9179: dataIn2 = 32'd0; 
32'd9180: dataIn2 = 32'd0; 
32'd9181: dataIn2 = 32'd1; 
32'd9182: dataIn2 = 32'd1; 
32'd9183: dataIn2 = 32'd0; 
32'd9184: dataIn2 = 32'd1; 
32'd9185: dataIn2 = 32'd1; 
32'd9186: dataIn2 = 32'd1; 
32'd9187: dataIn2 = 32'd1; 
32'd9188: dataIn2 = 32'd1; 
32'd9189: dataIn2 = 32'd0; 
32'd9190: dataIn2 = 32'd1; 
32'd9191: dataIn2 = 32'd0; 
32'd9192: dataIn2 = 32'd1; 
32'd9193: dataIn2 = 32'd0; 
32'd9194: dataIn2 = 32'd1; 
32'd9195: dataIn2 = 32'd0; 
32'd9196: dataIn2 = 32'd0; 
32'd9197: dataIn2 = 32'd0; 
32'd9198: dataIn2 = 32'd0; 
32'd9199: dataIn2 = 32'd1; 
32'd9200: dataIn2 = 32'd0; 
32'd9201: dataIn2 = 32'd0; 
32'd9202: dataIn2 = 32'd0; 
32'd9203: dataIn2 = 32'd0; 
32'd9204: dataIn2 = 32'd1; 
32'd9205: dataIn2 = 32'd1; 
32'd9206: dataIn2 = 32'd1; 
32'd9207: dataIn2 = 32'd0; 
32'd9208: dataIn2 = 32'd1; 
32'd9209: dataIn2 = 32'd0; 
32'd9210: dataIn2 = 32'd1; 
32'd9211: dataIn2 = 32'd0; 
32'd9212: dataIn2 = 32'd1; 
32'd9213: dataIn2 = 32'd0; 
32'd9214: dataIn2 = 32'd0; 
32'd9215: dataIn2 = 32'd1; 
32'd9216: dataIn2 = 32'd0; 
32'd9217: dataIn2 = 32'd0; 
32'd9218: dataIn2 = 32'd1; 
32'd9219: dataIn2 = 32'd1; 
32'd9220: dataIn2 = 32'd0; 
32'd9221: dataIn2 = 32'd0; 
32'd9222: dataIn2 = 32'd1; 
32'd9223: dataIn2 = 32'd0; 
32'd9224: dataIn2 = 32'd1; 
32'd9225: dataIn2 = 32'd1; 
32'd9226: dataIn2 = 32'd0; 
32'd9227: dataIn2 = 32'd0; 
32'd9228: dataIn2 = 32'd0; 
32'd9229: dataIn2 = 32'd1; 
32'd9230: dataIn2 = 32'd0; 
32'd9231: dataIn2 = 32'd1; 
32'd9232: dataIn2 = 32'd0; 
32'd9233: dataIn2 = 32'd1; 
32'd9234: dataIn2 = 32'd1; 
32'd9235: dataIn2 = 32'd0; 
32'd9236: dataIn2 = 32'd1; 
32'd9237: dataIn2 = 32'd1; 
32'd9238: dataIn2 = 32'd0; 
32'd9239: dataIn2 = 32'd1; 
32'd9240: dataIn2 = 32'd0; 
32'd9241: dataIn2 = 32'd1; 
32'd9242: dataIn2 = 32'd0; 
32'd9243: dataIn2 = 32'd1; 
32'd9244: dataIn2 = 32'd0; 
32'd9245: dataIn2 = 32'd0; 
32'd9246: dataIn2 = 32'd0; 
32'd9247: dataIn2 = 32'd1; 
32'd9248: dataIn2 = 32'd0; 
32'd9249: dataIn2 = 32'd1; 
32'd9250: dataIn2 = 32'd0; 
32'd9251: dataIn2 = 32'd0; 
32'd9252: dataIn2 = 32'd1; 
32'd9253: dataIn2 = 32'd0; 
32'd9254: dataIn2 = 32'd1; 
32'd9255: dataIn2 = 32'd0; 
32'd9256: dataIn2 = 32'd0; 
32'd9257: dataIn2 = 32'd1; 
32'd9258: dataIn2 = 32'd1; 
32'd9259: dataIn2 = 32'd0; 
32'd9260: dataIn2 = 32'd0; 
32'd9261: dataIn2 = 32'd0; 
32'd9262: dataIn2 = 32'd0; 
32'd9263: dataIn2 = 32'd1; 
32'd9264: dataIn2 = 32'd1; 
32'd9265: dataIn2 = 32'd1; 
32'd9266: dataIn2 = 32'd1; 
32'd9267: dataIn2 = 32'd1; 
32'd9268: dataIn2 = 32'd0; 
32'd9269: dataIn2 = 32'd1; 
32'd9270: dataIn2 = 32'd0; 
32'd9271: dataIn2 = 32'd1; 
32'd9272: dataIn2 = 32'd1; 
32'd9273: dataIn2 = 32'd0; 
32'd9274: dataIn2 = 32'd0; 
32'd9275: dataIn2 = 32'd1; 
32'd9276: dataIn2 = 32'd1; 
32'd9277: dataIn2 = 32'd1; 
32'd9278: dataIn2 = 32'd1; 
32'd9279: dataIn2 = 32'd0; 
32'd9280: dataIn2 = 32'd0; 
32'd9281: dataIn2 = 32'd0; 
32'd9282: dataIn2 = 32'd0; 
32'd9283: dataIn2 = 32'd0; 
32'd9284: dataIn2 = 32'd1; 
32'd9285: dataIn2 = 32'd0; 
32'd9286: dataIn2 = 32'd1; 
32'd9287: dataIn2 = 32'd0; 
32'd9288: dataIn2 = 32'd1; 
32'd9289: dataIn2 = 32'd0; 
32'd9290: dataIn2 = 32'd1; 
32'd9291: dataIn2 = 32'd0; 
32'd9292: dataIn2 = 32'd1; 
32'd9293: dataIn2 = 32'd0; 
32'd9294: dataIn2 = 32'd1; 
32'd9295: dataIn2 = 32'd0; 
32'd9296: dataIn2 = 32'd1; 
32'd9297: dataIn2 = 32'd0; 
32'd9298: dataIn2 = 32'd0; 
32'd9299: dataIn2 = 32'd1; 
32'd9300: dataIn2 = 32'd1; 
32'd9301: dataIn2 = 32'd0; 
32'd9302: dataIn2 = 32'd1; 
32'd9303: dataIn2 = 32'd1; 
32'd9304: dataIn2 = 32'd1; 
32'd9305: dataIn2 = 32'd1; 
32'd9306: dataIn2 = 32'd1; 
32'd9307: dataIn2 = 32'd0; 
32'd9308: dataIn2 = 32'd1; 
32'd9309: dataIn2 = 32'd1; 
32'd9310: dataIn2 = 32'd0; 
32'd9311: dataIn2 = 32'd0; 
32'd9312: dataIn2 = 32'd1; 
32'd9313: dataIn2 = 32'd1; 
32'd9314: dataIn2 = 32'd1; 
32'd9315: dataIn2 = 32'd0; 
32'd9316: dataIn2 = 32'd1; 
32'd9317: dataIn2 = 32'd0; 
32'd9318: dataIn2 = 32'd0; 
32'd9319: dataIn2 = 32'd0; 
32'd9320: dataIn2 = 32'd1; 
32'd9321: dataIn2 = 32'd1; 
32'd9322: dataIn2 = 32'd1; 
32'd9323: dataIn2 = 32'd1; 
32'd9324: dataIn2 = 32'd0; 
32'd9325: dataIn2 = 32'd1; 
32'd9326: dataIn2 = 32'd0; 
32'd9327: dataIn2 = 32'd0; 
32'd9328: dataIn2 = 32'd0; 
32'd9329: dataIn2 = 32'd1; 
32'd9330: dataIn2 = 32'd1; 
32'd9331: dataIn2 = 32'd1; 
32'd9332: dataIn2 = 32'd1; 
32'd9333: dataIn2 = 32'd1; 
32'd9334: dataIn2 = 32'd1; 
32'd9335: dataIn2 = 32'd1; 
32'd9336: dataIn2 = 32'd1; 
32'd9337: dataIn2 = 32'd1; 
32'd9338: dataIn2 = 32'd0; 
32'd9339: dataIn2 = 32'd0; 
32'd9340: dataIn2 = 32'd1; 
32'd9341: dataIn2 = 32'd1; 
32'd9342: dataIn2 = 32'd1; 
32'd9343: dataIn2 = 32'd1; 
32'd9344: dataIn2 = 32'd1; 
32'd9345: dataIn2 = 32'd0; 
32'd9346: dataIn2 = 32'd1; 
32'd9347: dataIn2 = 32'd1; 
32'd9348: dataIn2 = 32'd0; 
32'd9349: dataIn2 = 32'd0; 
32'd9350: dataIn2 = 32'd1; 
32'd9351: dataIn2 = 32'd1; 
32'd9352: dataIn2 = 32'd0; 
32'd9353: dataIn2 = 32'd1; 
32'd9354: dataIn2 = 32'd0; 
32'd9355: dataIn2 = 32'd1; 
32'd9356: dataIn2 = 32'd1; 
32'd9357: dataIn2 = 32'd0; 
32'd9358: dataIn2 = 32'd0; 
32'd9359: dataIn2 = 32'd0; 
32'd9360: dataIn2 = 32'd0; 
32'd9361: dataIn2 = 32'd1; 
32'd9362: dataIn2 = 32'd0; 
32'd9363: dataIn2 = 32'd1; 
32'd9364: dataIn2 = 32'd0; 
32'd9365: dataIn2 = 32'd1; 
32'd9366: dataIn2 = 32'd1; 
32'd9367: dataIn2 = 32'd0; 
32'd9368: dataIn2 = 32'd1; 
32'd9369: dataIn2 = 32'd1; 
32'd9370: dataIn2 = 32'd0; 
32'd9371: dataIn2 = 32'd0; 
32'd9372: dataIn2 = 32'd1; 
32'd9373: dataIn2 = 32'd1; 
32'd9374: dataIn2 = 32'd1; 
32'd9375: dataIn2 = 32'd0; 
32'd9376: dataIn2 = 32'd1; 
32'd9377: dataIn2 = 32'd0; 
32'd9378: dataIn2 = 32'd0; 
32'd9379: dataIn2 = 32'd1; 
32'd9380: dataIn2 = 32'd1; 
32'd9381: dataIn2 = 32'd0; 
32'd9382: dataIn2 = 32'd0; 
32'd9383: dataIn2 = 32'd1; 
32'd9384: dataIn2 = 32'd1; 
32'd9385: dataIn2 = 32'd0; 
32'd9386: dataIn2 = 32'd1; 
32'd9387: dataIn2 = 32'd1; 
32'd9388: dataIn2 = 32'd0; 
32'd9389: dataIn2 = 32'd1; 
32'd9390: dataIn2 = 32'd1; 
32'd9391: dataIn2 = 32'd1; 
32'd9392: dataIn2 = 32'd0; 
32'd9393: dataIn2 = 32'd1; 
32'd9394: dataIn2 = 32'd0; 
32'd9395: dataIn2 = 32'd0; 
32'd9396: dataIn2 = 32'd1; 
32'd9397: dataIn2 = 32'd1; 
32'd9398: dataIn2 = 32'd1; 
32'd9399: dataIn2 = 32'd0; 
32'd9400: dataIn2 = 32'd1; 
32'd9401: dataIn2 = 32'd0; 
32'd9402: dataIn2 = 32'd1; 
32'd9403: dataIn2 = 32'd1; 
32'd9404: dataIn2 = 32'd0; 
32'd9405: dataIn2 = 32'd0; 
32'd9406: dataIn2 = 32'd0; 
32'd9407: dataIn2 = 32'd1; 
32'd9408: dataIn2 = 32'd1; 
32'd9409: dataIn2 = 32'd0; 
32'd9410: dataIn2 = 32'd1; 
32'd9411: dataIn2 = 32'd0; 
32'd9412: dataIn2 = 32'd0; 
32'd9413: dataIn2 = 32'd0; 
32'd9414: dataIn2 = 32'd0; 
32'd9415: dataIn2 = 32'd0; 
32'd9416: dataIn2 = 32'd1; 
32'd9417: dataIn2 = 32'd1; 
32'd9418: dataIn2 = 32'd1; 
32'd9419: dataIn2 = 32'd0; 
32'd9420: dataIn2 = 32'd1; 
32'd9421: dataIn2 = 32'd0; 
32'd9422: dataIn2 = 32'd1; 
32'd9423: dataIn2 = 32'd0; 
32'd9424: dataIn2 = 32'd1; 
32'd9425: dataIn2 = 32'd0; 
32'd9426: dataIn2 = 32'd1; 
32'd9427: dataIn2 = 32'd1; 
32'd9428: dataIn2 = 32'd1; 
32'd9429: dataIn2 = 32'd0; 
32'd9430: dataIn2 = 32'd0; 
32'd9431: dataIn2 = 32'd1; 
32'd9432: dataIn2 = 32'd0; 
32'd9433: dataIn2 = 32'd0; 
32'd9434: dataIn2 = 32'd0; 
32'd9435: dataIn2 = 32'd1; 
32'd9436: dataIn2 = 32'd0; 
32'd9437: dataIn2 = 32'd0; 
32'd9438: dataIn2 = 32'd0; 
32'd9439: dataIn2 = 32'd0; 
32'd9440: dataIn2 = 32'd0; 
32'd9441: dataIn2 = 32'd1; 
32'd9442: dataIn2 = 32'd0; 
32'd9443: dataIn2 = 32'd0; 
32'd9444: dataIn2 = 32'd1; 
32'd9445: dataIn2 = 32'd0; 
32'd9446: dataIn2 = 32'd1; 
32'd9447: dataIn2 = 32'd1; 
32'd9448: dataIn2 = 32'd1; 
32'd9449: dataIn2 = 32'd1; 
32'd9450: dataIn2 = 32'd1; 
32'd9451: dataIn2 = 32'd1; 
32'd9452: dataIn2 = 32'd0; 
32'd9453: dataIn2 = 32'd0; 
32'd9454: dataIn2 = 32'd0; 
32'd9455: dataIn2 = 32'd1; 
32'd9456: dataIn2 = 32'd1; 
32'd9457: dataIn2 = 32'd0; 
32'd9458: dataIn2 = 32'd1; 
32'd9459: dataIn2 = 32'd0; 
32'd9460: dataIn2 = 32'd1; 
32'd9461: dataIn2 = 32'd0; 
32'd9462: dataIn2 = 32'd0; 
32'd9463: dataIn2 = 32'd1; 
32'd9464: dataIn2 = 32'd0; 
32'd9465: dataIn2 = 32'd1; 
32'd9466: dataIn2 = 32'd0; 
32'd9467: dataIn2 = 32'd1; 
32'd9468: dataIn2 = 32'd0; 
32'd9469: dataIn2 = 32'd1; 
32'd9470: dataIn2 = 32'd1; 
32'd9471: dataIn2 = 32'd1; 
32'd9472: dataIn2 = 32'd1; 
32'd9473: dataIn2 = 32'd0; 
32'd9474: dataIn2 = 32'd0; 
32'd9475: dataIn2 = 32'd0; 
32'd9476: dataIn2 = 32'd1; 
32'd9477: dataIn2 = 32'd0; 
32'd9478: dataIn2 = 32'd0; 
32'd9479: dataIn2 = 32'd0; 
32'd9480: dataIn2 = 32'd1; 
32'd9481: dataIn2 = 32'd1; 
32'd9482: dataIn2 = 32'd0; 
32'd9483: dataIn2 = 32'd0; 
32'd9484: dataIn2 = 32'd0; 
32'd9485: dataIn2 = 32'd1; 
32'd9486: dataIn2 = 32'd1; 
32'd9487: dataIn2 = 32'd0; 
32'd9488: dataIn2 = 32'd1; 
32'd9489: dataIn2 = 32'd0; 
32'd9490: dataIn2 = 32'd0; 
32'd9491: dataIn2 = 32'd1; 
32'd9492: dataIn2 = 32'd1; 
32'd9493: dataIn2 = 32'd0; 
32'd9494: dataIn2 = 32'd0; 
32'd9495: dataIn2 = 32'd0; 
32'd9496: dataIn2 = 32'd0; 
32'd9497: dataIn2 = 32'd0; 
32'd9498: dataIn2 = 32'd0; 
32'd9499: dataIn2 = 32'd1; 
32'd9500: dataIn2 = 32'd1; 
32'd9501: dataIn2 = 32'd1; 
32'd9502: dataIn2 = 32'd0; 
32'd9503: dataIn2 = 32'd0; 
32'd9504: dataIn2 = 32'd1; 
32'd9505: dataIn2 = 32'd0; 
32'd9506: dataIn2 = 32'd1; 
32'd9507: dataIn2 = 32'd1; 
32'd9508: dataIn2 = 32'd0; 
32'd9509: dataIn2 = 32'd1; 
32'd9510: dataIn2 = 32'd1; 
32'd9511: dataIn2 = 32'd0; 
32'd9512: dataIn2 = 32'd1; 
32'd9513: dataIn2 = 32'd0; 
32'd9514: dataIn2 = 32'd1; 
32'd9515: dataIn2 = 32'd0; 
32'd9516: dataIn2 = 32'd0; 
32'd9517: dataIn2 = 32'd0; 
32'd9518: dataIn2 = 32'd0; 
32'd9519: dataIn2 = 32'd0; 
32'd9520: dataIn2 = 32'd0; 
32'd9521: dataIn2 = 32'd0; 
32'd9522: dataIn2 = 32'd1; 
32'd9523: dataIn2 = 32'd0; 
32'd9524: dataIn2 = 32'd0; 
32'd9525: dataIn2 = 32'd1; 
32'd9526: dataIn2 = 32'd0; 
32'd9527: dataIn2 = 32'd0; 
32'd9528: dataIn2 = 32'd0; 
32'd9529: dataIn2 = 32'd0; 
32'd9530: dataIn2 = 32'd0; 
32'd9531: dataIn2 = 32'd0; 
32'd9532: dataIn2 = 32'd0; 
32'd9533: dataIn2 = 32'd0; 
32'd9534: dataIn2 = 32'd0; 
32'd9535: dataIn2 = 32'd1; 
32'd9536: dataIn2 = 32'd1; 
32'd9537: dataIn2 = 32'd0; 
32'd9538: dataIn2 = 32'd0; 
32'd9539: dataIn2 = 32'd0; 
32'd9540: dataIn2 = 32'd0; 
32'd9541: dataIn2 = 32'd0; 
32'd9542: dataIn2 = 32'd1; 
32'd9543: dataIn2 = 32'd1; 
32'd9544: dataIn2 = 32'd0; 
32'd9545: dataIn2 = 32'd0; 
32'd9546: dataIn2 = 32'd1; 
32'd9547: dataIn2 = 32'd0; 
32'd9548: dataIn2 = 32'd0; 
32'd9549: dataIn2 = 32'd0; 
32'd9550: dataIn2 = 32'd0; 
32'd9551: dataIn2 = 32'd0; 
32'd9552: dataIn2 = 32'd1; 
32'd9553: dataIn2 = 32'd1; 
32'd9554: dataIn2 = 32'd1; 
32'd9555: dataIn2 = 32'd1; 
32'd9556: dataIn2 = 32'd1; 
32'd9557: dataIn2 = 32'd1; 
32'd9558: dataIn2 = 32'd1; 
32'd9559: dataIn2 = 32'd1; 
32'd9560: dataIn2 = 32'd1; 
32'd9561: dataIn2 = 32'd0; 
32'd9562: dataIn2 = 32'd0; 
32'd9563: dataIn2 = 32'd1; 
32'd9564: dataIn2 = 32'd1; 
32'd9565: dataIn2 = 32'd0; 
32'd9566: dataIn2 = 32'd0; 
32'd9567: dataIn2 = 32'd1; 
32'd9568: dataIn2 = 32'd1; 
32'd9569: dataIn2 = 32'd1; 
32'd9570: dataIn2 = 32'd0; 
32'd9571: dataIn2 = 32'd1; 
32'd9572: dataIn2 = 32'd0; 
32'd9573: dataIn2 = 32'd1; 
32'd9574: dataIn2 = 32'd0; 
32'd9575: dataIn2 = 32'd0; 
32'd9576: dataIn2 = 32'd1; 
32'd9577: dataIn2 = 32'd0; 
32'd9578: dataIn2 = 32'd0; 
32'd9579: dataIn2 = 32'd1; 
32'd9580: dataIn2 = 32'd0; 
32'd9581: dataIn2 = 32'd1; 
32'd9582: dataIn2 = 32'd0; 
32'd9583: dataIn2 = 32'd0; 
32'd9584: dataIn2 = 32'd0; 
32'd9585: dataIn2 = 32'd0; 
32'd9586: dataIn2 = 32'd0; 
32'd9587: dataIn2 = 32'd0; 
32'd9588: dataIn2 = 32'd1; 
32'd9589: dataIn2 = 32'd0; 
32'd9590: dataIn2 = 32'd1; 
32'd9591: dataIn2 = 32'd1; 
32'd9592: dataIn2 = 32'd0; 
32'd9593: dataIn2 = 32'd1; 
32'd9594: dataIn2 = 32'd0; 
32'd9595: dataIn2 = 32'd0; 
32'd9596: dataIn2 = 32'd1; 
32'd9597: dataIn2 = 32'd1; 
32'd9598: dataIn2 = 32'd1; 
32'd9599: dataIn2 = 32'd0; 
32'd9600: dataIn2 = 32'd1; 
32'd9601: dataIn2 = 32'd0; 
32'd9602: dataIn2 = 32'd0; 
32'd9603: dataIn2 = 32'd0; 
32'd9604: dataIn2 = 32'd0; 
32'd9605: dataIn2 = 32'd1; 
32'd9606: dataIn2 = 32'd0; 
32'd9607: dataIn2 = 32'd1; 
32'd9608: dataIn2 = 32'd1; 
32'd9609: dataIn2 = 32'd0; 
32'd9610: dataIn2 = 32'd1; 
32'd9611: dataIn2 = 32'd0; 
32'd9612: dataIn2 = 32'd1; 
32'd9613: dataIn2 = 32'd0; 
32'd9614: dataIn2 = 32'd0; 
32'd9615: dataIn2 = 32'd1; 
32'd9616: dataIn2 = 32'd1; 
32'd9617: dataIn2 = 32'd0; 
32'd9618: dataIn2 = 32'd0; 
32'd9619: dataIn2 = 32'd0; 
32'd9620: dataIn2 = 32'd0; 
32'd9621: dataIn2 = 32'd0; 
32'd9622: dataIn2 = 32'd0; 
32'd9623: dataIn2 = 32'd0; 
32'd9624: dataIn2 = 32'd1; 
32'd9625: dataIn2 = 32'd0; 
32'd9626: dataIn2 = 32'd0; 
32'd9627: dataIn2 = 32'd0; 
32'd9628: dataIn2 = 32'd1; 
32'd9629: dataIn2 = 32'd1; 
32'd9630: dataIn2 = 32'd1; 
32'd9631: dataIn2 = 32'd1; 
32'd9632: dataIn2 = 32'd1; 
32'd9633: dataIn2 = 32'd1; 
32'd9634: dataIn2 = 32'd0; 
32'd9635: dataIn2 = 32'd1; 
32'd9636: dataIn2 = 32'd1; 
32'd9637: dataIn2 = 32'd1; 
32'd9638: dataIn2 = 32'd1; 
32'd9639: dataIn2 = 32'd0; 
32'd9640: dataIn2 = 32'd0; 
32'd9641: dataIn2 = 32'd1; 
32'd9642: dataIn2 = 32'd0; 
32'd9643: dataIn2 = 32'd1; 
32'd9644: dataIn2 = 32'd1; 
32'd9645: dataIn2 = 32'd1; 
32'd9646: dataIn2 = 32'd0; 
32'd9647: dataIn2 = 32'd0; 
32'd9648: dataIn2 = 32'd0; 
32'd9649: dataIn2 = 32'd0; 
32'd9650: dataIn2 = 32'd1; 
32'd9651: dataIn2 = 32'd0; 
32'd9652: dataIn2 = 32'd0; 
32'd9653: dataIn2 = 32'd1; 
32'd9654: dataIn2 = 32'd1; 
32'd9655: dataIn2 = 32'd0; 
32'd9656: dataIn2 = 32'd0; 
32'd9657: dataIn2 = 32'd0; 
32'd9658: dataIn2 = 32'd1; 
32'd9659: dataIn2 = 32'd1; 
32'd9660: dataIn2 = 32'd1; 
32'd9661: dataIn2 = 32'd1; 
32'd9662: dataIn2 = 32'd0; 
32'd9663: dataIn2 = 32'd0; 
32'd9664: dataIn2 = 32'd1; 
32'd9665: dataIn2 = 32'd1; 
32'd9666: dataIn2 = 32'd0; 
32'd9667: dataIn2 = 32'd0; 
32'd9668: dataIn2 = 32'd0; 
32'd9669: dataIn2 = 32'd1; 
32'd9670: dataIn2 = 32'd1; 
32'd9671: dataIn2 = 32'd1; 
32'd9672: dataIn2 = 32'd0; 
32'd9673: dataIn2 = 32'd0; 
32'd9674: dataIn2 = 32'd0; 
32'd9675: dataIn2 = 32'd0; 
32'd9676: dataIn2 = 32'd0; 
32'd9677: dataIn2 = 32'd1; 
32'd9678: dataIn2 = 32'd0; 
32'd9679: dataIn2 = 32'd0; 
32'd9680: dataIn2 = 32'd0; 
32'd9681: dataIn2 = 32'd0; 
32'd9682: dataIn2 = 32'd0; 
32'd9683: dataIn2 = 32'd1; 
32'd9684: dataIn2 = 32'd0; 
32'd9685: dataIn2 = 32'd1; 
32'd9686: dataIn2 = 32'd1; 
32'd9687: dataIn2 = 32'd1; 
32'd9688: dataIn2 = 32'd1; 
32'd9689: dataIn2 = 32'd1; 
32'd9690: dataIn2 = 32'd0; 
32'd9691: dataIn2 = 32'd0; 
32'd9692: dataIn2 = 32'd0; 
32'd9693: dataIn2 = 32'd0; 
32'd9694: dataIn2 = 32'd0; 
32'd9695: dataIn2 = 32'd0; 
32'd9696: dataIn2 = 32'd0; 
32'd9697: dataIn2 = 32'd0; 
32'd9698: dataIn2 = 32'd1; 
32'd9699: dataIn2 = 32'd0; 
32'd9700: dataIn2 = 32'd1; 
32'd9701: dataIn2 = 32'd1; 
32'd9702: dataIn2 = 32'd0; 
32'd9703: dataIn2 = 32'd1; 
32'd9704: dataIn2 = 32'd0; 
32'd9705: dataIn2 = 32'd1; 
32'd9706: dataIn2 = 32'd1; 
32'd9707: dataIn2 = 32'd0; 
32'd9708: dataIn2 = 32'd0; 
32'd9709: dataIn2 = 32'd1; 
32'd9710: dataIn2 = 32'd1; 
32'd9711: dataIn2 = 32'd0; 
32'd9712: dataIn2 = 32'd1; 
32'd9713: dataIn2 = 32'd1; 
32'd9714: dataIn2 = 32'd1; 
32'd9715: dataIn2 = 32'd0; 
32'd9716: dataIn2 = 32'd0; 
32'd9717: dataIn2 = 32'd0; 
32'd9718: dataIn2 = 32'd0; 
32'd9719: dataIn2 = 32'd1; 
32'd9720: dataIn2 = 32'd0; 
32'd9721: dataIn2 = 32'd1; 
32'd9722: dataIn2 = 32'd0; 
32'd9723: dataIn2 = 32'd0; 
32'd9724: dataIn2 = 32'd0; 
32'd9725: dataIn2 = 32'd1; 
32'd9726: dataIn2 = 32'd1; 
32'd9727: dataIn2 = 32'd0; 
32'd9728: dataIn2 = 32'd0; 
32'd9729: dataIn2 = 32'd0; 
32'd9730: dataIn2 = 32'd0; 
32'd9731: dataIn2 = 32'd0; 
32'd9732: dataIn2 = 32'd1; 
32'd9733: dataIn2 = 32'd0; 
32'd9734: dataIn2 = 32'd0; 
32'd9735: dataIn2 = 32'd0; 
32'd9736: dataIn2 = 32'd1; 
32'd9737: dataIn2 = 32'd0; 
32'd9738: dataIn2 = 32'd1; 
32'd9739: dataIn2 = 32'd0; 
32'd9740: dataIn2 = 32'd1; 
32'd9741: dataIn2 = 32'd0; 
32'd9742: dataIn2 = 32'd1; 
32'd9743: dataIn2 = 32'd0; 
32'd9744: dataIn2 = 32'd0; 
32'd9745: dataIn2 = 32'd1; 
32'd9746: dataIn2 = 32'd0; 
32'd9747: dataIn2 = 32'd0; 
32'd9748: dataIn2 = 32'd1; 
32'd9749: dataIn2 = 32'd0; 
32'd9750: dataIn2 = 32'd0; 
32'd9751: dataIn2 = 32'd1; 
32'd9752: dataIn2 = 32'd0; 
32'd9753: dataIn2 = 32'd0; 
32'd9754: dataIn2 = 32'd1; 
32'd9755: dataIn2 = 32'd0; 
32'd9756: dataIn2 = 32'd0; 
32'd9757: dataIn2 = 32'd0; 
32'd9758: dataIn2 = 32'd0; 
32'd9759: dataIn2 = 32'd1; 
32'd9760: dataIn2 = 32'd0; 
32'd9761: dataIn2 = 32'd1; 
32'd9762: dataIn2 = 32'd1; 
32'd9763: dataIn2 = 32'd1; 
32'd9764: dataIn2 = 32'd1; 
32'd9765: dataIn2 = 32'd1; 
32'd9766: dataIn2 = 32'd1; 
32'd9767: dataIn2 = 32'd0; 
32'd9768: dataIn2 = 32'd0; 
32'd9769: dataIn2 = 32'd0; 
32'd9770: dataIn2 = 32'd1; 
32'd9771: dataIn2 = 32'd1; 
32'd9772: dataIn2 = 32'd0; 
32'd9773: dataIn2 = 32'd0; 
32'd9774: dataIn2 = 32'd1; 
32'd9775: dataIn2 = 32'd0; 
32'd9776: dataIn2 = 32'd0; 
32'd9777: dataIn2 = 32'd1; 
32'd9778: dataIn2 = 32'd0; 
32'd9779: dataIn2 = 32'd1; 
32'd9780: dataIn2 = 32'd0; 
32'd9781: dataIn2 = 32'd0; 
32'd9782: dataIn2 = 32'd1; 
32'd9783: dataIn2 = 32'd0; 
32'd9784: dataIn2 = 32'd0; 
32'd9785: dataIn2 = 32'd1; 
32'd9786: dataIn2 = 32'd1; 
32'd9787: dataIn2 = 32'd0; 
32'd9788: dataIn2 = 32'd0; 
32'd9789: dataIn2 = 32'd0; 
32'd9790: dataIn2 = 32'd0; 
32'd9791: dataIn2 = 32'd1; 
32'd9792: dataIn2 = 32'd0; 
32'd9793: dataIn2 = 32'd1; 
32'd9794: dataIn2 = 32'd1; 
32'd9795: dataIn2 = 32'd1; 
32'd9796: dataIn2 = 32'd0; 
32'd9797: dataIn2 = 32'd1; 
32'd9798: dataIn2 = 32'd0; 
32'd9799: dataIn2 = 32'd1; 
32'd9800: dataIn2 = 32'd0; 
32'd9801: dataIn2 = 32'd1; 
32'd9802: dataIn2 = 32'd1; 
32'd9803: dataIn2 = 32'd1; 
32'd9804: dataIn2 = 32'd1; 
32'd9805: dataIn2 = 32'd0; 
32'd9806: dataIn2 = 32'd1; 
32'd9807: dataIn2 = 32'd1; 
32'd9808: dataIn2 = 32'd1; 
32'd9809: dataIn2 = 32'd1; 
32'd9810: dataIn2 = 32'd1; 
32'd9811: dataIn2 = 32'd0; 
32'd9812: dataIn2 = 32'd0; 
32'd9813: dataIn2 = 32'd0; 
32'd9814: dataIn2 = 32'd0; 
32'd9815: dataIn2 = 32'd0; 
32'd9816: dataIn2 = 32'd1; 
32'd9817: dataIn2 = 32'd0; 
32'd9818: dataIn2 = 32'd1; 
32'd9819: dataIn2 = 32'd1; 
32'd9820: dataIn2 = 32'd0; 
32'd9821: dataIn2 = 32'd0; 
32'd9822: dataIn2 = 32'd1; 
32'd9823: dataIn2 = 32'd1; 
32'd9824: dataIn2 = 32'd1; 
32'd9825: dataIn2 = 32'd0; 
32'd9826: dataIn2 = 32'd0; 
32'd9827: dataIn2 = 32'd1; 
32'd9828: dataIn2 = 32'd1; 
32'd9829: dataIn2 = 32'd0; 
32'd9830: dataIn2 = 32'd0; 
32'd9831: dataIn2 = 32'd1; 
32'd9832: dataIn2 = 32'd0; 
32'd9833: dataIn2 = 32'd1; 
32'd9834: dataIn2 = 32'd1; 
32'd9835: dataIn2 = 32'd1; 
32'd9836: dataIn2 = 32'd0; 
32'd9837: dataIn2 = 32'd0; 
32'd9838: dataIn2 = 32'd0; 
32'd9839: dataIn2 = 32'd0; 
32'd9840: dataIn2 = 32'd1; 
32'd9841: dataIn2 = 32'd0; 
32'd9842: dataIn2 = 32'd0; 
32'd9843: dataIn2 = 32'd0; 
32'd9844: dataIn2 = 32'd0; 
32'd9845: dataIn2 = 32'd0; 
32'd9846: dataIn2 = 32'd1; 
32'd9847: dataIn2 = 32'd1; 
32'd9848: dataIn2 = 32'd0; 
32'd9849: dataIn2 = 32'd1; 
32'd9850: dataIn2 = 32'd0; 
32'd9851: dataIn2 = 32'd1; 
32'd9852: dataIn2 = 32'd1; 
32'd9853: dataIn2 = 32'd1; 
32'd9854: dataIn2 = 32'd1; 
32'd9855: dataIn2 = 32'd0; 
32'd9856: dataIn2 = 32'd1; 
32'd9857: dataIn2 = 32'd0; 
32'd9858: dataIn2 = 32'd1; 
32'd9859: dataIn2 = 32'd1; 
32'd9860: dataIn2 = 32'd0; 
32'd9861: dataIn2 = 32'd1; 
32'd9862: dataIn2 = 32'd0; 
32'd9863: dataIn2 = 32'd0; 
32'd9864: dataIn2 = 32'd1; 
32'd9865: dataIn2 = 32'd0; 
32'd9866: dataIn2 = 32'd0; 
32'd9867: dataIn2 = 32'd0; 
32'd9868: dataIn2 = 32'd1; 
32'd9869: dataIn2 = 32'd0; 
32'd9870: dataIn2 = 32'd1; 
32'd9871: dataIn2 = 32'd1; 
32'd9872: dataIn2 = 32'd0; 
32'd9873: dataIn2 = 32'd0; 
32'd9874: dataIn2 = 32'd1; 
32'd9875: dataIn2 = 32'd0; 
32'd9876: dataIn2 = 32'd1; 
32'd9877: dataIn2 = 32'd1; 
32'd9878: dataIn2 = 32'd0; 
32'd9879: dataIn2 = 32'd1; 
32'd9880: dataIn2 = 32'd1; 
32'd9881: dataIn2 = 32'd1; 
32'd9882: dataIn2 = 32'd1; 
32'd9883: dataIn2 = 32'd0; 
32'd9884: dataIn2 = 32'd1; 
32'd9885: dataIn2 = 32'd0; 
32'd9886: dataIn2 = 32'd1; 
32'd9887: dataIn2 = 32'd0; 
32'd9888: dataIn2 = 32'd0; 
32'd9889: dataIn2 = 32'd1; 
32'd9890: dataIn2 = 32'd1; 
32'd9891: dataIn2 = 32'd0; 
32'd9892: dataIn2 = 32'd0; 
32'd9893: dataIn2 = 32'd0; 
32'd9894: dataIn2 = 32'd0; 
32'd9895: dataIn2 = 32'd1; 
32'd9896: dataIn2 = 32'd0; 
32'd9897: dataIn2 = 32'd0; 
32'd9898: dataIn2 = 32'd0; 
32'd9899: dataIn2 = 32'd1; 
32'd9900: dataIn2 = 32'd0; 
32'd9901: dataIn2 = 32'd0; 
32'd9902: dataIn2 = 32'd1; 
32'd9903: dataIn2 = 32'd0; 
32'd9904: dataIn2 = 32'd0; 
32'd9905: dataIn2 = 32'd1; 
32'd9906: dataIn2 = 32'd0; 
32'd9907: dataIn2 = 32'd0; 
32'd9908: dataIn2 = 32'd1; 
32'd9909: dataIn2 = 32'd1; 
32'd9910: dataIn2 = 32'd1; 
32'd9911: dataIn2 = 32'd0; 
32'd9912: dataIn2 = 32'd0; 
32'd9913: dataIn2 = 32'd1; 
32'd9914: dataIn2 = 32'd0; 
32'd9915: dataIn2 = 32'd0; 
32'd9916: dataIn2 = 32'd0; 
32'd9917: dataIn2 = 32'd0; 
32'd9918: dataIn2 = 32'd0; 
32'd9919: dataIn2 = 32'd1; 
32'd9920: dataIn2 = 32'd0; 
32'd9921: dataIn2 = 32'd0; 
32'd9922: dataIn2 = 32'd1; 
32'd9923: dataIn2 = 32'd1; 
32'd9924: dataIn2 = 32'd1; 
32'd9925: dataIn2 = 32'd0; 
32'd9926: dataIn2 = 32'd1; 
32'd9927: dataIn2 = 32'd0; 
32'd9928: dataIn2 = 32'd0; 
32'd9929: dataIn2 = 32'd1; 
32'd9930: dataIn2 = 32'd0; 
32'd9931: dataIn2 = 32'd0; 
32'd9932: dataIn2 = 32'd1; 
32'd9933: dataIn2 = 32'd0; 
32'd9934: dataIn2 = 32'd0; 
32'd9935: dataIn2 = 32'd1; 
32'd9936: dataIn2 = 32'd1; 
32'd9937: dataIn2 = 32'd1; 
32'd9938: dataIn2 = 32'd0; 
32'd9939: dataIn2 = 32'd0; 
32'd9940: dataIn2 = 32'd1; 
32'd9941: dataIn2 = 32'd1; 
32'd9942: dataIn2 = 32'd1; 
32'd9943: dataIn2 = 32'd1; 
32'd9944: dataIn2 = 32'd0; 
32'd9945: dataIn2 = 32'd1; 
32'd9946: dataIn2 = 32'd1; 
32'd9947: dataIn2 = 32'd0; 
32'd9948: dataIn2 = 32'd0; 
32'd9949: dataIn2 = 32'd1; 
32'd9950: dataIn2 = 32'd0; 
32'd9951: dataIn2 = 32'd1; 
32'd9952: dataIn2 = 32'd0; 
32'd9953: dataIn2 = 32'd0; 
32'd9954: dataIn2 = 32'd0; 
32'd9955: dataIn2 = 32'd1; 
32'd9956: dataIn2 = 32'd0; 
32'd9957: dataIn2 = 32'd1; 
32'd9958: dataIn2 = 32'd1; 
32'd9959: dataIn2 = 32'd1; 
32'd9960: dataIn2 = 32'd0; 
32'd9961: dataIn2 = 32'd1; 
32'd9962: dataIn2 = 32'd0; 
32'd9963: dataIn2 = 32'd0; 
32'd9964: dataIn2 = 32'd1; 
32'd9965: dataIn2 = 32'd0; 
32'd9966: dataIn2 = 32'd1; 
32'd9967: dataIn2 = 32'd1; 
32'd9968: dataIn2 = 32'd1; 
32'd9969: dataIn2 = 32'd1; 
32'd9970: dataIn2 = 32'd0; 
32'd9971: dataIn2 = 32'd1; 
32'd9972: dataIn2 = 32'd1; 
32'd9973: dataIn2 = 32'd0; 
32'd9974: dataIn2 = 32'd1; 
32'd9975: dataIn2 = 32'd1; 
32'd9976: dataIn2 = 32'd0; 
32'd9977: dataIn2 = 32'd0; 
32'd9978: dataIn2 = 32'd0; 
32'd9979: dataIn2 = 32'd1; 
32'd9980: dataIn2 = 32'd1; 
32'd9981: dataIn2 = 32'd1; 
32'd9982: dataIn2 = 32'd1; 
32'd9983: dataIn2 = 32'd1; 
32'd9984: dataIn2 = 32'd1; 
32'd9985: dataIn2 = 32'd0; 
32'd9986: dataIn2 = 32'd1; 
32'd9987: dataIn2 = 32'd1; 
32'd9988: dataIn2 = 32'd1; 
32'd9989: dataIn2 = 32'd1; 
32'd9990: dataIn2 = 32'd0; 
32'd9991: dataIn2 = 32'd0; 
32'd9992: dataIn2 = 32'd0; 
32'd9993: dataIn2 = 32'd0; 
32'd9994: dataIn2 = 32'd0; 
32'd9995: dataIn2 = 32'd1; 
32'd9996: dataIn2 = 32'd0; 
32'd9997: dataIn2 = 32'd1; 
32'd9998: dataIn2 = 32'd1; 
32'd9999: dataIn2 = 32'd1; 
32'd10000: dataIn2 = 32'd1; 
32'd10001: dataIn2 = 32'd1; 
32'd10002: dataIn2 = 32'd1; 
32'd10003: dataIn2 = 32'd0; 
32'd10004: dataIn2 = 32'd1; 
32'd10005: dataIn2 = 32'd0; 
32'd10006: dataIn2 = 32'd1; 
32'd10007: dataIn2 = 32'd0; 
32'd10008: dataIn2 = 32'd0; 
32'd10009: dataIn2 = 32'd1; 
32'd10010: dataIn2 = 32'd1; 
32'd10011: dataIn2 = 32'd1; 
32'd10012: dataIn2 = 32'd0; 
32'd10013: dataIn2 = 32'd0; 
32'd10014: dataIn2 = 32'd0; 
32'd10015: dataIn2 = 32'd0; 
32'd10016: dataIn2 = 32'd1; 
32'd10017: dataIn2 = 32'd0; 
32'd10018: dataIn2 = 32'd1; 
32'd10019: dataIn2 = 32'd1; 
32'd10020: dataIn2 = 32'd1; 
32'd10021: dataIn2 = 32'd1; 
32'd10022: dataIn2 = 32'd0; 
32'd10023: dataIn2 = 32'd0; 
32'd10024: dataIn2 = 32'd0; 
32'd10025: dataIn2 = 32'd0; 
32'd10026: dataIn2 = 32'd1; 
32'd10027: dataIn2 = 32'd1; 
32'd10028: dataIn2 = 32'd1; 
32'd10029: dataIn2 = 32'd0; 
32'd10030: dataIn2 = 32'd0; 
32'd10031: dataIn2 = 32'd1; 
32'd10032: dataIn2 = 32'd1; 
32'd10033: dataIn2 = 32'd1; 
32'd10034: dataIn2 = 32'd0; 
32'd10035: dataIn2 = 32'd0; 
32'd10036: dataIn2 = 32'd0; 
32'd10037: dataIn2 = 32'd1; 
32'd10038: dataIn2 = 32'd0; 
32'd10039: dataIn2 = 32'd1; 
32'd10040: dataIn2 = 32'd1; 
32'd10041: dataIn2 = 32'd1; 
32'd10042: dataIn2 = 32'd0; 
32'd10043: dataIn2 = 32'd1; 
32'd10044: dataIn2 = 32'd0; 
32'd10045: dataIn2 = 32'd0; 
32'd10046: dataIn2 = 32'd1; 
32'd10047: dataIn2 = 32'd1; 
32'd10048: dataIn2 = 32'd0; 
32'd10049: dataIn2 = 32'd1; 
32'd10050: dataIn2 = 32'd0; 
32'd10051: dataIn2 = 32'd0; 
32'd10052: dataIn2 = 32'd0; 
32'd10053: dataIn2 = 32'd0; 
32'd10054: dataIn2 = 32'd1; 
32'd10055: dataIn2 = 32'd1; 
32'd10056: dataIn2 = 32'd0; 
32'd10057: dataIn2 = 32'd0; 
32'd10058: dataIn2 = 32'd0; 
32'd10059: dataIn2 = 32'd1; 
32'd10060: dataIn2 = 32'd1; 
32'd10061: dataIn2 = 32'd0; 
32'd10062: dataIn2 = 32'd1; 
32'd10063: dataIn2 = 32'd1; 
32'd10064: dataIn2 = 32'd0; 
32'd10065: dataIn2 = 32'd1; 
32'd10066: dataIn2 = 32'd0; 
32'd10067: dataIn2 = 32'd1; 
32'd10068: dataIn2 = 32'd0; 
32'd10069: dataIn2 = 32'd1; 
32'd10070: dataIn2 = 32'd0; 
32'd10071: dataIn2 = 32'd1; 
32'd10072: dataIn2 = 32'd0; 
32'd10073: dataIn2 = 32'd1; 
32'd10074: dataIn2 = 32'd0; 
32'd10075: dataIn2 = 32'd1; 
32'd10076: dataIn2 = 32'd1; 
32'd10077: dataIn2 = 32'd1; 
32'd10078: dataIn2 = 32'd0; 
32'd10079: dataIn2 = 32'd0; 
32'd10080: dataIn2 = 32'd0; 
32'd10081: dataIn2 = 32'd1; 
32'd10082: dataIn2 = 32'd0; 
32'd10083: dataIn2 = 32'd0; 
32'd10084: dataIn2 = 32'd0; 
32'd10085: dataIn2 = 32'd0; 
32'd10086: dataIn2 = 32'd1; 
32'd10087: dataIn2 = 32'd1; 
32'd10088: dataIn2 = 32'd1; 
32'd10089: dataIn2 = 32'd1; 
32'd10090: dataIn2 = 32'd0; 
32'd10091: dataIn2 = 32'd0; 
32'd10092: dataIn2 = 32'd0; 
32'd10093: dataIn2 = 32'd1; 
32'd10094: dataIn2 = 32'd0; 
32'd10095: dataIn2 = 32'd0; 
32'd10096: dataIn2 = 32'd0; 
32'd10097: dataIn2 = 32'd1; 
32'd10098: dataIn2 = 32'd1; 
32'd10099: dataIn2 = 32'd1; 
32'd10100: dataIn2 = 32'd1; 
32'd10101: dataIn2 = 32'd1; 
32'd10102: dataIn2 = 32'd0; 
32'd10103: dataIn2 = 32'd0; 
32'd10104: dataIn2 = 32'd0; 
32'd10105: dataIn2 = 32'd1; 
32'd10106: dataIn2 = 32'd1; 
32'd10107: dataIn2 = 32'd0; 
32'd10108: dataIn2 = 32'd0; 
32'd10109: dataIn2 = 32'd1; 
32'd10110: dataIn2 = 32'd0; 
32'd10111: dataIn2 = 32'd1; 
32'd10112: dataIn2 = 32'd1; 
32'd10113: dataIn2 = 32'd1; 
32'd10114: dataIn2 = 32'd1; 
32'd10115: dataIn2 = 32'd1; 
32'd10116: dataIn2 = 32'd1; 
32'd10117: dataIn2 = 32'd0; 
32'd10118: dataIn2 = 32'd1; 
32'd10119: dataIn2 = 32'd0; 
32'd10120: dataIn2 = 32'd1; 
32'd10121: dataIn2 = 32'd0; 
32'd10122: dataIn2 = 32'd1; 
32'd10123: dataIn2 = 32'd0; 
32'd10124: dataIn2 = 32'd0; 
32'd10125: dataIn2 = 32'd0; 
32'd10126: dataIn2 = 32'd1; 
32'd10127: dataIn2 = 32'd1; 
32'd10128: dataIn2 = 32'd1; 
32'd10129: dataIn2 = 32'd0; 
32'd10130: dataIn2 = 32'd1; 
32'd10131: dataIn2 = 32'd0; 
32'd10132: dataIn2 = 32'd0; 
32'd10133: dataIn2 = 32'd1; 
32'd10134: dataIn2 = 32'd0; 
32'd10135: dataIn2 = 32'd0; 
32'd10136: dataIn2 = 32'd0; 
32'd10137: dataIn2 = 32'd1; 
32'd10138: dataIn2 = 32'd1; 
32'd10139: dataIn2 = 32'd1; 
32'd10140: dataIn2 = 32'd1; 
32'd10141: dataIn2 = 32'd0; 
32'd10142: dataIn2 = 32'd0; 
32'd10143: dataIn2 = 32'd0; 
32'd10144: dataIn2 = 32'd0; 
32'd10145: dataIn2 = 32'd0; 
32'd10146: dataIn2 = 32'd1; 
32'd10147: dataIn2 = 32'd0; 
32'd10148: dataIn2 = 32'd1; 
32'd10149: dataIn2 = 32'd1; 
32'd10150: dataIn2 = 32'd0; 
32'd10151: dataIn2 = 32'd0; 
32'd10152: dataIn2 = 32'd0; 
32'd10153: dataIn2 = 32'd1; 
32'd10154: dataIn2 = 32'd1; 
32'd10155: dataIn2 = 32'd0; 
32'd10156: dataIn2 = 32'd0; 
32'd10157: dataIn2 = 32'd1; 
32'd10158: dataIn2 = 32'd1; 
32'd10159: dataIn2 = 32'd0; 
32'd10160: dataIn2 = 32'd0; 
32'd10161: dataIn2 = 32'd1; 
32'd10162: dataIn2 = 32'd0; 
32'd10163: dataIn2 = 32'd0; 
32'd10164: dataIn2 = 32'd1; 
32'd10165: dataIn2 = 32'd1; 
32'd10166: dataIn2 = 32'd1; 
32'd10167: dataIn2 = 32'd1; 
32'd10168: dataIn2 = 32'd0; 
32'd10169: dataIn2 = 32'd0; 
32'd10170: dataIn2 = 32'd1; 
32'd10171: dataIn2 = 32'd0; 
32'd10172: dataIn2 = 32'd0; 
32'd10173: dataIn2 = 32'd0; 
32'd10174: dataIn2 = 32'd1; 
32'd10175: dataIn2 = 32'd0; 
32'd10176: dataIn2 = 32'd0; 
32'd10177: dataIn2 = 32'd1; 
32'd10178: dataIn2 = 32'd1; 
32'd10179: dataIn2 = 32'd1; 
32'd10180: dataIn2 = 32'd1; 
32'd10181: dataIn2 = 32'd0; 
32'd10182: dataIn2 = 32'd1; 
32'd10183: dataIn2 = 32'd0; 
32'd10184: dataIn2 = 32'd1; 
32'd10185: dataIn2 = 32'd1; 
32'd10186: dataIn2 = 32'd1; 
32'd10187: dataIn2 = 32'd0; 
32'd10188: dataIn2 = 32'd1; 
32'd10189: dataIn2 = 32'd0; 
32'd10190: dataIn2 = 32'd1; 
32'd10191: dataIn2 = 32'd1; 
32'd10192: dataIn2 = 32'd0; 
32'd10193: dataIn2 = 32'd1; 
32'd10194: dataIn2 = 32'd0; 
32'd10195: dataIn2 = 32'd0; 
32'd10196: dataIn2 = 32'd1; 
32'd10197: dataIn2 = 32'd1; 
32'd10198: dataIn2 = 32'd0; 
32'd10199: dataIn2 = 32'd0; 
32'd10200: dataIn2 = 32'd0; 
32'd10201: dataIn2 = 32'd0; 
32'd10202: dataIn2 = 32'd0; 
32'd10203: dataIn2 = 32'd0; 
32'd10204: dataIn2 = 32'd0; 
32'd10205: dataIn2 = 32'd1; 
32'd10206: dataIn2 = 32'd1; 
32'd10207: dataIn2 = 32'd0; 
32'd10208: dataIn2 = 32'd0; 
32'd10209: dataIn2 = 32'd1; 
32'd10210: dataIn2 = 32'd1; 
32'd10211: dataIn2 = 32'd0; 
32'd10212: dataIn2 = 32'd0; 
32'd10213: dataIn2 = 32'd0; 
32'd10214: dataIn2 = 32'd0; 
32'd10215: dataIn2 = 32'd0; 
32'd10216: dataIn2 = 32'd0; 
32'd10217: dataIn2 = 32'd1; 
32'd10218: dataIn2 = 32'd1; 
32'd10219: dataIn2 = 32'd1; 
32'd10220: dataIn2 = 32'd1; 
32'd10221: dataIn2 = 32'd1; 
32'd10222: dataIn2 = 32'd0; 
32'd10223: dataIn2 = 32'd0; 
32'd10224: dataIn2 = 32'd1; 
32'd10225: dataIn2 = 32'd1; 
32'd10226: dataIn2 = 32'd1; 
32'd10227: dataIn2 = 32'd1; 
32'd10228: dataIn2 = 32'd1; 
32'd10229: dataIn2 = 32'd0; 
32'd10230: dataIn2 = 32'd1; 
32'd10231: dataIn2 = 32'd1; 
32'd10232: dataIn2 = 32'd0; 
32'd10233: dataIn2 = 32'd1; 
32'd10234: dataIn2 = 32'd0; 
32'd10235: dataIn2 = 32'd1; 
32'd10236: dataIn2 = 32'd0; 
32'd10237: dataIn2 = 32'd0; 
32'd10238: dataIn2 = 32'd1; 
32'd10239: dataIn2 = 32'd1; 
32'd10240: dataIn2 = 32'd1; 
32'd10241: dataIn2 = 32'd1; 
32'd10242: dataIn2 = 32'd0; 
32'd10243: dataIn2 = 32'd1; 
32'd10244: dataIn2 = 32'd0; 
32'd10245: dataIn2 = 32'd1; 
32'd10246: dataIn2 = 32'd1; 
32'd10247: dataIn2 = 32'd0; 
32'd10248: dataIn2 = 32'd1; 
32'd10249: dataIn2 = 32'd1; 
32'd10250: dataIn2 = 32'd1; 
32'd10251: dataIn2 = 32'd1; 
32'd10252: dataIn2 = 32'd0; 
32'd10253: dataIn2 = 32'd1; 
32'd10254: dataIn2 = 32'd0; 
32'd10255: dataIn2 = 32'd0; 
32'd10256: dataIn2 = 32'd1; 
32'd10257: dataIn2 = 32'd1; 
32'd10258: dataIn2 = 32'd0; 
32'd10259: dataIn2 = 32'd1; 
32'd10260: dataIn2 = 32'd1; 
32'd10261: dataIn2 = 32'd1; 
32'd10262: dataIn2 = 32'd1; 
32'd10263: dataIn2 = 32'd1; 
32'd10264: dataIn2 = 32'd0; 
32'd10265: dataIn2 = 32'd1; 
32'd10266: dataIn2 = 32'd0; 
32'd10267: dataIn2 = 32'd1; 
32'd10268: dataIn2 = 32'd1; 
32'd10269: dataIn2 = 32'd1; 
32'd10270: dataIn2 = 32'd1; 
32'd10271: dataIn2 = 32'd0; 
32'd10272: dataIn2 = 32'd0; 
32'd10273: dataIn2 = 32'd0; 
32'd10274: dataIn2 = 32'd0; 
32'd10275: dataIn2 = 32'd0; 
32'd10276: dataIn2 = 32'd1; 
32'd10277: dataIn2 = 32'd0; 
32'd10278: dataIn2 = 32'd0; 
32'd10279: dataIn2 = 32'd0; 
32'd10280: dataIn2 = 32'd0; 
32'd10281: dataIn2 = 32'd0; 
32'd10282: dataIn2 = 32'd0; 
32'd10283: dataIn2 = 32'd0; 
32'd10284: dataIn2 = 32'd1; 
32'd10285: dataIn2 = 32'd0; 
32'd10286: dataIn2 = 32'd1; 
32'd10287: dataIn2 = 32'd1; 
32'd10288: dataIn2 = 32'd0; 
32'd10289: dataIn2 = 32'd1; 
32'd10290: dataIn2 = 32'd0; 
32'd10291: dataIn2 = 32'd0; 
32'd10292: dataIn2 = 32'd1; 
32'd10293: dataIn2 = 32'd0; 
32'd10294: dataIn2 = 32'd0; 
32'd10295: dataIn2 = 32'd0; 
32'd10296: dataIn2 = 32'd0; 
32'd10297: dataIn2 = 32'd0; 
32'd10298: dataIn2 = 32'd0; 
32'd10299: dataIn2 = 32'd1; 
32'd10300: dataIn2 = 32'd1; 
32'd10301: dataIn2 = 32'd1; 
32'd10302: dataIn2 = 32'd0; 
32'd10303: dataIn2 = 32'd1; 
32'd10304: dataIn2 = 32'd0; 
32'd10305: dataIn2 = 32'd1; 
32'd10306: dataIn2 = 32'd0; 
32'd10307: dataIn2 = 32'd0; 
32'd10308: dataIn2 = 32'd0; 
32'd10309: dataIn2 = 32'd0; 
32'd10310: dataIn2 = 32'd1; 
32'd10311: dataIn2 = 32'd0; 
32'd10312: dataIn2 = 32'd0; 
32'd10313: dataIn2 = 32'd0; 
32'd10314: dataIn2 = 32'd0; 
32'd10315: dataIn2 = 32'd0; 
32'd10316: dataIn2 = 32'd1; 
32'd10317: dataIn2 = 32'd0; 
32'd10318: dataIn2 = 32'd0; 
32'd10319: dataIn2 = 32'd0; 
32'd10320: dataIn2 = 32'd0; 
32'd10321: dataIn2 = 32'd0; 
32'd10322: dataIn2 = 32'd1; 
32'd10323: dataIn2 = 32'd0; 
32'd10324: dataIn2 = 32'd1; 
32'd10325: dataIn2 = 32'd1; 
32'd10326: dataIn2 = 32'd0; 
32'd10327: dataIn2 = 32'd0; 
32'd10328: dataIn2 = 32'd0; 
32'd10329: dataIn2 = 32'd0; 
32'd10330: dataIn2 = 32'd0; 
32'd10331: dataIn2 = 32'd1; 
32'd10332: dataIn2 = 32'd0; 
32'd10333: dataIn2 = 32'd1; 
32'd10334: dataIn2 = 32'd0; 
32'd10335: dataIn2 = 32'd1; 
32'd10336: dataIn2 = 32'd1; 
32'd10337: dataIn2 = 32'd1; 
32'd10338: dataIn2 = 32'd1; 
32'd10339: dataIn2 = 32'd1; 
32'd10340: dataIn2 = 32'd0; 
32'd10341: dataIn2 = 32'd0; 
32'd10342: dataIn2 = 32'd1; 
32'd10343: dataIn2 = 32'd0; 
32'd10344: dataIn2 = 32'd0; 
32'd10345: dataIn2 = 32'd0; 
32'd10346: dataIn2 = 32'd0; 
32'd10347: dataIn2 = 32'd0; 
32'd10348: dataIn2 = 32'd0; 
32'd10349: dataIn2 = 32'd1; 
32'd10350: dataIn2 = 32'd0; 
32'd10351: dataIn2 = 32'd1; 
32'd10352: dataIn2 = 32'd0; 
32'd10353: dataIn2 = 32'd1; 
32'd10354: dataIn2 = 32'd0; 
32'd10355: dataIn2 = 32'd0; 
32'd10356: dataIn2 = 32'd0; 
32'd10357: dataIn2 = 32'd1; 
32'd10358: dataIn2 = 32'd1; 
32'd10359: dataIn2 = 32'd1; 
32'd10360: dataIn2 = 32'd0; 
32'd10361: dataIn2 = 32'd0; 
32'd10362: dataIn2 = 32'd1; 
32'd10363: dataIn2 = 32'd1; 
32'd10364: dataIn2 = 32'd0; 
32'd10365: dataIn2 = 32'd0; 
32'd10366: dataIn2 = 32'd1; 
32'd10367: dataIn2 = 32'd0; 
32'd10368: dataIn2 = 32'd1; 
32'd10369: dataIn2 = 32'd1; 
32'd10370: dataIn2 = 32'd0; 
32'd10371: dataIn2 = 32'd0; 
32'd10372: dataIn2 = 32'd0; 
32'd10373: dataIn2 = 32'd1; 
32'd10374: dataIn2 = 32'd1; 
32'd10375: dataIn2 = 32'd1; 
32'd10376: dataIn2 = 32'd1; 
32'd10377: dataIn2 = 32'd1; 
32'd10378: dataIn2 = 32'd1; 
32'd10379: dataIn2 = 32'd0; 
32'd10380: dataIn2 = 32'd0; 
32'd10381: dataIn2 = 32'd0; 
32'd10382: dataIn2 = 32'd0; 
32'd10383: dataIn2 = 32'd1; 
32'd10384: dataIn2 = 32'd0; 
32'd10385: dataIn2 = 32'd1; 
32'd10386: dataIn2 = 32'd1; 
32'd10387: dataIn2 = 32'd1; 
32'd10388: dataIn2 = 32'd1; 
32'd10389: dataIn2 = 32'd0; 
32'd10390: dataIn2 = 32'd0; 
32'd10391: dataIn2 = 32'd0; 
32'd10392: dataIn2 = 32'd0; 
32'd10393: dataIn2 = 32'd1; 
32'd10394: dataIn2 = 32'd1; 
32'd10395: dataIn2 = 32'd0; 
32'd10396: dataIn2 = 32'd0; 
32'd10397: dataIn2 = 32'd0; 
32'd10398: dataIn2 = 32'd1; 
32'd10399: dataIn2 = 32'd0; 
32'd10400: dataIn2 = 32'd0; 
32'd10401: dataIn2 = 32'd1; 
32'd10402: dataIn2 = 32'd1; 
32'd10403: dataIn2 = 32'd1; 
32'd10404: dataIn2 = 32'd0; 
32'd10405: dataIn2 = 32'd1; 
32'd10406: dataIn2 = 32'd1; 
32'd10407: dataIn2 = 32'd0; 
32'd10408: dataIn2 = 32'd1; 
32'd10409: dataIn2 = 32'd0; 
32'd10410: dataIn2 = 32'd0; 
32'd10411: dataIn2 = 32'd0; 
32'd10412: dataIn2 = 32'd0; 
32'd10413: dataIn2 = 32'd1; 
32'd10414: dataIn2 = 32'd0; 
32'd10415: dataIn2 = 32'd1; 
32'd10416: dataIn2 = 32'd0; 
32'd10417: dataIn2 = 32'd1; 
32'd10418: dataIn2 = 32'd0; 
32'd10419: dataIn2 = 32'd0; 
32'd10420: dataIn2 = 32'd0; 
32'd10421: dataIn2 = 32'd1; 
32'd10422: dataIn2 = 32'd1; 
32'd10423: dataIn2 = 32'd1; 
32'd10424: dataIn2 = 32'd0; 
32'd10425: dataIn2 = 32'd1; 
32'd10426: dataIn2 = 32'd1; 
32'd10427: dataIn2 = 32'd1; 
32'd10428: dataIn2 = 32'd0; 
32'd10429: dataIn2 = 32'd1; 
32'd10430: dataIn2 = 32'd1; 
32'd10431: dataIn2 = 32'd0; 
32'd10432: dataIn2 = 32'd1; 
32'd10433: dataIn2 = 32'd1; 
32'd10434: dataIn2 = 32'd1; 
32'd10435: dataIn2 = 32'd1; 
32'd10436: dataIn2 = 32'd1; 
32'd10437: dataIn2 = 32'd0; 
32'd10438: dataIn2 = 32'd0; 
32'd10439: dataIn2 = 32'd1; 
32'd10440: dataIn2 = 32'd0; 
32'd10441: dataIn2 = 32'd1; 
32'd10442: dataIn2 = 32'd0; 
32'd10443: dataIn2 = 32'd0; 
32'd10444: dataIn2 = 32'd1; 
32'd10445: dataIn2 = 32'd1; 
32'd10446: dataIn2 = 32'd1; 
32'd10447: dataIn2 = 32'd1; 
32'd10448: dataIn2 = 32'd1; 
32'd10449: dataIn2 = 32'd0; 
32'd10450: dataIn2 = 32'd1; 
32'd10451: dataIn2 = 32'd1; 
32'd10452: dataIn2 = 32'd0; 
32'd10453: dataIn2 = 32'd0; 
32'd10454: dataIn2 = 32'd0; 
32'd10455: dataIn2 = 32'd1; 
32'd10456: dataIn2 = 32'd0; 
32'd10457: dataIn2 = 32'd0; 
32'd10458: dataIn2 = 32'd0; 
32'd10459: dataIn2 = 32'd0; 
32'd10460: dataIn2 = 32'd0; 
32'd10461: dataIn2 = 32'd0; 
32'd10462: dataIn2 = 32'd0; 
32'd10463: dataIn2 = 32'd0; 
32'd10464: dataIn2 = 32'd0; 
32'd10465: dataIn2 = 32'd0; 
32'd10466: dataIn2 = 32'd0; 
32'd10467: dataIn2 = 32'd0; 
32'd10468: dataIn2 = 32'd0; 
32'd10469: dataIn2 = 32'd0; 
32'd10470: dataIn2 = 32'd1; 
32'd10471: dataIn2 = 32'd0; 
32'd10472: dataIn2 = 32'd1; 
32'd10473: dataIn2 = 32'd0; 
32'd10474: dataIn2 = 32'd1; 
32'd10475: dataIn2 = 32'd1; 
32'd10476: dataIn2 = 32'd0; 
32'd10477: dataIn2 = 32'd1; 
32'd10478: dataIn2 = 32'd1; 
32'd10479: dataIn2 = 32'd1; 
32'd10480: dataIn2 = 32'd0; 
32'd10481: dataIn2 = 32'd1; 
32'd10482: dataIn2 = 32'd0; 
32'd10483: dataIn2 = 32'd1; 
32'd10484: dataIn2 = 32'd1; 
32'd10485: dataIn2 = 32'd0; 
32'd10486: dataIn2 = 32'd0; 
32'd10487: dataIn2 = 32'd1; 
32'd10488: dataIn2 = 32'd1; 
32'd10489: dataIn2 = 32'd1; 
32'd10490: dataIn2 = 32'd0; 
32'd10491: dataIn2 = 32'd1; 
32'd10492: dataIn2 = 32'd0; 
32'd10493: dataIn2 = 32'd0; 
32'd10494: dataIn2 = 32'd1; 
32'd10495: dataIn2 = 32'd1; 
32'd10496: dataIn2 = 32'd1; 
32'd10497: dataIn2 = 32'd1; 
32'd10498: dataIn2 = 32'd1; 
32'd10499: dataIn2 = 32'd0; 
32'd10500: dataIn2 = 32'd1; 
32'd10501: dataIn2 = 32'd1; 
32'd10502: dataIn2 = 32'd1; 
32'd10503: dataIn2 = 32'd1; 
32'd10504: dataIn2 = 32'd0; 
32'd10505: dataIn2 = 32'd1; 
32'd10506: dataIn2 = 32'd1; 
32'd10507: dataIn2 = 32'd1; 
32'd10508: dataIn2 = 32'd0; 
32'd10509: dataIn2 = 32'd0; 
32'd10510: dataIn2 = 32'd0; 
32'd10511: dataIn2 = 32'd1; 
32'd10512: dataIn2 = 32'd1; 
32'd10513: dataIn2 = 32'd0; 
32'd10514: dataIn2 = 32'd1; 
32'd10515: dataIn2 = 32'd0; 
32'd10516: dataIn2 = 32'd1; 
32'd10517: dataIn2 = 32'd1; 
32'd10518: dataIn2 = 32'd0; 
32'd10519: dataIn2 = 32'd0; 
32'd10520: dataIn2 = 32'd1; 
32'd10521: dataIn2 = 32'd1; 
32'd10522: dataIn2 = 32'd0; 
32'd10523: dataIn2 = 32'd0; 
32'd10524: dataIn2 = 32'd0; 
32'd10525: dataIn2 = 32'd0; 
32'd10526: dataIn2 = 32'd1; 
32'd10527: dataIn2 = 32'd0; 
32'd10528: dataIn2 = 32'd1; 
32'd10529: dataIn2 = 32'd1; 
32'd10530: dataIn2 = 32'd0; 
32'd10531: dataIn2 = 32'd1; 
32'd10532: dataIn2 = 32'd1; 
32'd10533: dataIn2 = 32'd0; 
32'd10534: dataIn2 = 32'd1; 
32'd10535: dataIn2 = 32'd1; 
32'd10536: dataIn2 = 32'd0; 
32'd10537: dataIn2 = 32'd0; 
32'd10538: dataIn2 = 32'd0; 
32'd10539: dataIn2 = 32'd0; 
32'd10540: dataIn2 = 32'd1; 
32'd10541: dataIn2 = 32'd0; 
32'd10542: dataIn2 = 32'd1; 
32'd10543: dataIn2 = 32'd1; 
32'd10544: dataIn2 = 32'd0; 
32'd10545: dataIn2 = 32'd1; 
32'd10546: dataIn2 = 32'd1; 
32'd10547: dataIn2 = 32'd1; 
32'd10548: dataIn2 = 32'd1; 
32'd10549: dataIn2 = 32'd0; 
32'd10550: dataIn2 = 32'd0; 
32'd10551: dataIn2 = 32'd1; 
32'd10552: dataIn2 = 32'd1; 
32'd10553: dataIn2 = 32'd0; 
32'd10554: dataIn2 = 32'd1; 
32'd10555: dataIn2 = 32'd1; 
32'd10556: dataIn2 = 32'd0; 
32'd10557: dataIn2 = 32'd1; 
32'd10558: dataIn2 = 32'd1; 
32'd10559: dataIn2 = 32'd0; 
32'd10560: dataIn2 = 32'd0; 
32'd10561: dataIn2 = 32'd1; 
32'd10562: dataIn2 = 32'd0; 
32'd10563: dataIn2 = 32'd0; 
32'd10564: dataIn2 = 32'd1; 
32'd10565: dataIn2 = 32'd1; 
32'd10566: dataIn2 = 32'd0; 
32'd10567: dataIn2 = 32'd0; 
32'd10568: dataIn2 = 32'd0; 
32'd10569: dataIn2 = 32'd1; 
32'd10570: dataIn2 = 32'd0; 
32'd10571: dataIn2 = 32'd0; 
32'd10572: dataIn2 = 32'd0; 
32'd10573: dataIn2 = 32'd1; 
32'd10574: dataIn2 = 32'd1; 
32'd10575: dataIn2 = 32'd1; 
32'd10576: dataIn2 = 32'd0; 
32'd10577: dataIn2 = 32'd0; 
32'd10578: dataIn2 = 32'd1; 
32'd10579: dataIn2 = 32'd1; 
32'd10580: dataIn2 = 32'd1; 
32'd10581: dataIn2 = 32'd1; 
32'd10582: dataIn2 = 32'd1; 
32'd10583: dataIn2 = 32'd1; 
32'd10584: dataIn2 = 32'd1; 
32'd10585: dataIn2 = 32'd1; 
32'd10586: dataIn2 = 32'd1; 
32'd10587: dataIn2 = 32'd0; 
32'd10588: dataIn2 = 32'd0; 
32'd10589: dataIn2 = 32'd1; 
32'd10590: dataIn2 = 32'd1; 
32'd10591: dataIn2 = 32'd1; 
32'd10592: dataIn2 = 32'd1; 
32'd10593: dataIn2 = 32'd1; 
32'd10594: dataIn2 = 32'd0; 
32'd10595: dataIn2 = 32'd1; 
32'd10596: dataIn2 = 32'd0; 
32'd10597: dataIn2 = 32'd0; 
32'd10598: dataIn2 = 32'd0; 
32'd10599: dataIn2 = 32'd1; 
32'd10600: dataIn2 = 32'd1; 
32'd10601: dataIn2 = 32'd0; 
32'd10602: dataIn2 = 32'd1; 
32'd10603: dataIn2 = 32'd1; 
32'd10604: dataIn2 = 32'd1; 
32'd10605: dataIn2 = 32'd1; 
32'd10606: dataIn2 = 32'd0; 
32'd10607: dataIn2 = 32'd1; 
32'd10608: dataIn2 = 32'd0; 
32'd10609: dataIn2 = 32'd0; 
32'd10610: dataIn2 = 32'd1; 
32'd10611: dataIn2 = 32'd1; 
32'd10612: dataIn2 = 32'd1; 
32'd10613: dataIn2 = 32'd0; 
32'd10614: dataIn2 = 32'd0; 
32'd10615: dataIn2 = 32'd0; 
32'd10616: dataIn2 = 32'd0; 
32'd10617: dataIn2 = 32'd1; 
32'd10618: dataIn2 = 32'd1; 
32'd10619: dataIn2 = 32'd0; 
32'd10620: dataIn2 = 32'd0; 
32'd10621: dataIn2 = 32'd0; 
32'd10622: dataIn2 = 32'd0; 
32'd10623: dataIn2 = 32'd0; 
32'd10624: dataIn2 = 32'd0; 
32'd10625: dataIn2 = 32'd0; 
32'd10626: dataIn2 = 32'd0; 
32'd10627: dataIn2 = 32'd0; 
32'd10628: dataIn2 = 32'd1; 
32'd10629: dataIn2 = 32'd0; 
32'd10630: dataIn2 = 32'd0; 
32'd10631: dataIn2 = 32'd1; 
32'd10632: dataIn2 = 32'd1; 
32'd10633: dataIn2 = 32'd1; 
32'd10634: dataIn2 = 32'd1; 
32'd10635: dataIn2 = 32'd1; 
32'd10636: dataIn2 = 32'd1; 
32'd10637: dataIn2 = 32'd1; 
32'd10638: dataIn2 = 32'd0; 
32'd10639: dataIn2 = 32'd0; 
32'd10640: dataIn2 = 32'd0; 
32'd10641: dataIn2 = 32'd1; 
32'd10642: dataIn2 = 32'd1; 
32'd10643: dataIn2 = 32'd1; 
32'd10644: dataIn2 = 32'd1; 
32'd10645: dataIn2 = 32'd0; 
32'd10646: dataIn2 = 32'd0; 
32'd10647: dataIn2 = 32'd1; 
32'd10648: dataIn2 = 32'd1; 
32'd10649: dataIn2 = 32'd0; 
32'd10650: dataIn2 = 32'd1; 
32'd10651: dataIn2 = 32'd1; 
32'd10652: dataIn2 = 32'd0; 
32'd10653: dataIn2 = 32'd0; 
32'd10654: dataIn2 = 32'd0; 
32'd10655: dataIn2 = 32'd1; 
32'd10656: dataIn2 = 32'd1; 
32'd10657: dataIn2 = 32'd1; 
32'd10658: dataIn2 = 32'd0; 
32'd10659: dataIn2 = 32'd1; 
32'd10660: dataIn2 = 32'd1; 
32'd10661: dataIn2 = 32'd0; 
32'd10662: dataIn2 = 32'd1; 
32'd10663: dataIn2 = 32'd0; 
32'd10664: dataIn2 = 32'd0; 
32'd10665: dataIn2 = 32'd0; 
32'd10666: dataIn2 = 32'd0; 
32'd10667: dataIn2 = 32'd1; 
32'd10668: dataIn2 = 32'd0; 
32'd10669: dataIn2 = 32'd1; 
32'd10670: dataIn2 = 32'd0; 
32'd10671: dataIn2 = 32'd1; 
32'd10672: dataIn2 = 32'd1; 
32'd10673: dataIn2 = 32'd1; 
32'd10674: dataIn2 = 32'd1; 
32'd10675: dataIn2 = 32'd0; 
32'd10676: dataIn2 = 32'd1; 
32'd10677: dataIn2 = 32'd1; 
32'd10678: dataIn2 = 32'd0; 
32'd10679: dataIn2 = 32'd0; 
32'd10680: dataIn2 = 32'd0; 
32'd10681: dataIn2 = 32'd0; 
32'd10682: dataIn2 = 32'd0; 
32'd10683: dataIn2 = 32'd1; 
32'd10684: dataIn2 = 32'd1; 
32'd10685: dataIn2 = 32'd1; 
32'd10686: dataIn2 = 32'd1; 
32'd10687: dataIn2 = 32'd0; 
32'd10688: dataIn2 = 32'd0; 
32'd10689: dataIn2 = 32'd1; 
32'd10690: dataIn2 = 32'd0; 
32'd10691: dataIn2 = 32'd1; 
32'd10692: dataIn2 = 32'd1; 
32'd10693: dataIn2 = 32'd0; 
32'd10694: dataIn2 = 32'd1; 
32'd10695: dataIn2 = 32'd0; 
32'd10696: dataIn2 = 32'd0; 
32'd10697: dataIn2 = 32'd1; 
32'd10698: dataIn2 = 32'd1; 
32'd10699: dataIn2 = 32'd1; 
32'd10700: dataIn2 = 32'd1; 
32'd10701: dataIn2 = 32'd1; 
32'd10702: dataIn2 = 32'd0; 
32'd10703: dataIn2 = 32'd1; 
32'd10704: dataIn2 = 32'd1; 
32'd10705: dataIn2 = 32'd0; 
32'd10706: dataIn2 = 32'd1; 
32'd10707: dataIn2 = 32'd0; 
32'd10708: dataIn2 = 32'd1; 
32'd10709: dataIn2 = 32'd1; 
32'd10710: dataIn2 = 32'd1; 
32'd10711: dataIn2 = 32'd0; 
32'd10712: dataIn2 = 32'd0; 
32'd10713: dataIn2 = 32'd1; 
32'd10714: dataIn2 = 32'd0; 
32'd10715: dataIn2 = 32'd0; 
32'd10716: dataIn2 = 32'd1; 
32'd10717: dataIn2 = 32'd0; 
32'd10718: dataIn2 = 32'd1; 
32'd10719: dataIn2 = 32'd0; 
32'd10720: dataIn2 = 32'd0; 
32'd10721: dataIn2 = 32'd1; 
32'd10722: dataIn2 = 32'd0; 
32'd10723: dataIn2 = 32'd0; 
32'd10724: dataIn2 = 32'd0; 
32'd10725: dataIn2 = 32'd1; 
32'd10726: dataIn2 = 32'd0; 
32'd10727: dataIn2 = 32'd1; 
32'd10728: dataIn2 = 32'd0; 
32'd10729: dataIn2 = 32'd0; 
32'd10730: dataIn2 = 32'd1; 
32'd10731: dataIn2 = 32'd0; 
32'd10732: dataIn2 = 32'd1; 
32'd10733: dataIn2 = 32'd0; 
32'd10734: dataIn2 = 32'd1; 
32'd10735: dataIn2 = 32'd1; 
32'd10736: dataIn2 = 32'd0; 
32'd10737: dataIn2 = 32'd1; 
32'd10738: dataIn2 = 32'd0; 
32'd10739: dataIn2 = 32'd1; 
32'd10740: dataIn2 = 32'd1; 
32'd10741: dataIn2 = 32'd0; 
32'd10742: dataIn2 = 32'd1; 
32'd10743: dataIn2 = 32'd1; 
32'd10744: dataIn2 = 32'd1; 
32'd10745: dataIn2 = 32'd0; 
32'd10746: dataIn2 = 32'd0; 
32'd10747: dataIn2 = 32'd0; 
32'd10748: dataIn2 = 32'd0; 
32'd10749: dataIn2 = 32'd0; 
32'd10750: dataIn2 = 32'd0; 
32'd10751: dataIn2 = 32'd1; 
32'd10752: dataIn2 = 32'd0; 
32'd10753: dataIn2 = 32'd0; 
32'd10754: dataIn2 = 32'd1; 
32'd10755: dataIn2 = 32'd0; 
32'd10756: dataIn2 = 32'd0; 
32'd10757: dataIn2 = 32'd1; 
32'd10758: dataIn2 = 32'd1; 
32'd10759: dataIn2 = 32'd0; 
32'd10760: dataIn2 = 32'd1; 
32'd10761: dataIn2 = 32'd0; 
32'd10762: dataIn2 = 32'd1; 
32'd10763: dataIn2 = 32'd1; 
32'd10764: dataIn2 = 32'd0; 
32'd10765: dataIn2 = 32'd1; 
32'd10766: dataIn2 = 32'd1; 
32'd10767: dataIn2 = 32'd0; 
32'd10768: dataIn2 = 32'd0; 
32'd10769: dataIn2 = 32'd1; 
32'd10770: dataIn2 = 32'd0; 
32'd10771: dataIn2 = 32'd1; 
32'd10772: dataIn2 = 32'd1; 
32'd10773: dataIn2 = 32'd1; 
32'd10774: dataIn2 = 32'd0; 
32'd10775: dataIn2 = 32'd0; 
32'd10776: dataIn2 = 32'd0; 
32'd10777: dataIn2 = 32'd1; 
32'd10778: dataIn2 = 32'd0; 
32'd10779: dataIn2 = 32'd0; 
32'd10780: dataIn2 = 32'd0; 
32'd10781: dataIn2 = 32'd0; 
32'd10782: dataIn2 = 32'd0; 
32'd10783: dataIn2 = 32'd1; 
32'd10784: dataIn2 = 32'd1; 
32'd10785: dataIn2 = 32'd1; 
32'd10786: dataIn2 = 32'd0; 
32'd10787: dataIn2 = 32'd0; 
32'd10788: dataIn2 = 32'd0; 
32'd10789: dataIn2 = 32'd1; 
32'd10790: dataIn2 = 32'd0; 
32'd10791: dataIn2 = 32'd1; 
32'd10792: dataIn2 = 32'd0; 
32'd10793: dataIn2 = 32'd1; 
32'd10794: dataIn2 = 32'd0; 
32'd10795: dataIn2 = 32'd0; 
32'd10796: dataIn2 = 32'd0; 
32'd10797: dataIn2 = 32'd1; 
32'd10798: dataIn2 = 32'd0; 
32'd10799: dataIn2 = 32'd0; 
32'd10800: dataIn2 = 32'd0; 
32'd10801: dataIn2 = 32'd0; 
32'd10802: dataIn2 = 32'd1; 
32'd10803: dataIn2 = 32'd0; 
32'd10804: dataIn2 = 32'd1; 
32'd10805: dataIn2 = 32'd1; 
32'd10806: dataIn2 = 32'd0; 
32'd10807: dataIn2 = 32'd1; 
32'd10808: dataIn2 = 32'd0; 
32'd10809: dataIn2 = 32'd1; 
32'd10810: dataIn2 = 32'd1; 
32'd10811: dataIn2 = 32'd0; 
32'd10812: dataIn2 = 32'd0; 
32'd10813: dataIn2 = 32'd1; 
32'd10814: dataIn2 = 32'd0; 
32'd10815: dataIn2 = 32'd0; 
32'd10816: dataIn2 = 32'd1; 
32'd10817: dataIn2 = 32'd0; 
32'd10818: dataIn2 = 32'd0; 
32'd10819: dataIn2 = 32'd0; 
32'd10820: dataIn2 = 32'd1; 
32'd10821: dataIn2 = 32'd1; 
32'd10822: dataIn2 = 32'd0; 
32'd10823: dataIn2 = 32'd1; 
32'd10824: dataIn2 = 32'd0; 
32'd10825: dataIn2 = 32'd1; 
32'd10826: dataIn2 = 32'd0; 
32'd10827: dataIn2 = 32'd1; 
32'd10828: dataIn2 = 32'd1; 
32'd10829: dataIn2 = 32'd0; 
32'd10830: dataIn2 = 32'd0; 
32'd10831: dataIn2 = 32'd0; 
32'd10832: dataIn2 = 32'd0; 
32'd10833: dataIn2 = 32'd1; 
32'd10834: dataIn2 = 32'd1; 
32'd10835: dataIn2 = 32'd0; 
32'd10836: dataIn2 = 32'd1; 
32'd10837: dataIn2 = 32'd0; 
32'd10838: dataIn2 = 32'd1; 
32'd10839: dataIn2 = 32'd0; 
32'd10840: dataIn2 = 32'd1; 
32'd10841: dataIn2 = 32'd0; 
32'd10842: dataIn2 = 32'd0; 
32'd10843: dataIn2 = 32'd1; 
32'd10844: dataIn2 = 32'd1; 
32'd10845: dataIn2 = 32'd0; 
32'd10846: dataIn2 = 32'd1; 
32'd10847: dataIn2 = 32'd0; 
32'd10848: dataIn2 = 32'd1; 
32'd10849: dataIn2 = 32'd0; 
32'd10850: dataIn2 = 32'd1; 
32'd10851: dataIn2 = 32'd1; 
32'd10852: dataIn2 = 32'd1; 
32'd10853: dataIn2 = 32'd1; 
32'd10854: dataIn2 = 32'd1; 
32'd10855: dataIn2 = 32'd0; 
32'd10856: dataIn2 = 32'd1; 
32'd10857: dataIn2 = 32'd1; 
32'd10858: dataIn2 = 32'd1; 
32'd10859: dataIn2 = 32'd0; 
32'd10860: dataIn2 = 32'd1; 
32'd10861: dataIn2 = 32'd1; 
32'd10862: dataIn2 = 32'd0; 
32'd10863: dataIn2 = 32'd0; 
32'd10864: dataIn2 = 32'd0; 
32'd10865: dataIn2 = 32'd0; 
32'd10866: dataIn2 = 32'd1; 
32'd10867: dataIn2 = 32'd1; 
32'd10868: dataIn2 = 32'd0; 
32'd10869: dataIn2 = 32'd1; 
32'd10870: dataIn2 = 32'd0; 
32'd10871: dataIn2 = 32'd0; 
32'd10872: dataIn2 = 32'd0; 
32'd10873: dataIn2 = 32'd0; 
32'd10874: dataIn2 = 32'd1; 
32'd10875: dataIn2 = 32'd1; 
32'd10876: dataIn2 = 32'd1; 
32'd10877: dataIn2 = 32'd0; 
32'd10878: dataIn2 = 32'd0; 
32'd10879: dataIn2 = 32'd1; 
32'd10880: dataIn2 = 32'd1; 
32'd10881: dataIn2 = 32'd0; 
32'd10882: dataIn2 = 32'd0; 
32'd10883: dataIn2 = 32'd1; 
32'd10884: dataIn2 = 32'd0; 
32'd10885: dataIn2 = 32'd0; 
32'd10886: dataIn2 = 32'd1; 
32'd10887: dataIn2 = 32'd0; 
32'd10888: dataIn2 = 32'd0; 
32'd10889: dataIn2 = 32'd0; 
32'd10890: dataIn2 = 32'd0; 
32'd10891: dataIn2 = 32'd1; 
32'd10892: dataIn2 = 32'd1; 
32'd10893: dataIn2 = 32'd0; 
32'd10894: dataIn2 = 32'd1; 
32'd10895: dataIn2 = 32'd0; 
32'd10896: dataIn2 = 32'd1; 
32'd10897: dataIn2 = 32'd1; 
32'd10898: dataIn2 = 32'd1; 
32'd10899: dataIn2 = 32'd1; 
32'd10900: dataIn2 = 32'd0; 
32'd10901: dataIn2 = 32'd0; 
32'd10902: dataIn2 = 32'd0; 
32'd10903: dataIn2 = 32'd0; 
32'd10904: dataIn2 = 32'd1; 
32'd10905: dataIn2 = 32'd0; 
32'd10906: dataIn2 = 32'd0; 
32'd10907: dataIn2 = 32'd0; 
32'd10908: dataIn2 = 32'd1; 
32'd10909: dataIn2 = 32'd1; 
32'd10910: dataIn2 = 32'd1; 
32'd10911: dataIn2 = 32'd1; 
32'd10912: dataIn2 = 32'd1; 
32'd10913: dataIn2 = 32'd0; 
32'd10914: dataIn2 = 32'd0; 
32'd10915: dataIn2 = 32'd1; 
32'd10916: dataIn2 = 32'd1; 
32'd10917: dataIn2 = 32'd0; 
32'd10918: dataIn2 = 32'd0; 
32'd10919: dataIn2 = 32'd0; 
32'd10920: dataIn2 = 32'd1; 
32'd10921: dataIn2 = 32'd0; 
32'd10922: dataIn2 = 32'd1; 
32'd10923: dataIn2 = 32'd1; 
32'd10924: dataIn2 = 32'd0; 
32'd10925: dataIn2 = 32'd1; 
32'd10926: dataIn2 = 32'd1; 
32'd10927: dataIn2 = 32'd1; 
32'd10928: dataIn2 = 32'd1; 
32'd10929: dataIn2 = 32'd1; 
32'd10930: dataIn2 = 32'd1; 
32'd10931: dataIn2 = 32'd1; 
32'd10932: dataIn2 = 32'd1; 
32'd10933: dataIn2 = 32'd1; 
32'd10934: dataIn2 = 32'd1; 
32'd10935: dataIn2 = 32'd0; 
32'd10936: dataIn2 = 32'd0; 
32'd10937: dataIn2 = 32'd1; 
32'd10938: dataIn2 = 32'd1; 
32'd10939: dataIn2 = 32'd0; 
32'd10940: dataIn2 = 32'd1; 
32'd10941: dataIn2 = 32'd0; 
32'd10942: dataIn2 = 32'd1; 
32'd10943: dataIn2 = 32'd1; 
32'd10944: dataIn2 = 32'd1; 
32'd10945: dataIn2 = 32'd1; 
32'd10946: dataIn2 = 32'd0; 
32'd10947: dataIn2 = 32'd1; 
32'd10948: dataIn2 = 32'd1; 
32'd10949: dataIn2 = 32'd0; 
32'd10950: dataIn2 = 32'd1; 
32'd10951: dataIn2 = 32'd0; 
32'd10952: dataIn2 = 32'd1; 
32'd10953: dataIn2 = 32'd0; 
32'd10954: dataIn2 = 32'd1; 
32'd10955: dataIn2 = 32'd1; 
32'd10956: dataIn2 = 32'd0; 
32'd10957: dataIn2 = 32'd0; 
32'd10958: dataIn2 = 32'd0; 
32'd10959: dataIn2 = 32'd1; 
32'd10960: dataIn2 = 32'd0; 
32'd10961: dataIn2 = 32'd1; 
32'd10962: dataIn2 = 32'd1; 
32'd10963: dataIn2 = 32'd0; 
32'd10964: dataIn2 = 32'd1; 
32'd10965: dataIn2 = 32'd0; 
32'd10966: dataIn2 = 32'd0; 
32'd10967: dataIn2 = 32'd1; 
32'd10968: dataIn2 = 32'd0; 
32'd10969: dataIn2 = 32'd0; 
32'd10970: dataIn2 = 32'd1; 
32'd10971: dataIn2 = 32'd1; 
32'd10972: dataIn2 = 32'd0; 
32'd10973: dataIn2 = 32'd0; 
32'd10974: dataIn2 = 32'd1; 
32'd10975: dataIn2 = 32'd1; 
32'd10976: dataIn2 = 32'd1; 
32'd10977: dataIn2 = 32'd0; 
32'd10978: dataIn2 = 32'd1; 
32'd10979: dataIn2 = 32'd1; 
32'd10980: dataIn2 = 32'd1; 
32'd10981: dataIn2 = 32'd1; 
32'd10982: dataIn2 = 32'd0; 
32'd10983: dataIn2 = 32'd0; 
32'd10984: dataIn2 = 32'd0; 
32'd10985: dataIn2 = 32'd1; 
32'd10986: dataIn2 = 32'd0; 
32'd10987: dataIn2 = 32'd0; 
32'd10988: dataIn2 = 32'd0; 
32'd10989: dataIn2 = 32'd1; 
32'd10990: dataIn2 = 32'd0; 
32'd10991: dataIn2 = 32'd1; 
32'd10992: dataIn2 = 32'd0; 
32'd10993: dataIn2 = 32'd1; 
32'd10994: dataIn2 = 32'd1; 
32'd10995: dataIn2 = 32'd1; 
32'd10996: dataIn2 = 32'd1; 
32'd10997: dataIn2 = 32'd0; 
32'd10998: dataIn2 = 32'd0; 
32'd10999: dataIn2 = 32'd1; 
32'd11000: dataIn2 = 32'd0; 
32'd11001: dataIn2 = 32'd0; 
32'd11002: dataIn2 = 32'd1; 
32'd11003: dataIn2 = 32'd1; 
32'd11004: dataIn2 = 32'd1; 
32'd11005: dataIn2 = 32'd1; 
32'd11006: dataIn2 = 32'd1; 
32'd11007: dataIn2 = 32'd0; 
32'd11008: dataIn2 = 32'd1; 
32'd11009: dataIn2 = 32'd0; 
32'd11010: dataIn2 = 32'd1; 
32'd11011: dataIn2 = 32'd0; 
32'd11012: dataIn2 = 32'd1; 
32'd11013: dataIn2 = 32'd1; 
32'd11014: dataIn2 = 32'd1; 
32'd11015: dataIn2 = 32'd1; 
32'd11016: dataIn2 = 32'd1; 
32'd11017: dataIn2 = 32'd1; 
32'd11018: dataIn2 = 32'd1; 
32'd11019: dataIn2 = 32'd1; 
32'd11020: dataIn2 = 32'd1; 
32'd11021: dataIn2 = 32'd0; 
32'd11022: dataIn2 = 32'd1; 
32'd11023: dataIn2 = 32'd1; 
32'd11024: dataIn2 = 32'd1; 
32'd11025: dataIn2 = 32'd0; 
32'd11026: dataIn2 = 32'd1; 
32'd11027: dataIn2 = 32'd1; 
32'd11028: dataIn2 = 32'd1; 
32'd11029: dataIn2 = 32'd1; 
32'd11030: dataIn2 = 32'd1; 
32'd11031: dataIn2 = 32'd1; 
32'd11032: dataIn2 = 32'd1; 
32'd11033: dataIn2 = 32'd1; 
32'd11034: dataIn2 = 32'd1; 
32'd11035: dataIn2 = 32'd1; 
32'd11036: dataIn2 = 32'd0; 
32'd11037: dataIn2 = 32'd0; 
32'd11038: dataIn2 = 32'd0; 
32'd11039: dataIn2 = 32'd0; 
32'd11040: dataIn2 = 32'd1; 
32'd11041: dataIn2 = 32'd1; 
32'd11042: dataIn2 = 32'd1; 
32'd11043: dataIn2 = 32'd1; 
32'd11044: dataIn2 = 32'd0; 
32'd11045: dataIn2 = 32'd1; 
32'd11046: dataIn2 = 32'd0; 
32'd11047: dataIn2 = 32'd0; 
32'd11048: dataIn2 = 32'd0; 
32'd11049: dataIn2 = 32'd1; 
32'd11050: dataIn2 = 32'd1; 
32'd11051: dataIn2 = 32'd0; 
32'd11052: dataIn2 = 32'd1; 
32'd11053: dataIn2 = 32'd0; 
32'd11054: dataIn2 = 32'd0; 
32'd11055: dataIn2 = 32'd1; 
32'd11056: dataIn2 = 32'd0; 
32'd11057: dataIn2 = 32'd0; 
32'd11058: dataIn2 = 32'd0; 
32'd11059: dataIn2 = 32'd0; 
32'd11060: dataIn2 = 32'd0; 
32'd11061: dataIn2 = 32'd0; 
32'd11062: dataIn2 = 32'd1; 
32'd11063: dataIn2 = 32'd1; 
32'd11064: dataIn2 = 32'd1; 
32'd11065: dataIn2 = 32'd0; 
32'd11066: dataIn2 = 32'd0; 
32'd11067: dataIn2 = 32'd0; 
32'd11068: dataIn2 = 32'd1; 
32'd11069: dataIn2 = 32'd0; 
32'd11070: dataIn2 = 32'd1; 
32'd11071: dataIn2 = 32'd1; 
32'd11072: dataIn2 = 32'd0; 
32'd11073: dataIn2 = 32'd1; 
32'd11074: dataIn2 = 32'd1; 
32'd11075: dataIn2 = 32'd0; 
32'd11076: dataIn2 = 32'd0; 
32'd11077: dataIn2 = 32'd1; 
32'd11078: dataIn2 = 32'd0; 
32'd11079: dataIn2 = 32'd0; 
32'd11080: dataIn2 = 32'd0; 
32'd11081: dataIn2 = 32'd0; 
32'd11082: dataIn2 = 32'd0; 
32'd11083: dataIn2 = 32'd0; 
32'd11084: dataIn2 = 32'd0; 
32'd11085: dataIn2 = 32'd1; 
32'd11086: dataIn2 = 32'd0; 
32'd11087: dataIn2 = 32'd0; 
32'd11088: dataIn2 = 32'd1; 
32'd11089: dataIn2 = 32'd0; 
32'd11090: dataIn2 = 32'd1; 
32'd11091: dataIn2 = 32'd1; 
32'd11092: dataIn2 = 32'd1; 
32'd11093: dataIn2 = 32'd0; 
32'd11094: dataIn2 = 32'd0; 
32'd11095: dataIn2 = 32'd0; 
32'd11096: dataIn2 = 32'd1; 
32'd11097: dataIn2 = 32'd1; 
32'd11098: dataIn2 = 32'd1; 
32'd11099: dataIn2 = 32'd0; 
32'd11100: dataIn2 = 32'd0; 
32'd11101: dataIn2 = 32'd0; 
32'd11102: dataIn2 = 32'd1; 
32'd11103: dataIn2 = 32'd1; 
32'd11104: dataIn2 = 32'd0; 
32'd11105: dataIn2 = 32'd1; 
32'd11106: dataIn2 = 32'd0; 
32'd11107: dataIn2 = 32'd0; 
32'd11108: dataIn2 = 32'd1; 
32'd11109: dataIn2 = 32'd1; 
32'd11110: dataIn2 = 32'd0; 
32'd11111: dataIn2 = 32'd0; 
32'd11112: dataIn2 = 32'd1; 
32'd11113: dataIn2 = 32'd0; 
32'd11114: dataIn2 = 32'd0; 
32'd11115: dataIn2 = 32'd1; 
32'd11116: dataIn2 = 32'd0; 
32'd11117: dataIn2 = 32'd1; 
32'd11118: dataIn2 = 32'd0; 
32'd11119: dataIn2 = 32'd0; 
32'd11120: dataIn2 = 32'd0; 
32'd11121: dataIn2 = 32'd1; 
32'd11122: dataIn2 = 32'd0; 
32'd11123: dataIn2 = 32'd0; 
32'd11124: dataIn2 = 32'd1; 
32'd11125: dataIn2 = 32'd1; 
32'd11126: dataIn2 = 32'd1; 
32'd11127: dataIn2 = 32'd1; 
32'd11128: dataIn2 = 32'd0; 
32'd11129: dataIn2 = 32'd1; 
32'd11130: dataIn2 = 32'd0; 
32'd11131: dataIn2 = 32'd0; 
32'd11132: dataIn2 = 32'd1; 
32'd11133: dataIn2 = 32'd1; 
32'd11134: dataIn2 = 32'd1; 
32'd11135: dataIn2 = 32'd0; 
32'd11136: dataIn2 = 32'd0; 
32'd11137: dataIn2 = 32'd0; 
32'd11138: dataIn2 = 32'd1; 
32'd11139: dataIn2 = 32'd0; 
32'd11140: dataIn2 = 32'd0; 
32'd11141: dataIn2 = 32'd0; 
32'd11142: dataIn2 = 32'd0; 
32'd11143: dataIn2 = 32'd1; 
32'd11144: dataIn2 = 32'd1; 
32'd11145: dataIn2 = 32'd0; 
32'd11146: dataIn2 = 32'd0; 
32'd11147: dataIn2 = 32'd0; 
32'd11148: dataIn2 = 32'd0; 
32'd11149: dataIn2 = 32'd1; 
32'd11150: dataIn2 = 32'd1; 
32'd11151: dataIn2 = 32'd0; 
32'd11152: dataIn2 = 32'd1; 
32'd11153: dataIn2 = 32'd0; 
32'd11154: dataIn2 = 32'd1; 
32'd11155: dataIn2 = 32'd1; 
32'd11156: dataIn2 = 32'd0; 
32'd11157: dataIn2 = 32'd1; 
32'd11158: dataIn2 = 32'd0; 
32'd11159: dataIn2 = 32'd1; 
32'd11160: dataIn2 = 32'd1; 
32'd11161: dataIn2 = 32'd1; 
32'd11162: dataIn2 = 32'd0; 
32'd11163: dataIn2 = 32'd0; 
32'd11164: dataIn2 = 32'd0; 
32'd11165: dataIn2 = 32'd1; 
32'd11166: dataIn2 = 32'd0; 
32'd11167: dataIn2 = 32'd0; 
32'd11168: dataIn2 = 32'd1; 
32'd11169: dataIn2 = 32'd1; 
32'd11170: dataIn2 = 32'd0; 
32'd11171: dataIn2 = 32'd1; 
32'd11172: dataIn2 = 32'd0; 
32'd11173: dataIn2 = 32'd0; 
32'd11174: dataIn2 = 32'd0; 
32'd11175: dataIn2 = 32'd1; 
32'd11176: dataIn2 = 32'd0; 
32'd11177: dataIn2 = 32'd1; 
32'd11178: dataIn2 = 32'd1; 
32'd11179: dataIn2 = 32'd0; 
32'd11180: dataIn2 = 32'd0; 
32'd11181: dataIn2 = 32'd0; 
32'd11182: dataIn2 = 32'd0; 
32'd11183: dataIn2 = 32'd1; 
32'd11184: dataIn2 = 32'd0; 
32'd11185: dataIn2 = 32'd1; 
32'd11186: dataIn2 = 32'd0; 
32'd11187: dataIn2 = 32'd0; 
32'd11188: dataIn2 = 32'd0; 
32'd11189: dataIn2 = 32'd0; 
32'd11190: dataIn2 = 32'd1; 
32'd11191: dataIn2 = 32'd0; 
32'd11192: dataIn2 = 32'd0; 
32'd11193: dataIn2 = 32'd1; 
32'd11194: dataIn2 = 32'd1; 
32'd11195: dataIn2 = 32'd1; 
32'd11196: dataIn2 = 32'd0; 
32'd11197: dataIn2 = 32'd1; 
32'd11198: dataIn2 = 32'd0; 
32'd11199: dataIn2 = 32'd1; 
32'd11200: dataIn2 = 32'd1; 
32'd11201: dataIn2 = 32'd0; 
32'd11202: dataIn2 = 32'd1; 
32'd11203: dataIn2 = 32'd0; 
32'd11204: dataIn2 = 32'd1; 
32'd11205: dataIn2 = 32'd1; 
32'd11206: dataIn2 = 32'd0; 
32'd11207: dataIn2 = 32'd0; 
32'd11208: dataIn2 = 32'd1; 
32'd11209: dataIn2 = 32'd1; 
32'd11210: dataIn2 = 32'd0; 
32'd11211: dataIn2 = 32'd0; 
32'd11212: dataIn2 = 32'd1; 
32'd11213: dataIn2 = 32'd1; 
32'd11214: dataIn2 = 32'd1; 
32'd11215: dataIn2 = 32'd0; 
32'd11216: dataIn2 = 32'd1; 
32'd11217: dataIn2 = 32'd0; 
32'd11218: dataIn2 = 32'd0; 
32'd11219: dataIn2 = 32'd1; 
32'd11220: dataIn2 = 32'd1; 
32'd11221: dataIn2 = 32'd1; 
32'd11222: dataIn2 = 32'd0; 
32'd11223: dataIn2 = 32'd1; 
32'd11224: dataIn2 = 32'd0; 
32'd11225: dataIn2 = 32'd1; 
32'd11226: dataIn2 = 32'd0; 
32'd11227: dataIn2 = 32'd1; 
32'd11228: dataIn2 = 32'd0; 
32'd11229: dataIn2 = 32'd0; 
32'd11230: dataIn2 = 32'd0; 
32'd11231: dataIn2 = 32'd0; 
32'd11232: dataIn2 = 32'd0; 
32'd11233: dataIn2 = 32'd0; 
32'd11234: dataIn2 = 32'd0; 
32'd11235: dataIn2 = 32'd1; 
32'd11236: dataIn2 = 32'd1; 
32'd11237: dataIn2 = 32'd0; 
32'd11238: dataIn2 = 32'd0; 
32'd11239: dataIn2 = 32'd1; 
32'd11240: dataIn2 = 32'd1; 
32'd11241: dataIn2 = 32'd0; 
32'd11242: dataIn2 = 32'd0; 
32'd11243: dataIn2 = 32'd0; 
32'd11244: dataIn2 = 32'd1; 
32'd11245: dataIn2 = 32'd0; 
32'd11246: dataIn2 = 32'd0; 
32'd11247: dataIn2 = 32'd1; 
32'd11248: dataIn2 = 32'd0; 
32'd11249: dataIn2 = 32'd1; 
32'd11250: dataIn2 = 32'd0; 
32'd11251: dataIn2 = 32'd0; 
32'd11252: dataIn2 = 32'd1; 
32'd11253: dataIn2 = 32'd0; 
32'd11254: dataIn2 = 32'd1; 
32'd11255: dataIn2 = 32'd1; 
32'd11256: dataIn2 = 32'd0; 
32'd11257: dataIn2 = 32'd0; 
32'd11258: dataIn2 = 32'd1; 
32'd11259: dataIn2 = 32'd0; 
32'd11260: dataIn2 = 32'd0; 
32'd11261: dataIn2 = 32'd1; 
32'd11262: dataIn2 = 32'd0; 
32'd11263: dataIn2 = 32'd0; 
32'd11264: dataIn2 = 32'd1; 
32'd11265: dataIn2 = 32'd0; 
32'd11266: dataIn2 = 32'd0; 
32'd11267: dataIn2 = 32'd0; 
32'd11268: dataIn2 = 32'd0; 
32'd11269: dataIn2 = 32'd1; 
32'd11270: dataIn2 = 32'd1; 
32'd11271: dataIn2 = 32'd0; 
32'd11272: dataIn2 = 32'd0; 
32'd11273: dataIn2 = 32'd1; 
32'd11274: dataIn2 = 32'd1; 
32'd11275: dataIn2 = 32'd0; 
32'd11276: dataIn2 = 32'd0; 
32'd11277: dataIn2 = 32'd0; 
32'd11278: dataIn2 = 32'd0; 
32'd11279: dataIn2 = 32'd0; 
32'd11280: dataIn2 = 32'd1; 
32'd11281: dataIn2 = 32'd1; 
32'd11282: dataIn2 = 32'd0; 
32'd11283: dataIn2 = 32'd1; 
32'd11284: dataIn2 = 32'd0; 
32'd11285: dataIn2 = 32'd1; 
32'd11286: dataIn2 = 32'd1; 
32'd11287: dataIn2 = 32'd0; 
32'd11288: dataIn2 = 32'd0; 
32'd11289: dataIn2 = 32'd0; 
32'd11290: dataIn2 = 32'd0; 
32'd11291: dataIn2 = 32'd1; 
32'd11292: dataIn2 = 32'd0; 
32'd11293: dataIn2 = 32'd1; 
32'd11294: dataIn2 = 32'd0; 
32'd11295: dataIn2 = 32'd1; 
32'd11296: dataIn2 = 32'd1; 
32'd11297: dataIn2 = 32'd1; 
32'd11298: dataIn2 = 32'd1; 
32'd11299: dataIn2 = 32'd0; 
32'd11300: dataIn2 = 32'd0; 
32'd11301: dataIn2 = 32'd0; 
32'd11302: dataIn2 = 32'd0; 
32'd11303: dataIn2 = 32'd0; 
32'd11304: dataIn2 = 32'd1; 
32'd11305: dataIn2 = 32'd0; 
32'd11306: dataIn2 = 32'd0; 
32'd11307: dataIn2 = 32'd1; 
32'd11308: dataIn2 = 32'd0; 
32'd11309: dataIn2 = 32'd0; 
32'd11310: dataIn2 = 32'd0; 
32'd11311: dataIn2 = 32'd0; 
32'd11312: dataIn2 = 32'd1; 
32'd11313: dataIn2 = 32'd1; 
32'd11314: dataIn2 = 32'd1; 
32'd11315: dataIn2 = 32'd0; 
32'd11316: dataIn2 = 32'd1; 
32'd11317: dataIn2 = 32'd0; 
32'd11318: dataIn2 = 32'd0; 
32'd11319: dataIn2 = 32'd1; 
32'd11320: dataIn2 = 32'd0; 
32'd11321: dataIn2 = 32'd0; 
32'd11322: dataIn2 = 32'd1; 
32'd11323: dataIn2 = 32'd0; 
32'd11324: dataIn2 = 32'd1; 
32'd11325: dataIn2 = 32'd1; 
32'd11326: dataIn2 = 32'd0; 
32'd11327: dataIn2 = 32'd1; 
32'd11328: dataIn2 = 32'd1; 
32'd11329: dataIn2 = 32'd1; 
32'd11330: dataIn2 = 32'd0; 
32'd11331: dataIn2 = 32'd1; 
32'd11332: dataIn2 = 32'd1; 
32'd11333: dataIn2 = 32'd0; 
32'd11334: dataIn2 = 32'd1; 
32'd11335: dataIn2 = 32'd1; 
32'd11336: dataIn2 = 32'd1; 
32'd11337: dataIn2 = 32'd1; 
32'd11338: dataIn2 = 32'd1; 
32'd11339: dataIn2 = 32'd1; 
32'd11340: dataIn2 = 32'd0; 
32'd11341: dataIn2 = 32'd0; 
32'd11342: dataIn2 = 32'd1; 
32'd11343: dataIn2 = 32'd0; 
32'd11344: dataIn2 = 32'd0; 
32'd11345: dataIn2 = 32'd1; 
32'd11346: dataIn2 = 32'd0; 
32'd11347: dataIn2 = 32'd1; 
32'd11348: dataIn2 = 32'd0; 
32'd11349: dataIn2 = 32'd1; 
32'd11350: dataIn2 = 32'd1; 
32'd11351: dataIn2 = 32'd0; 
32'd11352: dataIn2 = 32'd0; 
32'd11353: dataIn2 = 32'd0; 
32'd11354: dataIn2 = 32'd0; 
32'd11355: dataIn2 = 32'd1; 
32'd11356: dataIn2 = 32'd0; 
32'd11357: dataIn2 = 32'd0; 
32'd11358: dataIn2 = 32'd1; 
32'd11359: dataIn2 = 32'd0; 
32'd11360: dataIn2 = 32'd0; 
32'd11361: dataIn2 = 32'd0; 
32'd11362: dataIn2 = 32'd1; 
32'd11363: dataIn2 = 32'd1; 
32'd11364: dataIn2 = 32'd1; 
32'd11365: dataIn2 = 32'd0; 
32'd11366: dataIn2 = 32'd0; 
32'd11367: dataIn2 = 32'd1; 
32'd11368: dataIn2 = 32'd0; 
32'd11369: dataIn2 = 32'd0; 
32'd11370: dataIn2 = 32'd0; 
32'd11371: dataIn2 = 32'd1; 
32'd11372: dataIn2 = 32'd0; 
32'd11373: dataIn2 = 32'd1; 
32'd11374: dataIn2 = 32'd1; 
32'd11375: dataIn2 = 32'd1; 
32'd11376: dataIn2 = 32'd1; 
32'd11377: dataIn2 = 32'd1; 
32'd11378: dataIn2 = 32'd1; 
32'd11379: dataIn2 = 32'd0; 
32'd11380: dataIn2 = 32'd0; 
32'd11381: dataIn2 = 32'd0; 
32'd11382: dataIn2 = 32'd1; 
32'd11383: dataIn2 = 32'd0; 
32'd11384: dataIn2 = 32'd0; 
32'd11385: dataIn2 = 32'd0; 
32'd11386: dataIn2 = 32'd0; 
32'd11387: dataIn2 = 32'd0; 
32'd11388: dataIn2 = 32'd1; 
32'd11389: dataIn2 = 32'd0; 
32'd11390: dataIn2 = 32'd0; 
32'd11391: dataIn2 = 32'd1; 
32'd11392: dataIn2 = 32'd1; 
32'd11393: dataIn2 = 32'd0; 
32'd11394: dataIn2 = 32'd0; 
32'd11395: dataIn2 = 32'd0; 
32'd11396: dataIn2 = 32'd0; 
32'd11397: dataIn2 = 32'd1; 
32'd11398: dataIn2 = 32'd1; 
32'd11399: dataIn2 = 32'd0; 
32'd11400: dataIn2 = 32'd1; 
32'd11401: dataIn2 = 32'd0; 
32'd11402: dataIn2 = 32'd0; 
32'd11403: dataIn2 = 32'd0; 
32'd11404: dataIn2 = 32'd0; 
32'd11405: dataIn2 = 32'd0; 
32'd11406: dataIn2 = 32'd1; 
32'd11407: dataIn2 = 32'd1; 
32'd11408: dataIn2 = 32'd1; 
32'd11409: dataIn2 = 32'd1; 
32'd11410: dataIn2 = 32'd1; 
32'd11411: dataIn2 = 32'd0; 
32'd11412: dataIn2 = 32'd0; 
32'd11413: dataIn2 = 32'd0; 
32'd11414: dataIn2 = 32'd0; 
32'd11415: dataIn2 = 32'd1; 
32'd11416: dataIn2 = 32'd1; 
32'd11417: dataIn2 = 32'd1; 
32'd11418: dataIn2 = 32'd0; 
32'd11419: dataIn2 = 32'd0; 
32'd11420: dataIn2 = 32'd0; 
32'd11421: dataIn2 = 32'd0; 
32'd11422: dataIn2 = 32'd1; 
32'd11423: dataIn2 = 32'd0; 
32'd11424: dataIn2 = 32'd1; 
32'd11425: dataIn2 = 32'd1; 
32'd11426: dataIn2 = 32'd1; 
32'd11427: dataIn2 = 32'd0; 
32'd11428: dataIn2 = 32'd0; 
32'd11429: dataIn2 = 32'd0; 
32'd11430: dataIn2 = 32'd1; 
32'd11431: dataIn2 = 32'd0; 
32'd11432: dataIn2 = 32'd0; 
32'd11433: dataIn2 = 32'd1; 
32'd11434: dataIn2 = 32'd1; 
32'd11435: dataIn2 = 32'd1; 
32'd11436: dataIn2 = 32'd0; 
32'd11437: dataIn2 = 32'd1; 
32'd11438: dataIn2 = 32'd1; 
32'd11439: dataIn2 = 32'd1; 
32'd11440: dataIn2 = 32'd1; 
32'd11441: dataIn2 = 32'd1; 
32'd11442: dataIn2 = 32'd1; 
32'd11443: dataIn2 = 32'd1; 
32'd11444: dataIn2 = 32'd1; 
32'd11445: dataIn2 = 32'd0; 
32'd11446: dataIn2 = 32'd1; 
32'd11447: dataIn2 = 32'd1; 
32'd11448: dataIn2 = 32'd1; 
32'd11449: dataIn2 = 32'd1; 
32'd11450: dataIn2 = 32'd0; 
32'd11451: dataIn2 = 32'd0; 
32'd11452: dataIn2 = 32'd0; 
32'd11453: dataIn2 = 32'd0; 
32'd11454: dataIn2 = 32'd1; 
32'd11455: dataIn2 = 32'd0; 
32'd11456: dataIn2 = 32'd0; 
32'd11457: dataIn2 = 32'd1; 
32'd11458: dataIn2 = 32'd0; 
32'd11459: dataIn2 = 32'd1; 
32'd11460: dataIn2 = 32'd0; 
32'd11461: dataIn2 = 32'd0; 
32'd11462: dataIn2 = 32'd1; 
32'd11463: dataIn2 = 32'd1; 
32'd11464: dataIn2 = 32'd0; 
32'd11465: dataIn2 = 32'd0; 
32'd11466: dataIn2 = 32'd0; 
32'd11467: dataIn2 = 32'd0; 
32'd11468: dataIn2 = 32'd1; 
32'd11469: dataIn2 = 32'd1; 
32'd11470: dataIn2 = 32'd1; 
32'd11471: dataIn2 = 32'd0; 
32'd11472: dataIn2 = 32'd1; 
32'd11473: dataIn2 = 32'd0; 
32'd11474: dataIn2 = 32'd1; 
32'd11475: dataIn2 = 32'd0; 
32'd11476: dataIn2 = 32'd1; 
32'd11477: dataIn2 = 32'd0; 
32'd11478: dataIn2 = 32'd1; 
32'd11479: dataIn2 = 32'd1; 
32'd11480: dataIn2 = 32'd1; 
32'd11481: dataIn2 = 32'd0; 
32'd11482: dataIn2 = 32'd0; 
32'd11483: dataIn2 = 32'd0; 
32'd11484: dataIn2 = 32'd0; 
32'd11485: dataIn2 = 32'd1; 
32'd11486: dataIn2 = 32'd1; 
32'd11487: dataIn2 = 32'd0; 
32'd11488: dataIn2 = 32'd1; 
32'd11489: dataIn2 = 32'd1; 
32'd11490: dataIn2 = 32'd0; 
32'd11491: dataIn2 = 32'd0; 
32'd11492: dataIn2 = 32'd1; 
32'd11493: dataIn2 = 32'd1; 
32'd11494: dataIn2 = 32'd1; 
32'd11495: dataIn2 = 32'd0; 
32'd11496: dataIn2 = 32'd0; 
32'd11497: dataIn2 = 32'd0; 
32'd11498: dataIn2 = 32'd1; 
32'd11499: dataIn2 = 32'd0; 
32'd11500: dataIn2 = 32'd1; 
32'd11501: dataIn2 = 32'd0; 
32'd11502: dataIn2 = 32'd1; 
32'd11503: dataIn2 = 32'd0; 
32'd11504: dataIn2 = 32'd0; 
32'd11505: dataIn2 = 32'd0; 
32'd11506: dataIn2 = 32'd1; 
32'd11507: dataIn2 = 32'd1; 
32'd11508: dataIn2 = 32'd0; 
32'd11509: dataIn2 = 32'd1; 
32'd11510: dataIn2 = 32'd0; 
32'd11511: dataIn2 = 32'd1; 
32'd11512: dataIn2 = 32'd1; 
32'd11513: dataIn2 = 32'd0; 
32'd11514: dataIn2 = 32'd0; 
32'd11515: dataIn2 = 32'd1; 
32'd11516: dataIn2 = 32'd1; 
32'd11517: dataIn2 = 32'd1; 
32'd11518: dataIn2 = 32'd1; 
32'd11519: dataIn2 = 32'd0; 
32'd11520: dataIn2 = 32'd1; 
32'd11521: dataIn2 = 32'd0; 
32'd11522: dataIn2 = 32'd1; 
32'd11523: dataIn2 = 32'd0; 
32'd11524: dataIn2 = 32'd0; 
32'd11525: dataIn2 = 32'd1; 
32'd11526: dataIn2 = 32'd0; 
32'd11527: dataIn2 = 32'd0; 
32'd11528: dataIn2 = 32'd0; 
32'd11529: dataIn2 = 32'd0; 
32'd11530: dataIn2 = 32'd1; 
32'd11531: dataIn2 = 32'd0; 
32'd11532: dataIn2 = 32'd1; 
32'd11533: dataIn2 = 32'd0; 
32'd11534: dataIn2 = 32'd1; 
32'd11535: dataIn2 = 32'd1; 
32'd11536: dataIn2 = 32'd0; 
32'd11537: dataIn2 = 32'd1; 
32'd11538: dataIn2 = 32'd0; 
32'd11539: dataIn2 = 32'd0; 
32'd11540: dataIn2 = 32'd1; 
32'd11541: dataIn2 = 32'd0; 
32'd11542: dataIn2 = 32'd1; 
32'd11543: dataIn2 = 32'd1; 
32'd11544: dataIn2 = 32'd1; 
32'd11545: dataIn2 = 32'd1; 
32'd11546: dataIn2 = 32'd0; 
32'd11547: dataIn2 = 32'd1; 
32'd11548: dataIn2 = 32'd0; 
32'd11549: dataIn2 = 32'd1; 
32'd11550: dataIn2 = 32'd1; 
32'd11551: dataIn2 = 32'd0; 
32'd11552: dataIn2 = 32'd1; 
32'd11553: dataIn2 = 32'd0; 
32'd11554: dataIn2 = 32'd1; 
32'd11555: dataIn2 = 32'd0; 
32'd11556: dataIn2 = 32'd1; 
32'd11557: dataIn2 = 32'd1; 
32'd11558: dataIn2 = 32'd0; 
32'd11559: dataIn2 = 32'd1; 
32'd11560: dataIn2 = 32'd0; 
32'd11561: dataIn2 = 32'd1; 
32'd11562: dataIn2 = 32'd0; 
32'd11563: dataIn2 = 32'd0; 
32'd11564: dataIn2 = 32'd0; 
32'd11565: dataIn2 = 32'd0; 
32'd11566: dataIn2 = 32'd0; 
32'd11567: dataIn2 = 32'd0; 
32'd11568: dataIn2 = 32'd1; 
32'd11569: dataIn2 = 32'd0; 
32'd11570: dataIn2 = 32'd0; 
32'd11571: dataIn2 = 32'd1; 
32'd11572: dataIn2 = 32'd1; 
32'd11573: dataIn2 = 32'd1; 
32'd11574: dataIn2 = 32'd0; 
32'd11575: dataIn2 = 32'd0; 
32'd11576: dataIn2 = 32'd0; 
32'd11577: dataIn2 = 32'd1; 
32'd11578: dataIn2 = 32'd1; 
32'd11579: dataIn2 = 32'd0; 
32'd11580: dataIn2 = 32'd1; 
32'd11581: dataIn2 = 32'd0; 
32'd11582: dataIn2 = 32'd0; 
32'd11583: dataIn2 = 32'd1; 
32'd11584: dataIn2 = 32'd0; 
32'd11585: dataIn2 = 32'd1; 
32'd11586: dataIn2 = 32'd1; 
32'd11587: dataIn2 = 32'd1; 
32'd11588: dataIn2 = 32'd1; 
32'd11589: dataIn2 = 32'd1; 
32'd11590: dataIn2 = 32'd0; 
32'd11591: dataIn2 = 32'd0; 
32'd11592: dataIn2 = 32'd1; 
32'd11593: dataIn2 = 32'd0; 
32'd11594: dataIn2 = 32'd1; 
32'd11595: dataIn2 = 32'd0; 
32'd11596: dataIn2 = 32'd0; 
32'd11597: dataIn2 = 32'd0; 
32'd11598: dataIn2 = 32'd1; 
32'd11599: dataIn2 = 32'd0; 
32'd11600: dataIn2 = 32'd0; 
32'd11601: dataIn2 = 32'd0; 
32'd11602: dataIn2 = 32'd0; 
32'd11603: dataIn2 = 32'd1; 
32'd11604: dataIn2 = 32'd0; 
32'd11605: dataIn2 = 32'd1; 
32'd11606: dataIn2 = 32'd1; 
32'd11607: dataIn2 = 32'd1; 
32'd11608: dataIn2 = 32'd1; 
32'd11609: dataIn2 = 32'd0; 
32'd11610: dataIn2 = 32'd0; 
32'd11611: dataIn2 = 32'd1; 
32'd11612: dataIn2 = 32'd0; 
32'd11613: dataIn2 = 32'd1; 
32'd11614: dataIn2 = 32'd0; 
32'd11615: dataIn2 = 32'd1; 
32'd11616: dataIn2 = 32'd1; 
32'd11617: dataIn2 = 32'd0; 
32'd11618: dataIn2 = 32'd0; 
32'd11619: dataIn2 = 32'd1; 
32'd11620: dataIn2 = 32'd1; 
32'd11621: dataIn2 = 32'd1; 
32'd11622: dataIn2 = 32'd1; 
32'd11623: dataIn2 = 32'd1; 
32'd11624: dataIn2 = 32'd1; 
32'd11625: dataIn2 = 32'd1; 
32'd11626: dataIn2 = 32'd1; 
32'd11627: dataIn2 = 32'd1; 
32'd11628: dataIn2 = 32'd0; 
32'd11629: dataIn2 = 32'd0; 
32'd11630: dataIn2 = 32'd1; 
32'd11631: dataIn2 = 32'd1; 
32'd11632: dataIn2 = 32'd1; 
32'd11633: dataIn2 = 32'd1; 
32'd11634: dataIn2 = 32'd1; 
32'd11635: dataIn2 = 32'd1; 
32'd11636: dataIn2 = 32'd0; 
32'd11637: dataIn2 = 32'd1; 
32'd11638: dataIn2 = 32'd1; 
32'd11639: dataIn2 = 32'd0; 
32'd11640: dataIn2 = 32'd1; 
32'd11641: dataIn2 = 32'd0; 
32'd11642: dataIn2 = 32'd1; 
32'd11643: dataIn2 = 32'd1; 
32'd11644: dataIn2 = 32'd1; 
32'd11645: dataIn2 = 32'd1; 
32'd11646: dataIn2 = 32'd0; 
32'd11647: dataIn2 = 32'd1; 
32'd11648: dataIn2 = 32'd1; 
32'd11649: dataIn2 = 32'd0; 
32'd11650: dataIn2 = 32'd0; 
32'd11651: dataIn2 = 32'd1; 
32'd11652: dataIn2 = 32'd0; 
32'd11653: dataIn2 = 32'd1; 
32'd11654: dataIn2 = 32'd0; 
32'd11655: dataIn2 = 32'd0; 
32'd11656: dataIn2 = 32'd1; 
32'd11657: dataIn2 = 32'd0; 
32'd11658: dataIn2 = 32'd1; 
32'd11659: dataIn2 = 32'd0; 
32'd11660: dataIn2 = 32'd1; 
32'd11661: dataIn2 = 32'd1; 
32'd11662: dataIn2 = 32'd1; 
32'd11663: dataIn2 = 32'd0; 
32'd11664: dataIn2 = 32'd0; 
32'd11665: dataIn2 = 32'd0; 
32'd11666: dataIn2 = 32'd0; 
32'd11667: dataIn2 = 32'd0; 
32'd11668: dataIn2 = 32'd1; 
32'd11669: dataIn2 = 32'd1; 
32'd11670: dataIn2 = 32'd0; 
32'd11671: dataIn2 = 32'd1; 
32'd11672: dataIn2 = 32'd1; 
32'd11673: dataIn2 = 32'd0; 
32'd11674: dataIn2 = 32'd1; 
32'd11675: dataIn2 = 32'd0; 
32'd11676: dataIn2 = 32'd1; 
32'd11677: dataIn2 = 32'd0; 
32'd11678: dataIn2 = 32'd0; 
32'd11679: dataIn2 = 32'd0; 
32'd11680: dataIn2 = 32'd1; 
32'd11681: dataIn2 = 32'd0; 
32'd11682: dataIn2 = 32'd1; 
32'd11683: dataIn2 = 32'd0; 
32'd11684: dataIn2 = 32'd1; 
32'd11685: dataIn2 = 32'd1; 
32'd11686: dataIn2 = 32'd0; 
32'd11687: dataIn2 = 32'd0; 
32'd11688: dataIn2 = 32'd1; 
32'd11689: dataIn2 = 32'd0; 
32'd11690: dataIn2 = 32'd0; 
32'd11691: dataIn2 = 32'd1; 
32'd11692: dataIn2 = 32'd0; 
32'd11693: dataIn2 = 32'd1; 
32'd11694: dataIn2 = 32'd1; 
32'd11695: dataIn2 = 32'd0; 
32'd11696: dataIn2 = 32'd0; 
32'd11697: dataIn2 = 32'd0; 
32'd11698: dataIn2 = 32'd0; 
32'd11699: dataIn2 = 32'd1; 
32'd11700: dataIn2 = 32'd0; 
32'd11701: dataIn2 = 32'd0; 
32'd11702: dataIn2 = 32'd0; 
32'd11703: dataIn2 = 32'd1; 
32'd11704: dataIn2 = 32'd0; 
32'd11705: dataIn2 = 32'd0; 
32'd11706: dataIn2 = 32'd1; 
32'd11707: dataIn2 = 32'd1; 
32'd11708: dataIn2 = 32'd0; 
32'd11709: dataIn2 = 32'd1; 
32'd11710: dataIn2 = 32'd0; 
32'd11711: dataIn2 = 32'd0; 
32'd11712: dataIn2 = 32'd0; 
32'd11713: dataIn2 = 32'd1; 
32'd11714: dataIn2 = 32'd1; 
32'd11715: dataIn2 = 32'd1; 
32'd11716: dataIn2 = 32'd0; 
32'd11717: dataIn2 = 32'd0; 
32'd11718: dataIn2 = 32'd1; 
32'd11719: dataIn2 = 32'd1; 
32'd11720: dataIn2 = 32'd0; 
32'd11721: dataIn2 = 32'd1; 
32'd11722: dataIn2 = 32'd0; 
32'd11723: dataIn2 = 32'd0; 
32'd11724: dataIn2 = 32'd1; 
32'd11725: dataIn2 = 32'd0; 
32'd11726: dataIn2 = 32'd0; 
32'd11727: dataIn2 = 32'd1; 
32'd11728: dataIn2 = 32'd0; 
32'd11729: dataIn2 = 32'd0; 
32'd11730: dataIn2 = 32'd1; 
32'd11731: dataIn2 = 32'd1; 
32'd11732: dataIn2 = 32'd0; 
32'd11733: dataIn2 = 32'd0; 
32'd11734: dataIn2 = 32'd0; 
32'd11735: dataIn2 = 32'd0; 
32'd11736: dataIn2 = 32'd1; 
32'd11737: dataIn2 = 32'd0; 
32'd11738: dataIn2 = 32'd0; 
32'd11739: dataIn2 = 32'd0; 
default: 
	dataIn2 = 32'd99999; 
endcase 
end 
always begin 
#10 Clk = ~Clk; 
end 
//========== VCD ============ 
`ifdef VCD 
initial 
begin 
	$dumpfile("pesa.vcd");  
	$dumpvars; 
end 
`endif 
//===========RTLVCD ========== 
`ifdef RTLVCD 
initial 
begin 
	$dumpfile("hht_rtl.vcd"); 
	$dumpvars; 
end 
`endif 
endmodule 
